magic
tech sky130A
magscale 1 2
timestamp 1653997641
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 219342 700408 219348 700460
rect 219400 700448 219406 700460
rect 267642 700448 267648 700460
rect 219400 700420 267648 700448
rect 219400 700408 219406 700420
rect 267642 700408 267648 700420
rect 267700 700408 267706 700460
rect 217962 700340 217968 700392
rect 218020 700380 218026 700392
rect 283834 700380 283840 700392
rect 218020 700352 283840 700380
rect 218020 700340 218026 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 348786 700340 348792 700392
rect 348844 700380 348850 700392
rect 358814 700380 358820 700392
rect 348844 700352 358820 700380
rect 348844 700340 348850 700352
rect 358814 700340 358820 700352
rect 358872 700340 358878 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 98638 700312 98644 700324
rect 8168 700284 98644 700312
rect 8168 700272 8174 700284
rect 98638 700272 98644 700284
rect 98696 700272 98702 700324
rect 217870 700272 217876 700324
rect 217928 700312 217934 700324
rect 300118 700312 300124 700324
rect 217928 700284 300124 700312
rect 217928 700272 217934 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 357434 700312 357440 700324
rect 332560 700284 357440 700312
rect 332560 700272 332566 700284
rect 357434 700272 357440 700284
rect 357492 700272 357498 700324
rect 359458 700272 359464 700324
rect 359516 700312 359522 700324
rect 429838 700312 429844 700324
rect 359516 700284 429844 700312
rect 359516 700272 359522 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 442258 700272 442264 700324
rect 442316 700312 442322 700324
rect 559650 700312 559656 700324
rect 442316 700284 559656 700312
rect 442316 700272 442322 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 105446 699728 105452 699780
rect 105504 699768 105510 699780
rect 108298 699768 108304 699780
rect 105504 699740 108304 699768
rect 105504 699728 105510 699740
rect 108298 699728 108304 699740
rect 108356 699728 108362 699780
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 137830 699660 137836 699712
rect 137888 699700 137894 699712
rect 140038 699700 140044 699712
rect 137888 699672 140044 699700
rect 137888 699660 137894 699672
rect 140038 699660 140044 699672
rect 140096 699660 140102 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 391198 696940 391204 696992
rect 391256 696980 391262 696992
rect 580166 696980 580172 696992
rect 391256 696952 580172 696980
rect 391256 696940 391262 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 21358 683176 21364 683188
rect 3476 683148 21364 683176
rect 3476 683136 3482 683148
rect 21358 683136 21364 683148
rect 21416 683136 21422 683188
rect 381538 683136 381544 683188
rect 381596 683176 381602 683188
rect 580166 683176 580172 683188
rect 381596 683148 580172 683176
rect 381596 683136 381602 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 215938 670732 215944 670744
rect 3568 670704 215944 670732
rect 3568 670692 3574 670704
rect 215938 670692 215944 670704
rect 215996 670692 216002 670744
rect 377398 670692 377404 670744
rect 377456 670732 377462 670744
rect 580166 670732 580172 670744
rect 377456 670704 580172 670732
rect 377456 670692 377462 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 28258 656928 28264 656940
rect 3476 656900 28264 656928
rect 3476 656888 3482 656900
rect 28258 656888 28264 656900
rect 28316 656888 28322 656940
rect 373258 643084 373264 643136
rect 373316 643124 373322 643136
rect 580166 643124 580172 643136
rect 373316 643096 580172 643124
rect 373316 643084 373322 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 214558 618304 214564 618316
rect 3200 618276 214564 618304
rect 3200 618264 3206 618276
rect 214558 618264 214564 618276
rect 214616 618264 214622 618316
rect 363598 616836 363604 616888
rect 363656 616876 363662 616888
rect 580166 616876 580172 616888
rect 363656 616848 580172 616876
rect 363656 616836 363662 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 606024 3424 606076
rect 3476 606064 3482 606076
rect 7558 606064 7564 606076
rect 3476 606036 7564 606064
rect 3476 606024 3482 606036
rect 7558 606024 7564 606036
rect 7616 606024 7622 606076
rect 374638 590656 374644 590708
rect 374696 590696 374702 590708
rect 580166 590696 580172 590708
rect 374696 590668 580172 590696
rect 374696 590656 374702 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 57238 579680 57244 579692
rect 3384 579652 57244 579680
rect 3384 579640 3390 579652
rect 57238 579640 57244 579652
rect 57296 579640 57302 579692
rect 378778 576852 378784 576904
rect 378836 576892 378842 576904
rect 580166 576892 580172 576904
rect 378836 576864 580172 576892
rect 378836 576852 378842 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 211798 565876 211804 565888
rect 3476 565848 211804 565876
rect 3476 565836 3482 565848
rect 211798 565836 211804 565848
rect 211856 565836 211862 565888
rect 217778 565088 217784 565140
rect 217836 565128 217842 565140
rect 234614 565128 234620 565140
rect 217836 565100 234620 565128
rect 217836 565088 217842 565100
rect 234614 565088 234620 565100
rect 234672 565088 234678 565140
rect 367738 563048 367744 563100
rect 367796 563088 367802 563100
rect 580166 563088 580172 563100
rect 367796 563060 580172 563088
rect 367796 563048 367802 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3418 553664 3424 553716
rect 3476 553704 3482 553716
rect 8938 553704 8944 553716
rect 3476 553676 8944 553704
rect 3476 553664 3482 553676
rect 8938 553664 8944 553676
rect 8996 553664 9002 553716
rect 369118 536800 369124 536852
rect 369176 536840 369182 536852
rect 579890 536840 579896 536852
rect 369176 536812 579896 536840
rect 369176 536800 369182 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 35158 527184 35164 527196
rect 3476 527156 35164 527184
rect 3476 527144 3482 527156
rect 35158 527144 35164 527156
rect 35216 527144 35222 527196
rect 371878 524424 371884 524476
rect 371936 524464 371942 524476
rect 580166 524464 580172 524476
rect 371936 524436 580172 524464
rect 371936 524424 371942 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 210418 514808 210424 514820
rect 3476 514780 210424 514808
rect 3476 514768 3482 514780
rect 210418 514768 210424 514780
rect 210476 514768 210482 514820
rect 358078 510620 358084 510672
rect 358136 510660 358142 510672
rect 580166 510660 580172 510672
rect 358136 510632 580172 510660
rect 358136 510620 358142 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 13078 501004 13084 501016
rect 3108 500976 13084 501004
rect 3108 500964 3114 500976
rect 13078 500964 13084 500976
rect 13136 500964 13142 501016
rect 360838 484372 360844 484424
rect 360896 484412 360902 484424
rect 580166 484412 580172 484424
rect 360896 484384 580172 484412
rect 360896 484372 360902 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 217870 478592 217876 478644
rect 217928 478632 217934 478644
rect 269942 478632 269948 478644
rect 217928 478604 269948 478632
rect 217928 478592 217934 478604
rect 269942 478592 269948 478604
rect 270000 478592 270006 478644
rect 217962 478524 217968 478576
rect 218020 478564 218026 478576
rect 271230 478564 271236 478576
rect 218020 478536 271236 478564
rect 218020 478524 218026 478536
rect 271230 478524 271236 478536
rect 271288 478524 271294 478576
rect 268654 478456 268660 478508
rect 268712 478496 268718 478508
rect 357434 478496 357440 478508
rect 268712 478468 357440 478496
rect 268712 478456 268718 478468
rect 357434 478456 357440 478468
rect 357492 478456 357498 478508
rect 269298 478388 269304 478440
rect 269356 478428 269362 478440
rect 358814 478428 358820 478440
rect 269356 478400 358820 478428
rect 269356 478388 269362 478400
rect 358814 478388 358820 478400
rect 358872 478388 358878 478440
rect 217410 478320 217416 478372
rect 217468 478360 217474 478372
rect 308582 478360 308588 478372
rect 217468 478332 308588 478360
rect 217468 478320 217474 478332
rect 308582 478320 308588 478332
rect 308640 478320 308646 478372
rect 218974 478252 218980 478304
rect 219032 478292 219038 478304
rect 314470 478292 314476 478304
rect 219032 478264 314476 478292
rect 219032 478252 219038 478264
rect 314470 478252 314476 478264
rect 314528 478252 314534 478304
rect 256878 478184 256884 478236
rect 256936 478224 256942 478236
rect 374638 478224 374644 478236
rect 256936 478196 374644 478224
rect 256936 478184 256942 478196
rect 374638 478184 374644 478196
rect 374696 478184 374702 478236
rect 7558 478116 7564 478168
rect 7616 478156 7622 478168
rect 282362 478156 282368 478168
rect 7616 478128 282368 478156
rect 7616 478116 7622 478128
rect 282362 478116 282368 478128
rect 282420 478116 282426 478168
rect 241422 476824 241428 476876
rect 241480 476864 241486 476876
rect 241480 476836 248414 476864
rect 241480 476824 241486 476836
rect 238478 476756 238484 476808
rect 238536 476796 238542 476808
rect 248386 476796 248414 476836
rect 316402 476796 316408 476808
rect 238536 476768 243584 476796
rect 248386 476768 316408 476796
rect 238536 476756 238542 476768
rect 237282 476688 237288 476740
rect 237340 476728 237346 476740
rect 239398 476728 239404 476740
rect 237340 476700 239404 476728
rect 237340 476688 237346 476700
rect 239398 476688 239404 476700
rect 239456 476688 239462 476740
rect 243556 476728 243584 476768
rect 316402 476756 316408 476768
rect 316460 476756 316466 476808
rect 311250 476728 311256 476740
rect 243556 476700 311256 476728
rect 311250 476688 311256 476700
rect 311308 476688 311314 476740
rect 242802 476620 242808 476672
rect 242860 476660 242866 476672
rect 319070 476660 319076 476672
rect 242860 476632 319076 476660
rect 242860 476620 242866 476632
rect 319070 476620 319076 476632
rect 319128 476620 319134 476672
rect 271782 476552 271788 476604
rect 271840 476592 271846 476604
rect 330202 476592 330208 476604
rect 271840 476564 330208 476592
rect 271840 476552 271846 476564
rect 330202 476552 330208 476564
rect 330260 476552 330266 476604
rect 266262 476484 266268 476536
rect 266320 476524 266326 476536
rect 326890 476524 326896 476536
rect 266320 476496 326896 476524
rect 266320 476484 266326 476496
rect 326890 476484 326896 476496
rect 326948 476484 326954 476536
rect 256602 476416 256608 476468
rect 256660 476456 256666 476468
rect 318426 476456 318432 476468
rect 256660 476428 318432 476456
rect 256660 476416 256666 476428
rect 318426 476416 318432 476428
rect 318484 476416 318490 476468
rect 318702 476416 318708 476468
rect 318760 476456 318766 476468
rect 335998 476456 336004 476468
rect 318760 476428 336004 476456
rect 318760 476416 318766 476428
rect 335998 476416 336004 476428
rect 336056 476416 336062 476468
rect 262122 476348 262128 476400
rect 262180 476388 262186 476400
rect 323026 476388 323032 476400
rect 262180 476360 323032 476388
rect 262180 476348 262186 476360
rect 323026 476348 323032 476360
rect 323084 476348 323090 476400
rect 326982 476348 326988 476400
rect 327040 476388 327046 476400
rect 338758 476388 338764 476400
rect 327040 476360 338764 476388
rect 327040 476348 327046 476360
rect 338758 476348 338764 476360
rect 338816 476348 338822 476400
rect 309042 476280 309048 476332
rect 309100 476320 309106 476332
rect 329098 476320 329104 476332
rect 309100 476292 329104 476320
rect 309100 476280 309106 476292
rect 329098 476280 329104 476292
rect 329156 476280 329162 476332
rect 311802 476212 311808 476264
rect 311860 476252 311866 476264
rect 331858 476252 331864 476264
rect 311860 476224 331864 476252
rect 311860 476212 311866 476224
rect 331858 476212 331864 476224
rect 331916 476212 331922 476264
rect 315942 476144 315948 476196
rect 316000 476184 316006 476196
rect 334618 476184 334624 476196
rect 316000 476156 334624 476184
rect 316000 476144 316006 476156
rect 334618 476144 334624 476156
rect 334676 476144 334682 476196
rect 240042 476076 240048 476128
rect 240100 476116 240106 476128
rect 313826 476116 313832 476128
rect 240100 476088 313832 476116
rect 240100 476076 240106 476088
rect 313826 476076 313832 476088
rect 313884 476076 313890 476128
rect 314562 476076 314568 476128
rect 314620 476116 314626 476128
rect 333238 476116 333244 476128
rect 314620 476088 333244 476116
rect 314620 476076 314626 476088
rect 333238 476076 333244 476088
rect 333296 476076 333302 476128
rect 321462 475532 321468 475584
rect 321520 475572 321526 475584
rect 355318 475572 355324 475584
rect 321520 475544 355324 475572
rect 321520 475532 321526 475544
rect 355318 475532 355324 475544
rect 355376 475532 355382 475584
rect 274542 475464 274548 475516
rect 274600 475504 274606 475516
rect 331490 475504 331496 475516
rect 274600 475476 331496 475504
rect 274600 475464 274606 475476
rect 331490 475464 331496 475476
rect 331548 475464 331554 475516
rect 219158 475396 219164 475448
rect 219216 475436 219222 475448
rect 321646 475436 321652 475448
rect 219216 475408 321652 475436
rect 219216 475396 219222 475408
rect 321646 475396 321652 475408
rect 321704 475396 321710 475448
rect 255590 475328 255596 475380
rect 255648 475368 255654 475380
rect 371878 475368 371884 475380
rect 255648 475340 371884 475368
rect 255648 475328 255654 475340
rect 371878 475328 371884 475340
rect 371936 475328 371942 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 287606 474756 287612 474768
rect 3476 474728 287612 474756
rect 3476 474716 3482 474728
rect 287606 474716 287612 474728
rect 287664 474716 287670 474768
rect 264790 474240 264796 474292
rect 264848 474280 264854 474292
rect 297358 474280 297364 474292
rect 264848 474252 297364 474280
rect 264848 474240 264854 474252
rect 297358 474240 297364 474252
rect 297416 474240 297422 474292
rect 274450 474172 274456 474224
rect 274508 474212 274514 474224
rect 353110 474212 353116 474224
rect 274508 474184 353116 474212
rect 274508 474172 274514 474184
rect 353110 474172 353116 474184
rect 353168 474172 353174 474224
rect 219066 474104 219072 474156
rect 219124 474144 219130 474156
rect 317138 474144 317144 474156
rect 219124 474116 317144 474144
rect 219124 474104 219130 474116
rect 317138 474104 317144 474116
rect 317196 474104 317202 474156
rect 252922 474036 252928 474088
rect 252980 474076 252986 474088
rect 360838 474076 360844 474088
rect 252980 474048 360844 474076
rect 252980 474036 252986 474048
rect 360838 474036 360844 474048
rect 360896 474036 360902 474088
rect 153194 473968 153200 474020
rect 153252 474008 153258 474020
rect 275186 474008 275192 474020
rect 153252 473980 275192 474008
rect 153252 473968 153258 473980
rect 275186 473968 275192 473980
rect 275244 473968 275250 474020
rect 253750 472812 253756 472864
rect 253808 472852 253814 472864
rect 329558 472852 329564 472864
rect 253808 472824 329564 472852
rect 253808 472812 253814 472824
rect 329558 472812 329564 472824
rect 329616 472812 329622 472864
rect 217502 472744 217508 472796
rect 217560 472784 217566 472796
rect 323670 472784 323676 472796
rect 217560 472756 323676 472784
rect 217560 472744 217566 472756
rect 323670 472744 323676 472756
rect 323728 472744 323734 472796
rect 254854 472676 254860 472728
rect 254912 472716 254918 472728
rect 369118 472716 369124 472728
rect 254912 472688 369124 472716
rect 254912 472676 254918 472688
rect 369118 472676 369124 472688
rect 369176 472676 369182 472728
rect 8938 472608 8944 472660
rect 8996 472648 9002 472660
rect 284386 472648 284392 472660
rect 8996 472620 284392 472648
rect 8996 472608 9002 472620
rect 284386 472608 284392 472620
rect 284444 472608 284450 472660
rect 302142 472608 302148 472660
rect 302200 472648 302206 472660
rect 345934 472648 345940 472660
rect 302200 472620 345940 472648
rect 302200 472608 302206 472620
rect 345934 472608 345940 472620
rect 345992 472608 345998 472660
rect 259270 471384 259276 471436
rect 259328 471424 259334 471436
rect 294598 471424 294604 471436
rect 259328 471396 294604 471424
rect 259328 471384 259334 471396
rect 294598 471384 294604 471396
rect 294656 471384 294662 471436
rect 217594 471316 217600 471368
rect 217652 471356 217658 471368
rect 327534 471356 327540 471368
rect 217652 471328 327540 471356
rect 217652 471316 217658 471328
rect 327534 471316 327540 471328
rect 327592 471316 327598 471368
rect 13078 471248 13084 471300
rect 13136 471288 13142 471300
rect 286318 471288 286324 471300
rect 13136 471260 286324 471288
rect 13136 471248 13142 471260
rect 286318 471248 286324 471260
rect 286376 471248 286382 471300
rect 286502 471248 286508 471300
rect 286560 471288 286566 471300
rect 338022 471288 338028 471300
rect 286560 471260 338028 471288
rect 286560 471248 286566 471260
rect 338022 471248 338028 471260
rect 338080 471248 338086 471300
rect 253566 470568 253572 470620
rect 253624 470608 253630 470620
rect 580166 470608 580172 470620
rect 253624 470580 580172 470608
rect 253624 470568 253630 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 248230 470024 248236 470076
rect 248288 470064 248294 470076
rect 310514 470064 310520 470076
rect 248288 470036 310520 470064
rect 248288 470024 248294 470036
rect 310514 470024 310520 470036
rect 310572 470024 310578 470076
rect 257982 469956 257988 470008
rect 258040 469996 258046 470008
rect 333422 469996 333428 470008
rect 258040 469968 333428 469996
rect 258040 469956 258046 469968
rect 333422 469956 333428 469968
rect 333480 469956 333486 470008
rect 257522 469888 257528 469940
rect 257580 469928 257586 469940
rect 378778 469928 378784 469940
rect 257580 469900 378784 469928
rect 257580 469888 257586 469900
rect 378778 469888 378784 469900
rect 378836 469888 378842 469940
rect 35158 469820 35164 469872
rect 35216 469860 35222 469872
rect 285674 469860 285680 469872
rect 35216 469832 285680 469860
rect 35216 469820 35222 469832
rect 285674 469820 285680 469832
rect 285732 469820 285738 469872
rect 293862 469820 293868 469872
rect 293920 469860 293926 469872
rect 341978 469860 341984 469872
rect 293920 469832 341984 469860
rect 293920 469820 293926 469832
rect 341978 469820 341984 469832
rect 342036 469820 342042 469872
rect 253842 468732 253848 468784
rect 253900 468772 253906 468784
rect 301498 468772 301504 468784
rect 253900 468744 301504 468772
rect 253900 468732 253906 468744
rect 301498 468732 301504 468744
rect 301556 468732 301562 468784
rect 280062 468664 280068 468716
rect 280120 468704 280126 468716
rect 356698 468704 356704 468716
rect 280120 468676 356704 468704
rect 280120 468664 280126 468676
rect 356698 468664 356704 468676
rect 356756 468664 356762 468716
rect 219250 468596 219256 468648
rect 219308 468636 219314 468648
rect 319714 468636 319720 468648
rect 219308 468608 319720 468636
rect 219308 468596 219314 468608
rect 319714 468596 319720 468608
rect 319772 468596 319778 468648
rect 264698 468528 264704 468580
rect 264756 468568 264762 468580
rect 462314 468568 462320 468580
rect 264756 468540 462320 468568
rect 264756 468528 264762 468540
rect 462314 468528 462320 468540
rect 462372 468528 462378 468580
rect 57238 468460 57244 468512
rect 57296 468500 57302 468512
rect 283742 468500 283748 468512
rect 57296 468472 283748 468500
rect 57296 468460 57302 468472
rect 283742 468460 283748 468472
rect 283800 468460 283806 468512
rect 248322 467304 248328 467356
rect 248380 467344 248386 467356
rect 320358 467344 320364 467356
rect 248380 467316 320364 467344
rect 248380 467304 248386 467316
rect 320358 467304 320364 467316
rect 320416 467304 320422 467356
rect 217686 467236 217692 467288
rect 217744 467276 217750 467288
rect 325602 467276 325608 467288
rect 217744 467248 325608 467276
rect 217744 467236 217750 467248
rect 325602 467236 325608 467248
rect 325660 467236 325666 467288
rect 262766 467168 262772 467220
rect 262824 467208 262830 467220
rect 527174 467208 527180 467220
rect 262824 467180 527180 467208
rect 262824 467168 262830 467180
rect 527174 467168 527180 467180
rect 527232 467168 527238 467220
rect 4798 467100 4804 467152
rect 4856 467140 4862 467152
rect 281718 467140 281724 467152
rect 4856 467112 281724 467140
rect 4856 467100 4862 467112
rect 281718 467100 281724 467112
rect 281776 467100 281782 467152
rect 299382 467100 299388 467152
rect 299440 467140 299446 467152
rect 344554 467140 344560 467152
rect 299440 467112 344560 467140
rect 299440 467100 299446 467112
rect 344554 467100 344560 467112
rect 344612 467100 344618 467152
rect 275922 465876 275928 465928
rect 275980 465916 275986 465928
rect 354398 465916 354404 465928
rect 275980 465888 354404 465916
rect 275980 465876 275986 465888
rect 354398 465876 354404 465888
rect 354456 465876 354462 465928
rect 218882 465808 218888 465860
rect 218940 465848 218946 465860
rect 307294 465848 307300 465860
rect 218940 465820 307300 465848
rect 218940 465808 218946 465820
rect 307294 465808 307300 465820
rect 307352 465808 307358 465860
rect 258810 465740 258816 465792
rect 258868 465780 258874 465792
rect 373258 465780 373264 465792
rect 258868 465752 373264 465780
rect 258868 465740 258874 465752
rect 373258 465740 373264 465752
rect 373316 465740 373322 465792
rect 21358 465672 21364 465724
rect 21416 465712 21422 465724
rect 279786 465712 279792 465724
rect 21416 465684 279792 465712
rect 21416 465672 21422 465684
rect 279786 465672 279792 465684
rect 279844 465672 279850 465724
rect 291102 465672 291108 465724
rect 291160 465712 291166 465724
rect 340690 465712 340696 465724
rect 291160 465684 340696 465712
rect 291160 465672 291166 465684
rect 340690 465672 340696 465684
rect 340748 465672 340754 465724
rect 246942 464448 246948 464500
rect 247000 464488 247006 464500
rect 317782 464488 317788 464500
rect 247000 464460 317788 464488
rect 247000 464448 247006 464460
rect 317782 464448 317788 464460
rect 317840 464448 317846 464500
rect 218054 464380 218060 464432
rect 218112 464420 218118 464432
rect 273254 464420 273260 464432
rect 218112 464392 273260 464420
rect 218112 464380 218118 464392
rect 273254 464380 273260 464392
rect 273312 464380 273318 464432
rect 274358 464380 274364 464432
rect 274416 464420 274422 464432
rect 351822 464420 351828 464432
rect 274416 464392 351828 464420
rect 274416 464380 274422 464392
rect 351822 464380 351828 464392
rect 351880 464380 351886 464432
rect 266722 464312 266728 464364
rect 266780 464352 266786 464364
rect 396718 464352 396724 464364
rect 266780 464324 396724 464352
rect 266780 464312 266786 464324
rect 396718 464312 396724 464324
rect 396776 464312 396782 464364
rect 324222 463156 324228 463208
rect 324280 463196 324286 463208
rect 357710 463196 357716 463208
rect 324280 463168 357716 463196
rect 324280 463156 324286 463168
rect 357710 463156 357716 463168
rect 357768 463156 357774 463208
rect 252370 463088 252376 463140
rect 252428 463128 252434 463140
rect 326246 463128 326252 463140
rect 252428 463100 326252 463128
rect 252428 463088 252434 463100
rect 326246 463088 326252 463100
rect 326304 463088 326310 463140
rect 255222 463020 255228 463072
rect 255280 463060 255286 463072
rect 330846 463060 330852 463072
rect 255280 463032 330852 463060
rect 255280 463020 255286 463032
rect 330846 463020 330852 463032
rect 330904 463020 330910 463072
rect 260834 462952 260840 463004
rect 260892 462992 260898 463004
rect 391198 462992 391204 463004
rect 260892 462964 391204 462992
rect 260892 462952 260898 462964
rect 391198 462952 391204 462964
rect 391256 462952 391262 463004
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 288986 462380 288992 462392
rect 3292 462352 288992 462380
rect 3292 462340 3298 462352
rect 288986 462340 288992 462352
rect 289044 462340 289050 462392
rect 211798 461796 211804 461848
rect 211856 461836 211862 461848
rect 285030 461836 285036 461848
rect 211856 461808 285036 461836
rect 211856 461796 211862 461808
rect 285030 461796 285036 461808
rect 285088 461796 285094 461848
rect 262030 461728 262036 461780
rect 262088 461768 262094 461780
rect 338666 461768 338672 461780
rect 262088 461740 338672 461768
rect 262088 461728 262094 461740
rect 338666 461728 338672 461740
rect 338724 461728 338730 461780
rect 268010 461660 268016 461712
rect 268068 461700 268074 461712
rect 364334 461700 364340 461712
rect 268068 461672 364340 461700
rect 268068 461660 268074 461672
rect 364334 461660 364340 461672
rect 364392 461660 364398 461712
rect 71774 461592 71780 461644
rect 71832 461632 71838 461644
rect 276474 461632 276480 461644
rect 71832 461604 276480 461632
rect 71832 461592 71838 461604
rect 276474 461592 276480 461604
rect 276532 461592 276538 461644
rect 288342 461592 288348 461644
rect 288400 461632 288406 461644
rect 339402 461632 339408 461644
rect 288400 461604 339408 461632
rect 288400 461592 288406 461604
rect 339402 461592 339408 461604
rect 339460 461592 339466 461644
rect 250990 460436 250996 460488
rect 251048 460476 251054 460488
rect 313182 460476 313188 460488
rect 251048 460448 313188 460476
rect 251048 460436 251054 460448
rect 313182 460436 313188 460448
rect 313240 460436 313246 460488
rect 239398 460368 239404 460420
rect 239456 460408 239462 460420
rect 309226 460408 309232 460420
rect 239456 460380 309232 460408
rect 239456 460368 239462 460380
rect 309226 460368 309232 460380
rect 309284 460368 309290 460420
rect 277210 460300 277216 460352
rect 277268 460340 277274 460352
rect 355686 460340 355692 460352
rect 277268 460312 355692 460340
rect 277268 460300 277274 460312
rect 355686 460300 355692 460312
rect 355744 460300 355750 460352
rect 265986 460232 265992 460284
rect 266044 460272 266050 460284
rect 359458 460272 359464 460284
rect 266044 460244 359464 460272
rect 266044 460232 266050 460244
rect 359458 460232 359464 460244
rect 359516 460232 359522 460284
rect 98638 460164 98644 460216
rect 98696 460204 98702 460216
rect 278498 460204 278504 460216
rect 98696 460176 278504 460204
rect 98696 460164 98702 460176
rect 278498 460164 278504 460176
rect 278556 460164 278562 460216
rect 215938 459008 215944 459060
rect 215996 459048 216002 459060
rect 281074 459048 281080 459060
rect 215996 459020 281080 459048
rect 215996 459008 216002 459020
rect 281074 459008 281080 459020
rect 281132 459008 281138 459060
rect 260650 458940 260656 458992
rect 260708 458980 260714 458992
rect 337378 458980 337384 458992
rect 260708 458952 337384 458980
rect 260708 458940 260714 458952
rect 337378 458940 337384 458952
rect 337436 458940 337442 458992
rect 140038 458872 140044 458924
rect 140096 458912 140102 458924
rect 274542 458912 274548 458924
rect 140096 458884 274548 458912
rect 140096 458872 140102 458884
rect 274542 458872 274548 458884
rect 274600 458872 274606 458924
rect 281442 458872 281448 458924
rect 281500 458912 281506 458924
rect 335446 458912 335452 458924
rect 281500 458884 335452 458912
rect 281500 458872 281506 458884
rect 335446 458872 335452 458884
rect 335504 458872 335510 458924
rect 264054 458804 264060 458856
rect 264112 458844 264118 458856
rect 494054 458844 494060 458856
rect 264112 458816 494060 458844
rect 264112 458804 264118 458816
rect 494054 458804 494060 458816
rect 494112 458804 494118 458856
rect 249702 457580 249708 457632
rect 249760 457620 249766 457632
rect 322290 457620 322296 457632
rect 249760 457592 322296 457620
rect 249760 457580 249766 457592
rect 322290 457580 322296 457592
rect 322348 457580 322354 457632
rect 256510 457512 256516 457564
rect 256568 457552 256574 457564
rect 332134 457552 332140 457564
rect 256568 457524 332140 457552
rect 256568 457512 256574 457524
rect 332134 457512 332140 457524
rect 332192 457512 332198 457564
rect 28258 457444 28264 457496
rect 28316 457484 28322 457496
rect 280430 457484 280436 457496
rect 28316 457456 280436 457484
rect 28316 457444 28322 457456
rect 280430 457444 280436 457456
rect 280488 457444 280494 457496
rect 306282 457444 306288 457496
rect 306340 457484 306346 457496
rect 348510 457484 348516 457496
rect 306340 457456 348516 457484
rect 306340 457444 306346 457456
rect 348510 457444 348516 457456
rect 348568 457444 348574 457496
rect 252278 456764 252284 456816
rect 252336 456804 252342 456816
rect 580166 456804 580172 456816
rect 252336 456776 580172 456804
rect 252336 456764 252342 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 201494 456220 201500 456272
rect 201552 456260 201558 456272
rect 272610 456260 272616 456272
rect 201552 456232 272616 456260
rect 201552 456220 201558 456232
rect 272610 456220 272616 456232
rect 272668 456220 272674 456272
rect 259362 456152 259368 456204
rect 259420 456192 259426 456204
rect 334802 456192 334808 456204
rect 259420 456164 334808 456192
rect 259420 456152 259426 456164
rect 334802 456152 334808 456164
rect 334860 456152 334866 456204
rect 262122 456084 262128 456136
rect 262180 456124 262186 456136
rect 442258 456124 442264 456136
rect 262180 456096 442264 456124
rect 262180 456084 262186 456096
rect 442258 456084 442264 456096
rect 442316 456084 442322 456136
rect 88334 456016 88340 456068
rect 88392 456056 88398 456068
rect 277118 456056 277124 456068
rect 88392 456028 277124 456056
rect 88392 456016 88398 456028
rect 277118 456016 277124 456028
rect 277176 456016 277182 456068
rect 277302 456016 277308 456068
rect 277360 456056 277366 456068
rect 332778 456056 332784 456068
rect 277360 456028 332784 456056
rect 277360 456016 277366 456028
rect 332778 456016 332784 456028
rect 332836 456016 332842 456068
rect 268930 454860 268936 454912
rect 268988 454900 268994 454912
rect 293218 454900 293224 454912
rect 268988 454872 293224 454900
rect 268988 454860 268994 454872
rect 293218 454860 293224 454872
rect 293276 454860 293282 454912
rect 296622 454860 296628 454912
rect 296680 454900 296686 454912
rect 343266 454900 343272 454912
rect 296680 454872 343272 454900
rect 296680 454860 296686 454872
rect 343266 454860 343272 454872
rect 343324 454860 343330 454912
rect 244182 454792 244188 454844
rect 244240 454832 244246 454844
rect 309870 454832 309876 454844
rect 244240 454804 309876 454832
rect 244240 454792 244246 454804
rect 309870 454792 309876 454804
rect 309928 454792 309934 454844
rect 260098 454724 260104 454776
rect 260156 454764 260162 454776
rect 377398 454764 377404 454776
rect 260156 454736 377404 454764
rect 260156 454724 260162 454736
rect 377398 454724 377404 454736
rect 377456 454724 377462 454776
rect 40034 454656 40040 454708
rect 40092 454696 40098 454708
rect 277854 454696 277860 454708
rect 40092 454668 277860 454696
rect 40092 454656 40098 454668
rect 277854 454656 277860 454668
rect 277912 454656 277918 454708
rect 278590 454656 278596 454708
rect 278648 454696 278654 454708
rect 357066 454696 357072 454708
rect 278648 454668 357072 454696
rect 278648 454656 278654 454668
rect 357066 454656 357072 454668
rect 357124 454656 357130 454708
rect 214558 453568 214564 453620
rect 214616 453608 214622 453620
rect 283006 453608 283012 453620
rect 214616 453580 283012 453608
rect 214616 453568 214622 453580
rect 283006 453568 283012 453580
rect 283064 453568 283070 453620
rect 251082 453500 251088 453552
rect 251140 453540 251146 453552
rect 324314 453540 324320 453552
rect 251140 453512 324320 453540
rect 251140 453500 251146 453512
rect 324314 453500 324320 453512
rect 324372 453500 324378 453552
rect 271690 453432 271696 453484
rect 271748 453472 271754 453484
rect 349154 453472 349160 453484
rect 271748 453444 349160 453472
rect 271748 453432 271754 453444
rect 349154 453432 349160 453444
rect 349212 453432 349218 453484
rect 169754 453364 169760 453416
rect 169812 453404 169818 453416
rect 273898 453404 273904 453416
rect 169812 453376 273904 453404
rect 169812 453364 169818 453376
rect 273898 453364 273904 453376
rect 273956 453364 273962 453416
rect 258166 453296 258172 453348
rect 258224 453336 258230 453348
rect 363598 453336 363604 453348
rect 258224 453308 363604 453336
rect 258224 453296 258230 453308
rect 363598 453296 363604 453308
rect 363656 453296 363662 453348
rect 252462 452140 252468 452192
rect 252520 452180 252526 452192
rect 328270 452180 328276 452192
rect 252520 452152 328276 452180
rect 252520 452140 252526 452152
rect 328270 452140 328276 452152
rect 328328 452140 328334 452192
rect 210418 452072 210424 452124
rect 210476 452112 210482 452124
rect 286962 452112 286968 452124
rect 210476 452084 286968 452112
rect 210476 452072 210482 452084
rect 286962 452072 286968 452084
rect 287020 452072 287026 452124
rect 273162 452004 273168 452056
rect 273220 452044 273226 452056
rect 350534 452044 350540 452056
rect 273220 452016 350540 452044
rect 273220 452004 273226 452016
rect 350534 452004 350540 452016
rect 350592 452004 350598 452056
rect 255958 451936 255964 451988
rect 256016 451976 256022 451988
rect 367738 451976 367744 451988
rect 256016 451948 367744 451976
rect 256016 451936 256022 451948
rect 367738 451936 367744 451948
rect 367796 451936 367802 451988
rect 108298 451868 108304 451920
rect 108356 451908 108362 451920
rect 275830 451908 275836 451920
rect 108356 451880 275836 451908
rect 108356 451868 108362 451880
rect 275830 451868 275836 451880
rect 275888 451868 275894 451920
rect 278682 450712 278688 450764
rect 278740 450752 278746 450764
rect 334158 450752 334164 450764
rect 278740 450724 334164 450752
rect 278740 450712 278746 450724
rect 334158 450712 334164 450724
rect 334216 450712 334222 450764
rect 254210 450644 254216 450696
rect 254268 450684 254274 450696
rect 358078 450684 358084 450696
rect 254268 450656 358084 450684
rect 254268 450644 254274 450656
rect 358078 450644 358084 450656
rect 358136 450644 358142 450696
rect 261478 450576 261484 450628
rect 261536 450616 261542 450628
rect 381538 450616 381544 450628
rect 261536 450588 381544 450616
rect 261536 450576 261542 450588
rect 381538 450576 381544 450588
rect 381596 450576 381602 450628
rect 25498 450508 25504 450560
rect 25556 450548 25562 450560
rect 279142 450548 279148 450560
rect 25556 450520 279148 450548
rect 25556 450508 25562 450520
rect 279142 450508 279148 450520
rect 279200 450508 279206 450560
rect 245470 449692 245476 449744
rect 245528 449732 245534 449744
rect 312538 449732 312544 449744
rect 245528 449704 312544 449732
rect 245528 449692 245534 449704
rect 312538 449692 312544 449704
rect 312596 449692 312602 449744
rect 245562 449624 245568 449676
rect 245620 449664 245626 449676
rect 315114 449664 315120 449676
rect 245620 449636 315120 449664
rect 245620 449624 245626 449636
rect 315114 449624 315120 449636
rect 315172 449624 315178 449676
rect 267642 449556 267648 449608
rect 267700 449596 267706 449608
rect 343910 449596 343916 449608
rect 267700 449568 343916 449596
rect 267700 449556 267706 449568
rect 343910 449556 343916 449568
rect 343968 449556 343974 449608
rect 266170 449488 266176 449540
rect 266228 449528 266234 449540
rect 342622 449528 342628 449540
rect 266228 449500 342628 449528
rect 266228 449488 266234 449500
rect 342622 449488 342628 449500
rect 342680 449488 342686 449540
rect 263502 449420 263508 449472
rect 263560 449460 263566 449472
rect 340046 449460 340052 449472
rect 263560 449432 340052 449460
rect 263560 449420 263566 449432
rect 340046 449420 340052 449432
rect 340104 449420 340110 449472
rect 264882 449352 264888 449404
rect 264940 449392 264946 449404
rect 341334 449392 341340 449404
rect 264940 449364 341340 449392
rect 264940 449352 264946 449364
rect 341334 449352 341340 449364
rect 341392 449352 341398 449404
rect 269022 449284 269028 449336
rect 269080 449324 269086 449336
rect 346578 449324 346584 449336
rect 269080 449296 346584 449324
rect 269080 449284 269086 449296
rect 346578 449284 346584 449296
rect 346636 449284 346642 449336
rect 270402 449216 270408 449268
rect 270460 449256 270466 449268
rect 347866 449256 347872 449268
rect 270460 449228 347872 449256
rect 270460 449216 270466 449228
rect 347866 449216 347872 449228
rect 347924 449216 347930 449268
rect 267550 449148 267556 449200
rect 267608 449188 267614 449200
rect 345290 449188 345296 449200
rect 267608 449160 345296 449188
rect 267608 449148 267614 449160
rect 345290 449148 345296 449160
rect 345348 449148 345354 449200
rect 303522 448060 303528 448112
rect 303580 448100 303586 448112
rect 347222 448100 347228 448112
rect 303580 448072 347228 448100
rect 303580 448060 303586 448072
rect 347222 448060 347228 448072
rect 347280 448060 347286 448112
rect 284202 447992 284208 448044
rect 284260 448032 284266 448044
rect 336734 448032 336740 448044
rect 284260 448004 336740 448032
rect 284260 447992 284266 448004
rect 336734 447992 336740 448004
rect 336792 447992 336798 448044
rect 237190 447924 237196 447976
rect 237248 447964 237254 447976
rect 311894 447964 311900 447976
rect 237248 447936 311900 447964
rect 237248 447924 237254 447936
rect 311894 447924 311900 447936
rect 311952 447924 311958 447976
rect 260742 447856 260748 447908
rect 260800 447896 260806 447908
rect 336090 447896 336096 447908
rect 260800 447868 336096 447896
rect 260800 447856 260806 447868
rect 336090 447856 336096 447868
rect 336148 447856 336154 447908
rect 217318 447788 217324 447840
rect 217376 447828 217382 447840
rect 307938 447828 307944 447840
rect 217376 447800 307944 447828
rect 217376 447788 217382 447800
rect 307938 447788 307944 447800
rect 307996 447788 308002 447840
rect 267366 446632 267372 446684
rect 267424 446672 267430 446684
rect 412634 446672 412640 446684
rect 267424 446644 412640 446672
rect 267424 446632 267430 446644
rect 412634 446632 412640 446644
rect 412692 446632 412698 446684
rect 265342 446564 265348 446616
rect 265400 446604 265406 446616
rect 477494 446604 477500 446616
rect 265400 446576 477500 446604
rect 265400 446564 265406 446576
rect 477494 446564 477500 446576
rect 477552 446564 477558 446616
rect 263410 446496 263416 446548
rect 263468 446536 263474 446548
rect 542354 446536 542360 446548
rect 263468 446508 542360 446536
rect 263468 446496 263474 446508
rect 542354 446496 542360 446508
rect 542412 446496 542418 446548
rect 4154 446428 4160 446480
rect 4212 446468 4218 446480
rect 288250 446468 288256 446480
rect 4212 446440 288256 446468
rect 4212 446428 4218 446440
rect 288250 446428 288256 446440
rect 288308 446428 288314 446480
rect 259454 446360 259460 446412
rect 259512 446400 259518 446412
rect 580258 446400 580264 446412
rect 259512 446372 580264 446400
rect 259512 446360 259518 446372
rect 580258 446360 580264 446372
rect 580316 446360 580322 446412
rect 203518 446156 203524 446208
rect 203576 446196 203582 446208
rect 300118 446196 300124 446208
rect 203576 446168 300124 446196
rect 203576 446156 203582 446168
rect 300118 446156 300124 446168
rect 300176 446156 300182 446208
rect 199378 446088 199384 446140
rect 199436 446128 199442 446140
rect 300762 446128 300768 446140
rect 199436 446100 300768 446128
rect 199436 446088 199442 446100
rect 300762 446088 300768 446100
rect 300820 446088 300826 446140
rect 200758 446020 200764 446072
rect 200816 446060 200822 446072
rect 306006 446060 306012 446072
rect 200816 446032 306012 446060
rect 200816 446020 200822 446032
rect 306006 446020 306012 446032
rect 306064 446020 306070 446072
rect 250990 445952 250996 446004
rect 251048 445992 251054 446004
rect 362586 445992 362592 446004
rect 251048 445964 362592 445992
rect 251048 445952 251054 445964
rect 362586 445952 362592 445964
rect 362644 445952 362650 446004
rect 249702 445884 249708 445936
rect 249760 445924 249766 445936
rect 363598 445924 363604 445936
rect 249760 445896 363604 445924
rect 249760 445884 249766 445896
rect 363598 445884 363604 445896
rect 363656 445884 363662 445936
rect 235902 445816 235908 445868
rect 235960 445856 235966 445868
rect 378778 445856 378784 445868
rect 235960 445828 378784 445856
rect 235960 445816 235966 445828
rect 378778 445816 378784 445828
rect 378836 445816 378842 445868
rect 82078 445748 82084 445800
rect 82136 445788 82142 445800
rect 303982 445788 303988 445800
rect 82136 445760 303988 445788
rect 82136 445748 82142 445760
rect 303982 445748 303988 445760
rect 304040 445748 304046 445800
rect 231118 444932 231124 444984
rect 231176 444972 231182 444984
rect 290274 444972 290280 444984
rect 231176 444944 290280 444972
rect 231176 444932 231182 444944
rect 290274 444932 290280 444944
rect 290332 444932 290338 444984
rect 225598 444864 225604 444916
rect 225656 444904 225662 444916
rect 295518 444904 295524 444916
rect 225656 444876 295524 444904
rect 225656 444864 225662 444876
rect 295518 444864 295524 444876
rect 295576 444864 295582 444916
rect 215938 444796 215944 444848
rect 215996 444836 216002 444848
rect 297450 444836 297456 444848
rect 215996 444808 297456 444836
rect 215996 444796 216002 444808
rect 297450 444796 297456 444808
rect 297508 444796 297514 444848
rect 245746 444728 245752 444780
rect 245804 444768 245810 444780
rect 374638 444768 374644 444780
rect 245804 444740 374644 444768
rect 245804 444728 245810 444740
rect 374638 444728 374644 444740
rect 374696 444728 374702 444780
rect 240502 444660 240508 444712
rect 240560 444700 240566 444712
rect 371970 444700 371976 444712
rect 240560 444672 371976 444700
rect 240560 444660 240566 444672
rect 371970 444660 371976 444672
rect 372028 444660 372034 444712
rect 100018 444592 100024 444644
rect 100076 444632 100082 444644
rect 291562 444632 291568 444644
rect 100076 444604 291568 444632
rect 100076 444592 100082 444604
rect 291562 444592 291568 444604
rect 291620 444592 291626 444644
rect 95878 444524 95884 444576
rect 95936 444564 95942 444576
rect 293494 444564 293500 444576
rect 95936 444536 293500 444564
rect 95936 444524 95942 444536
rect 293494 444524 293500 444536
rect 293552 444524 293558 444576
rect 7558 444456 7564 444508
rect 7616 444496 7622 444508
rect 289630 444496 289636 444508
rect 7616 444468 289636 444496
rect 7616 444456 7622 444468
rect 289630 444456 289636 444468
rect 289688 444456 289694 444508
rect 244458 444388 244464 444440
rect 244516 444428 244522 444440
rect 578878 444428 578884 444440
rect 244516 444400 578884 444428
rect 244516 444388 244522 444400
rect 578878 444388 578884 444400
rect 578936 444388 578942 444440
rect 355318 444320 355324 444372
rect 355376 444360 355382 444372
rect 356422 444360 356428 444372
rect 355376 444332 356428 444360
rect 355376 444320 355382 444332
rect 356422 444320 356428 444332
rect 356480 444320 356486 444372
rect 356698 444320 356704 444372
rect 356756 444360 356762 444372
rect 358354 444360 358360 444372
rect 356756 444332 358360 444360
rect 356756 444320 356762 444332
rect 358354 444320 358360 444332
rect 358412 444320 358418 444372
rect 248322 444116 248328 444168
rect 248380 444156 248386 444168
rect 362402 444156 362408 444168
rect 248380 444128 362408 444156
rect 248380 444116 248386 444128
rect 362402 444116 362408 444128
rect 362460 444116 362466 444168
rect 245102 444048 245108 444100
rect 245160 444088 245166 444100
rect 362218 444088 362224 444100
rect 245160 444060 362224 444088
rect 245160 444048 245166 444060
rect 362218 444048 362224 444060
rect 362276 444048 362282 444100
rect 334618 443980 334624 444032
rect 334676 444020 334682 444032
rect 353754 444020 353760 444032
rect 334676 443992 353760 444020
rect 334676 443980 334682 443992
rect 353754 443980 353760 443992
rect 353812 443980 353818 444032
rect 243078 443912 243084 443964
rect 243136 443952 243142 443964
rect 251174 443952 251180 443964
rect 243136 443924 251180 443952
rect 243136 443912 243142 443924
rect 251174 443912 251180 443924
rect 251232 443912 251238 443964
rect 333238 443912 333244 443964
rect 333296 443952 333302 443964
rect 352466 443952 352472 443964
rect 333296 443924 352472 443952
rect 333296 443912 333302 443924
rect 352466 443912 352472 443924
rect 352524 443912 352530 443964
rect 94498 443844 94504 443896
rect 94556 443884 94562 443896
rect 294874 443884 294880 443896
rect 94556 443856 294880 443884
rect 94556 443844 94562 443856
rect 294874 443844 294880 443856
rect 294932 443844 294938 443896
rect 301498 443844 301504 443896
rect 301556 443884 301562 443896
rect 315758 443884 315764 443896
rect 301556 443856 315764 443884
rect 301556 443844 301562 443856
rect 315758 443844 315764 443856
rect 315816 443844 315822 443896
rect 331858 443844 331864 443896
rect 331916 443884 331922 443896
rect 351178 443884 351184 443896
rect 331916 443856 351184 443884
rect 331916 443844 331922 443856
rect 351178 443844 351184 443856
rect 351236 443844 351242 443896
rect 230474 443776 230480 443828
rect 230532 443816 230538 443828
rect 259454 443816 259460 443828
rect 230532 443788 259460 443816
rect 230532 443776 230538 443788
rect 259454 443776 259460 443788
rect 259512 443776 259518 443828
rect 294598 443776 294604 443828
rect 294656 443816 294662 443828
rect 321002 443816 321008 443828
rect 294656 443788 321008 443816
rect 294656 443776 294662 443788
rect 321002 443776 321008 443788
rect 321060 443776 321066 443828
rect 335998 443776 336004 443828
rect 336056 443816 336062 443828
rect 355042 443816 355048 443828
rect 336056 443788 355048 443816
rect 336056 443776 336062 443788
rect 355042 443776 355048 443788
rect 355100 443776 355106 443828
rect 219342 443708 219348 443760
rect 219400 443748 219406 443760
rect 270586 443748 270592 443760
rect 219400 443720 270592 443748
rect 219400 443708 219406 443720
rect 270586 443708 270592 443720
rect 270644 443708 270650 443760
rect 297358 443708 297364 443760
rect 297416 443748 297422 443760
rect 324958 443748 324964 443760
rect 297416 443720 324964 443748
rect 297416 443708 297422 443720
rect 324958 443708 324964 443720
rect 325016 443708 325022 443760
rect 329098 443708 329104 443760
rect 329156 443748 329162 443760
rect 349798 443748 349804 443760
rect 329156 443720 349804 443748
rect 329156 443708 329162 443720
rect 349798 443708 349804 443720
rect 349856 443708 349862 443760
rect 217778 443640 217784 443692
rect 217836 443680 217842 443692
rect 271966 443680 271972 443692
rect 217836 443652 271972 443680
rect 217836 443640 217842 443652
rect 271966 443640 271972 443652
rect 272024 443640 272030 443692
rect 293218 443640 293224 443692
rect 293276 443680 293282 443692
rect 328914 443680 328920 443692
rect 293276 443652 328920 443680
rect 293276 443640 293282 443652
rect 328914 443640 328920 443652
rect 328972 443640 328978 443692
rect 338758 443640 338764 443692
rect 338816 443680 338822 443692
rect 358998 443680 359004 443692
rect 338816 443652 359004 443680
rect 338816 443640 338822 443652
rect 358998 443640 359004 443652
rect 359056 443640 359062 443692
rect 243722 443572 243728 443624
rect 243780 443612 243786 443624
rect 276106 443612 276112 443624
rect 243780 443584 276112 443612
rect 243780 443572 243786 443584
rect 276106 443572 276112 443584
rect 276164 443572 276170 443624
rect 251266 443504 251272 443556
rect 251324 443544 251330 443556
rect 301406 443544 301412 443556
rect 251324 443516 301412 443544
rect 251324 443504 251330 443516
rect 301406 443504 301412 443516
rect 301464 443504 301470 443556
rect 229738 443436 229744 443488
rect 229796 443476 229802 443488
rect 292850 443476 292856 443488
rect 229796 443448 292856 443476
rect 229796 443436 229802 443448
rect 292850 443436 292856 443448
rect 292908 443436 292914 443488
rect 228358 443368 228364 443420
rect 228416 443408 228422 443420
rect 294138 443408 294144 443420
rect 228416 443380 294144 443408
rect 228416 443368 228422 443380
rect 294138 443368 294144 443380
rect 294196 443368 294202 443420
rect 239214 443300 239220 443352
rect 239272 443340 239278 443352
rect 329742 443340 329748 443352
rect 239272 443312 329748 443340
rect 239272 443300 239278 443312
rect 329742 443300 329748 443312
rect 329800 443300 329806 443352
rect 196710 443232 196716 443284
rect 196768 443272 196774 443284
rect 298738 443272 298744 443284
rect 196768 443244 298744 443272
rect 196768 443232 196774 443244
rect 298738 443232 298744 443244
rect 298796 443232 298802 443284
rect 250346 443164 250352 443216
rect 250404 443204 250410 443216
rect 362494 443204 362500 443216
rect 250404 443176 362500 443204
rect 250404 443164 250410 443176
rect 362494 443164 362500 443176
rect 362552 443164 362558 443216
rect 237190 443096 237196 443148
rect 237248 443136 237254 443148
rect 245562 443136 245568 443148
rect 237248 443108 245568 443136
rect 237248 443096 237254 443108
rect 245562 443096 245568 443108
rect 245620 443096 245626 443148
rect 359642 443096 359648 443148
rect 359700 443136 359706 443148
rect 388438 443136 388444 443148
rect 359700 443108 388444 443136
rect 359700 443096 359706 443108
rect 388438 443096 388444 443108
rect 388496 443096 388502 443148
rect 276014 443028 276020 443080
rect 276072 443068 276078 443080
rect 292206 443068 292212 443080
rect 276072 443040 292212 443068
rect 276072 443028 276078 443040
rect 292206 443028 292212 443040
rect 292264 443028 292270 443080
rect 360286 443028 360292 443080
rect 360344 443068 360350 443080
rect 581086 443068 581092 443080
rect 360344 443040 581092 443068
rect 360344 443028 360350 443040
rect 581086 443028 581092 443040
rect 581144 443028 581150 443080
rect 235258 442960 235264 443012
rect 235316 443000 235322 443012
rect 242894 443000 242900 443012
rect 235316 442972 242900 443000
rect 235316 442960 235322 442972
rect 242894 442960 242900 442972
rect 242952 442960 242958 443012
rect 246390 442960 246396 443012
rect 246448 443000 246454 443012
rect 277394 443000 277400 443012
rect 246448 442972 277400 443000
rect 246448 442960 246454 442972
rect 277394 442960 277400 442972
rect 277452 442960 277458 443012
rect 280062 442960 280068 443012
rect 280120 443000 280126 443012
rect 296162 443000 296168 443012
rect 280120 442972 296168 443000
rect 280120 442960 280126 442972
rect 296162 442960 296168 442972
rect 296220 442960 296226 443012
rect 360930 442960 360936 443012
rect 360988 443000 360994 443012
rect 582374 443000 582380 443012
rect 360988 442972 582380 443000
rect 360988 442960 360994 442972
rect 582374 442960 582380 442972
rect 582432 442960 582438 443012
rect 329742 442620 329748 442672
rect 329800 442660 329806 442672
rect 580718 442660 580724 442672
rect 329800 442632 580724 442660
rect 329800 442620 329806 442632
rect 580718 442620 580724 442632
rect 580776 442620 580782 442672
rect 3510 442552 3516 442604
rect 3568 442592 3574 442604
rect 280062 442592 280068 442604
rect 3568 442564 280068 442592
rect 3568 442552 3574 442564
rect 280062 442552 280068 442564
rect 280120 442552 280126 442604
rect 300854 442552 300860 442604
rect 300912 442592 300918 442604
rect 580626 442592 580632 442604
rect 300912 442564 580632 442592
rect 300912 442552 300918 442564
rect 580626 442552 580632 442564
rect 580684 442552 580690 442604
rect 3602 442484 3608 442536
rect 3660 442524 3666 442536
rect 276014 442524 276020 442536
rect 3660 442496 276020 442524
rect 3660 442484 3666 442496
rect 276014 442484 276020 442496
rect 276072 442484 276078 442536
rect 279970 442484 279976 442536
rect 280028 442524 280034 442536
rect 580258 442524 580264 442536
rect 280028 442496 580264 442524
rect 280028 442484 280034 442496
rect 580258 442484 580264 442496
rect 580316 442484 580322 442536
rect 276106 442416 276112 442468
rect 276164 442456 276170 442468
rect 580810 442456 580816 442468
rect 276164 442428 580816 442456
rect 276164 442416 276170 442428
rect 580810 442416 580816 442428
rect 580868 442416 580874 442468
rect 251174 442348 251180 442400
rect 251232 442388 251238 442400
rect 580902 442388 580908 442400
rect 251232 442360 580908 442388
rect 251232 442348 251238 442360
rect 580902 442348 580908 442360
rect 580960 442348 580966 442400
rect 245562 442280 245568 442332
rect 245620 442320 245626 442332
rect 580534 442320 580540 442332
rect 245620 442292 580540 442320
rect 245620 442280 245626 442292
rect 580534 442280 580540 442292
rect 580592 442280 580598 442332
rect 242894 442212 242900 442264
rect 242952 442252 242958 442264
rect 580442 442252 580448 442264
rect 242952 442224 580448 442252
rect 242952 442212 242958 442224
rect 580442 442212 580448 442224
rect 580500 442212 580506 442264
rect 231210 442144 231216 442196
rect 231268 442184 231274 442196
rect 290918 442184 290924 442196
rect 231268 442156 290924 442184
rect 231268 442144 231274 442156
rect 290918 442144 290924 442156
rect 290976 442144 290982 442196
rect 206278 442076 206284 442128
rect 206336 442116 206342 442128
rect 302050 442116 302056 442128
rect 206336 442088 302056 442116
rect 206336 442076 206342 442088
rect 302050 442076 302056 442088
rect 302108 442076 302114 442128
rect 197998 442008 198004 442060
rect 198056 442048 198062 442060
rect 302694 442048 302700 442060
rect 198056 442020 302700 442048
rect 198056 442008 198062 442020
rect 302694 442008 302700 442020
rect 302752 442008 302758 442060
rect 192570 441940 192576 441992
rect 192628 441980 192634 441992
rect 306650 441980 306656 441992
rect 192628 441952 306656 441980
rect 192628 441940 192634 441952
rect 306650 441940 306656 441952
rect 306708 441940 306714 441992
rect 248966 441872 248972 441924
rect 249024 441912 249030 441924
rect 363690 441912 363696 441924
rect 249024 441884 363696 441912
rect 249024 441872 249030 441884
rect 363690 441872 363696 441884
rect 363748 441872 363754 441924
rect 140774 441804 140780 441856
rect 140832 441844 140838 441856
rect 255958 441844 255964 441856
rect 140832 441816 255964 441844
rect 140832 441804 140838 441816
rect 255958 441804 255964 441816
rect 256016 441804 256022 441856
rect 247034 441736 247040 441788
rect 247092 441776 247098 441788
rect 362310 441776 362316 441788
rect 247092 441748 362316 441776
rect 247092 441736 247098 441748
rect 362310 441736 362316 441748
rect 362368 441736 362374 441788
rect 8938 441668 8944 441720
rect 8996 441708 9002 441720
rect 296806 441708 296812 441720
rect 8996 441680 296812 441708
rect 8996 441668 9002 441680
rect 296806 441668 296812 441680
rect 296864 441668 296870 441720
rect 241146 441600 241152 441652
rect 241204 441640 241210 441652
rect 577590 441640 577596 441652
rect 241204 441612 577596 441640
rect 241204 441600 241210 441612
rect 577590 441600 577596 441612
rect 577648 441600 577654 441652
rect 289262 441436 289268 441448
rect 283944 441408 289268 441436
rect 283834 441192 283840 441244
rect 283892 441192 283898 441244
rect 242342 441124 242348 441176
rect 242400 441164 242406 441176
rect 248046 441164 248052 441176
rect 242400 441136 248052 441164
rect 242400 441124 242406 441136
rect 248046 441124 248052 441136
rect 248104 441124 248110 441176
rect 283852 441164 283880 441192
rect 283208 441136 283880 441164
rect 251266 441096 251272 441108
rect 234586 441068 251272 441096
rect 3418 440852 3424 440904
rect 3476 440892 3482 440904
rect 234586 440892 234614 441068
rect 251266 441056 251272 441068
rect 251324 441056 251330 441108
rect 251928 441068 260834 441096
rect 242342 441028 242348 441040
rect 3476 440864 234614 440892
rect 240106 441000 242348 441028
rect 3476 440852 3482 440864
rect 207658 440648 207664 440700
rect 207716 440688 207722 440700
rect 207716 440660 234614 440688
rect 207716 440648 207722 440660
rect 234586 440620 234614 440660
rect 240106 440620 240134 441000
rect 242342 440988 242348 441000
rect 242400 440988 242406 441040
rect 242710 440988 242716 441040
rect 242768 440988 242774 441040
rect 247862 440988 247868 441040
rect 247920 440988 247926 441040
rect 248046 440988 248052 441040
rect 248104 441028 248110 441040
rect 248104 441000 249794 441028
rect 248104 440988 248110 441000
rect 234586 440592 240134 440620
rect 242728 440484 242756 440988
rect 247880 440552 247908 440988
rect 249766 440960 249794 441000
rect 251928 440960 251956 441068
rect 252002 440988 252008 441040
rect 252060 440988 252066 441040
rect 249766 440932 251956 440960
rect 252020 440620 252048 440988
rect 260806 440688 260834 441068
rect 277394 440988 277400 441040
rect 277452 440988 277458 441040
rect 283098 441028 283104 441040
rect 280126 441000 283104 441028
rect 277412 440892 277440 440988
rect 280126 440892 280154 441000
rect 283098 440988 283104 441000
rect 283156 440988 283162 441040
rect 277412 440864 280154 440892
rect 283208 440688 283236 441136
rect 283834 441096 283840 441108
rect 283668 441068 283840 441096
rect 283558 440988 283564 441040
rect 283616 440988 283622 441040
rect 283576 440756 283604 440988
rect 260806 440660 283236 440688
rect 283392 440728 283604 440756
rect 283392 440620 283420 440728
rect 252020 440592 283420 440620
rect 283668 440552 283696 441068
rect 283834 441056 283840 441068
rect 283892 441056 283898 441108
rect 247880 440524 283696 440552
rect 283944 440484 283972 441408
rect 289262 441396 289268 441408
rect 289320 441396 289326 441448
rect 284570 441328 284576 441380
rect 284628 441368 284634 441380
rect 304902 441368 304908 441380
rect 284628 441340 304908 441368
rect 284628 441328 284634 441340
rect 304902 441328 304908 441340
rect 304960 441328 304966 441380
rect 284846 441260 284852 441312
rect 284904 441300 284910 441312
rect 288894 441300 288900 441312
rect 284904 441272 288900 441300
rect 284904 441260 284910 441272
rect 288894 441260 288900 441272
rect 288952 441260 288958 441312
rect 303062 441300 303068 441312
rect 293926 441272 303068 441300
rect 284018 441192 284024 441244
rect 284076 441232 284082 441244
rect 293926 441232 293954 441272
rect 303062 441260 303068 441272
rect 303120 441260 303126 441312
rect 284076 441204 293954 441232
rect 284076 441192 284082 441204
rect 298646 441192 298652 441244
rect 298704 441232 298710 441244
rect 298704 441204 309134 441232
rect 298704 441192 298710 441204
rect 288894 441124 288900 441176
rect 288952 441164 288958 441176
rect 288952 441136 298094 441164
rect 288952 441124 288958 441136
rect 284018 441056 284024 441108
rect 284076 441096 284082 441108
rect 284076 441068 294736 441096
rect 284076 441056 284082 441068
rect 284570 440988 284576 441040
rect 284628 440988 284634 441040
rect 284846 440988 284852 441040
rect 284904 440988 284910 441040
rect 289262 440988 289268 441040
rect 289320 440988 289326 441040
rect 284588 440960 284616 440988
rect 284496 440932 284616 440960
rect 284496 440756 284524 440932
rect 284864 440892 284892 440988
rect 242728 440456 283972 440484
rect 284404 440728 284524 440756
rect 284588 440864 284892 440892
rect 88978 440376 88984 440428
rect 89036 440416 89042 440428
rect 284404 440416 284432 440728
rect 89036 440388 284432 440416
rect 89036 440376 89042 440388
rect 25498 440308 25504 440360
rect 25556 440348 25562 440360
rect 284588 440348 284616 440864
rect 289280 440620 289308 440988
rect 289280 440592 294644 440620
rect 294616 440484 294644 440592
rect 294708 440552 294736 441068
rect 298066 440620 298094 441136
rect 304350 441028 304356 441040
rect 303586 441000 304356 441028
rect 303586 440756 303614 441000
rect 304350 440988 304356 441000
rect 304408 440988 304414 441040
rect 304994 440988 305000 441040
rect 305052 441028 305058 441040
rect 305052 441000 306374 441028
rect 305052 440988 305058 441000
rect 300826 440728 303614 440756
rect 300826 440688 300854 440728
rect 299446 440660 300854 440688
rect 299446 440620 299474 440660
rect 298066 440592 299474 440620
rect 306346 440620 306374 441000
rect 309106 440892 309134 441204
rect 580166 440892 580172 440904
rect 309106 440864 580172 440892
rect 580166 440852 580172 440864
rect 580224 440852 580230 440904
rect 364978 440620 364984 440632
rect 306346 440592 364984 440620
rect 364978 440580 364984 440592
rect 365036 440580 365042 440632
rect 377398 440552 377404 440564
rect 294708 440524 377404 440552
rect 377398 440512 377404 440524
rect 377456 440512 377462 440564
rect 373350 440484 373356 440496
rect 294616 440456 299474 440484
rect 25556 440320 284616 440348
rect 299446 440348 299474 440456
rect 306346 440456 373356 440484
rect 306346 440348 306374 440456
rect 373350 440444 373356 440456
rect 373408 440444 373414 440496
rect 299446 440320 306374 440348
rect 25556 440308 25562 440320
rect 97626 438132 97632 438184
rect 97684 438172 97690 438184
rect 230474 438172 230480 438184
rect 97684 438144 230480 438172
rect 97684 438132 97690 438144
rect 230474 438132 230480 438144
rect 230532 438132 230538 438184
rect 362586 431876 362592 431928
rect 362644 431916 362650 431928
rect 579798 431916 579804 431928
rect 362644 431888 579804 431916
rect 362644 431876 362650 431888
rect 579798 431876 579804 431888
rect 579856 431876 579862 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 7558 423620 7564 423632
rect 3384 423592 7564 423620
rect 3384 423580 3390 423592
rect 7558 423580 7564 423592
rect 7616 423580 7622 423632
rect 364978 419432 364984 419484
rect 365036 419472 365042 419484
rect 579982 419472 579988 419484
rect 365036 419444 579988 419472
rect 365036 419432 365042 419444
rect 579982 419432 579988 419444
rect 580040 419432 580046 419484
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 231210 411244 231216 411256
rect 3384 411216 231216 411244
rect 3384 411204 3390 411216
rect 231210 411204 231216 411216
rect 231268 411204 231274 411256
rect 362494 405628 362500 405680
rect 362552 405668 362558 405680
rect 579798 405668 579804 405680
rect 362552 405640 579804 405668
rect 362552 405628 362558 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 231118 398800 231124 398812
rect 3384 398772 231124 398800
rect 3384 398760 3390 398772
rect 231118 398760 231124 398772
rect 231176 398760 231182 398812
rect 363690 379448 363696 379500
rect 363748 379488 363754 379500
rect 580074 379488 580080 379500
rect 363748 379460 580080 379488
rect 363748 379448 363754 379460
rect 580074 379448 580080 379460
rect 580132 379448 580138 379500
rect 3694 375980 3700 376032
rect 3752 376020 3758 376032
rect 229738 376020 229744 376032
rect 3752 375992 229744 376020
rect 3752 375980 3758 375992
rect 229738 375980 229744 375992
rect 229796 375980 229802 376032
rect 154758 374892 154764 374944
rect 154816 374932 154822 374944
rect 170398 374932 170404 374944
rect 154816 374904 170404 374932
rect 154816 374892 154822 374904
rect 170398 374892 170404 374904
rect 170456 374892 170462 374944
rect 116118 374824 116124 374876
rect 116176 374864 116182 374876
rect 170950 374864 170956 374876
rect 116176 374836 170956 374864
rect 116176 374824 116182 374836
rect 170950 374824 170956 374836
rect 171008 374824 171014 374876
rect 103238 374756 103244 374808
rect 103296 374796 103302 374808
rect 225690 374796 225696 374808
rect 103296 374768 225696 374796
rect 103296 374756 103302 374768
rect 225690 374756 225696 374768
rect 225748 374756 225754 374808
rect 100662 374688 100668 374740
rect 100720 374728 100726 374740
rect 229830 374728 229836 374740
rect 100720 374700 229836 374728
rect 100720 374688 100726 374700
rect 229830 374688 229836 374700
rect 229888 374688 229894 374740
rect 147030 374620 147036 374672
rect 147088 374660 147094 374672
rect 174722 374660 174728 374672
rect 147088 374632 174728 374660
rect 147088 374620 147094 374632
rect 174722 374620 174728 374632
rect 174780 374620 174786 374672
rect 139302 374552 139308 374604
rect 139360 374592 139366 374604
rect 171778 374592 171784 374604
rect 139360 374564 171784 374592
rect 139360 374552 139366 374564
rect 171778 374552 171784 374564
rect 171836 374552 171842 374604
rect 121270 374484 121276 374536
rect 121328 374524 121334 374536
rect 170766 374524 170772 374536
rect 121328 374496 170772 374524
rect 121328 374484 121334 374496
rect 170766 374484 170772 374496
rect 170824 374484 170830 374536
rect 165522 374416 165528 374468
rect 165580 374456 165586 374468
rect 226978 374456 226984 374468
rect 165580 374428 226984 374456
rect 165580 374416 165586 374428
rect 226978 374416 226984 374428
rect 227036 374416 227042 374468
rect 167638 374348 167644 374400
rect 167696 374388 167702 374400
rect 229738 374388 229744 374400
rect 167696 374360 229744 374388
rect 167696 374348 167702 374360
rect 229738 374348 229744 374360
rect 229796 374348 229802 374400
rect 108390 374280 108396 374332
rect 108448 374320 108454 374332
rect 175918 374320 175924 374332
rect 108448 374292 175924 374320
rect 108448 374280 108454 374292
rect 175918 374280 175924 374292
rect 175976 374280 175982 374332
rect 131574 374212 131580 374264
rect 131632 374252 131638 374264
rect 228450 374252 228456 374264
rect 131632 374224 228456 374252
rect 131632 374212 131638 374224
rect 228450 374212 228456 374224
rect 228508 374212 228514 374264
rect 126422 374144 126428 374196
rect 126480 374184 126486 374196
rect 231118 374184 231124 374196
rect 126480 374156 231124 374184
rect 126480 374144 126486 374156
rect 231118 374144 231124 374156
rect 231176 374144 231182 374196
rect 162486 374008 162492 374060
rect 162544 374048 162550 374060
rect 170490 374048 170496 374060
rect 162544 374020 170496 374048
rect 162544 374008 162550 374020
rect 170490 374008 170496 374020
rect 170548 374008 170554 374060
rect 32398 373056 32404 373108
rect 32456 373096 32462 373108
rect 165062 373096 165068 373108
rect 32456 373068 165068 373096
rect 32456 373056 32462 373068
rect 165062 373056 165068 373068
rect 165120 373096 165126 373108
rect 165522 373096 165528 373108
rect 165120 373068 165528 373096
rect 165120 373056 165126 373068
rect 165522 373056 165528 373068
rect 165580 373056 165586 373108
rect 123846 372988 123852 373040
rect 123904 373028 123910 373040
rect 170582 373028 170588 373040
rect 123904 373000 170588 373028
rect 123904 372988 123910 373000
rect 170582 372988 170588 373000
rect 170640 372988 170646 373040
rect 118694 372920 118700 372972
rect 118752 372960 118758 372972
rect 174538 372960 174544 372972
rect 118752 372932 174544 372960
rect 118752 372920 118758 372932
rect 174538 372920 174544 372932
rect 174596 372920 174602 372972
rect 105814 372852 105820 372904
rect 105872 372892 105878 372904
rect 174630 372892 174636 372904
rect 105872 372864 174636 372892
rect 105872 372852 105878 372864
rect 174630 372852 174636 372864
rect 174688 372852 174694 372904
rect 149606 372784 149612 372836
rect 149664 372824 149670 372836
rect 228542 372824 228548 372836
rect 149664 372796 228548 372824
rect 149664 372784 149670 372796
rect 228542 372784 228548 372796
rect 228600 372784 228606 372836
rect 136726 372716 136732 372768
rect 136784 372756 136790 372768
rect 224218 372756 224224 372768
rect 136784 372728 224224 372756
rect 136784 372716 136790 372728
rect 224218 372716 224224 372728
rect 224276 372716 224282 372768
rect 110966 372648 110972 372700
rect 111024 372688 111030 372700
rect 228634 372688 228640 372700
rect 111024 372660 228640 372688
rect 111024 372648 111030 372660
rect 228634 372648 228640 372660
rect 228692 372648 228698 372700
rect 157334 372580 157340 372632
rect 157392 372620 157398 372632
rect 173158 372620 173164 372632
rect 157392 372592 173164 372620
rect 157392 372580 157398 372592
rect 173158 372580 173164 372592
rect 173216 372580 173222 372632
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 100018 372552 100024 372564
rect 3384 372524 100024 372552
rect 3384 372512 3390 372524
rect 100018 372512 100024 372524
rect 100076 372512 100082 372564
rect 103486 371844 161474 371872
rect 97810 371696 97816 371748
rect 97868 371736 97874 371748
rect 103486 371736 103514 371844
rect 97868 371708 103514 371736
rect 109006 371776 118694 371804
rect 97868 371696 97874 371708
rect 97718 371628 97724 371680
rect 97776 371668 97782 371680
rect 109006 371668 109034 371776
rect 113450 371696 113456 371748
rect 113508 371736 113514 371748
rect 115750 371736 115756 371748
rect 113508 371708 115756 371736
rect 113508 371696 113514 371708
rect 115750 371696 115756 371708
rect 115808 371696 115814 371748
rect 118666 371668 118694 371776
rect 134058 371764 134064 371816
rect 134116 371804 134122 371816
rect 134116 371776 157334 371804
rect 134116 371764 134122 371776
rect 133828 371736 133834 371748
rect 121426 371708 133834 371736
rect 121426 371668 121454 371708
rect 133828 371696 133834 371708
rect 133886 371696 133892 371748
rect 143166 371696 143172 371748
rect 143224 371736 143230 371748
rect 144362 371736 144368 371748
rect 143224 371708 144368 371736
rect 143224 371696 143230 371708
rect 144362 371696 144368 371708
rect 144420 371696 144426 371748
rect 144886 371708 153148 371736
rect 97776 371640 109034 371668
rect 111076 371640 115934 371668
rect 118666 371640 121454 371668
rect 128326 371640 129412 371668
rect 97776 371628 97782 371640
rect 99834 371560 99840 371612
rect 99892 371600 99898 371612
rect 111076 371600 111104 371640
rect 113450 371600 113456 371612
rect 99892 371572 111104 371600
rect 113146 371572 113456 371600
rect 99892 371560 99898 371572
rect 97902 371492 97908 371544
rect 97960 371532 97966 371544
rect 97960 371504 103514 371532
rect 97960 371492 97966 371504
rect 103486 371464 103514 371504
rect 103486 371436 106274 371464
rect 106246 371260 106274 371436
rect 113146 371260 113174 371572
rect 113450 371560 113456 371572
rect 113508 371560 113514 371612
rect 113818 371560 113824 371612
rect 113876 371560 113882 371612
rect 115750 371560 115756 371612
rect 115808 371560 115814 371612
rect 106246 371232 113174 371260
rect 113836 371056 113864 371560
rect 115768 371464 115796 371560
rect 115906 371532 115934 371640
rect 128326 371600 128354 371640
rect 118666 371572 128354 371600
rect 118666 371532 118694 371572
rect 129182 371560 129188 371612
rect 129240 371560 129246 371612
rect 129384 371600 129412 371640
rect 135162 371628 135168 371680
rect 135220 371668 135226 371680
rect 144886 371668 144914 371708
rect 135220 371640 144914 371668
rect 135220 371628 135226 371640
rect 145006 371628 145012 371680
rect 145064 371668 145070 371680
rect 145064 371640 145788 371668
rect 145064 371628 145070 371640
rect 133828 371600 133834 371612
rect 129384 371572 133834 371600
rect 133828 371560 133834 371572
rect 133886 371560 133892 371612
rect 143166 371600 143172 371612
rect 133984 371572 143172 371600
rect 115906 371504 118694 371532
rect 129200 371464 129228 371560
rect 133984 371532 134012 371572
rect 143166 371560 143172 371572
rect 143224 371560 143230 371612
rect 143258 371560 143264 371612
rect 143316 371560 143322 371612
rect 144362 371560 144368 371612
rect 144420 371560 144426 371612
rect 144730 371560 144736 371612
rect 144788 371600 144794 371612
rect 144914 371600 144920 371612
rect 144788 371572 144920 371600
rect 144788 371560 144794 371572
rect 144914 371560 144920 371572
rect 144972 371560 144978 371612
rect 143276 371532 143304 371560
rect 132466 371504 134012 371532
rect 142126 371504 143304 371532
rect 144380 371532 144408 371560
rect 144380 371504 144868 371532
rect 132466 371464 132494 371504
rect 142126 371464 142154 371504
rect 115768 371436 122834 371464
rect 129200 371436 132494 371464
rect 140746 371436 142154 371464
rect 122806 371124 122834 371436
rect 140746 371396 140774 371436
rect 135226 371368 136634 371396
rect 135226 371192 135254 371368
rect 136606 371328 136634 371368
rect 137986 371368 140774 371396
rect 137986 371328 138014 371368
rect 144840 371328 144868 371504
rect 145760 371396 145788 371640
rect 153010 371628 153016 371680
rect 153068 371628 153074 371680
rect 152550 371560 152556 371612
rect 152608 371600 152614 371612
rect 152608 371572 152688 371600
rect 152608 371560 152614 371572
rect 152660 371464 152688 371572
rect 153028 371532 153056 371628
rect 153120 371600 153148 371708
rect 157306 371668 157334 371776
rect 161446 371736 161474 371844
rect 173250 371736 173256 371748
rect 161446 371708 173256 371736
rect 173250 371696 173256 371708
rect 173308 371696 173314 371748
rect 229922 371668 229928 371680
rect 157306 371640 229928 371668
rect 229922 371628 229928 371640
rect 229980 371628 229986 371680
rect 231210 371600 231216 371612
rect 153120 371572 231216 371600
rect 231210 371560 231216 371572
rect 231268 371560 231274 371612
rect 231394 371532 231400 371544
rect 153028 371504 231400 371532
rect 231394 371492 231400 371504
rect 231452 371492 231458 371544
rect 231302 371464 231308 371476
rect 152660 371436 231308 371464
rect 231302 371424 231308 371436
rect 231360 371424 231366 371476
rect 230014 371396 230020 371408
rect 145760 371368 230020 371396
rect 230014 371356 230020 371368
rect 230072 371356 230078 371408
rect 230106 371328 230112 371340
rect 136606 371300 138014 371328
rect 142126 371300 143534 371328
rect 144840 371300 230112 371328
rect 142126 371260 142154 371300
rect 140746 371232 142154 371260
rect 140746 371192 140774 371232
rect 124186 371164 125594 371192
rect 124186 371124 124214 371164
rect 122806 371096 124214 371124
rect 125566 371124 125594 371164
rect 129706 371164 132494 371192
rect 129706 371124 129734 371164
rect 125566 371096 129734 371124
rect 132466 371124 132494 371164
rect 133846 371164 135254 371192
rect 137986 371164 140774 371192
rect 133846 371124 133874 371164
rect 137986 371124 138014 371164
rect 132466 371096 133874 371124
rect 136606 371096 138014 371124
rect 143506 371124 143534 371300
rect 230106 371288 230112 371300
rect 230164 371288 230170 371340
rect 231486 371260 231492 371272
rect 144886 371232 231492 371260
rect 144886 371124 144914 371232
rect 231486 371220 231492 371232
rect 231544 371220 231550 371272
rect 143506 371096 144914 371124
rect 136606 371056 136634 371096
rect 113836 371028 124214 371056
rect 124186 370988 124214 371028
rect 128326 371028 129734 371056
rect 128326 370988 128354 371028
rect 124186 370960 128354 370988
rect 129706 370988 129734 371028
rect 131086 371028 133874 371056
rect 131086 370988 131114 371028
rect 129706 370960 131114 370988
rect 133846 370988 133874 371028
rect 135226 371028 136634 371056
rect 135226 370988 135254 371028
rect 133846 370960 135254 370988
rect 172330 368500 172336 368552
rect 172388 368540 172394 368552
rect 227070 368540 227076 368552
rect 172388 368512 227076 368540
rect 172388 368500 172394 368512
rect 227070 368500 227076 368512
rect 227128 368500 227134 368552
rect 169938 367888 169944 367940
rect 169996 367928 170002 367940
rect 170674 367928 170680 367940
rect 169996 367900 170680 367928
rect 169996 367888 170002 367900
rect 170674 367888 170680 367900
rect 170732 367888 170738 367940
rect 172422 365712 172428 365764
rect 172480 365752 172486 365764
rect 231578 365752 231584 365764
rect 172480 365724 231584 365752
rect 172480 365712 172486 365724
rect 231578 365712 231584 365724
rect 231636 365712 231642 365764
rect 363598 365644 363604 365696
rect 363656 365684 363662 365696
rect 580074 365684 580080 365696
rect 363656 365656 580080 365684
rect 363656 365644 363662 365656
rect 580074 365644 580080 365656
rect 580132 365644 580138 365696
rect 171686 357416 171692 357468
rect 171744 357456 171750 357468
rect 228726 357456 228732 357468
rect 171744 357428 228732 357456
rect 171744 357416 171750 357428
rect 228726 357416 228732 357428
rect 228784 357416 228790 357468
rect 172422 354696 172428 354748
rect 172480 354736 172486 354748
rect 230198 354736 230204 354748
rect 172480 354708 230204 354736
rect 172480 354696 172486 354708
rect 230198 354696 230204 354708
rect 230256 354696 230262 354748
rect 362402 353200 362408 353252
rect 362460 353240 362466 353252
rect 579982 353240 579988 353252
rect 362460 353212 579988 353240
rect 362460 353200 362466 353212
rect 579982 353200 579988 353212
rect 580040 353200 580046 353252
rect 172422 351908 172428 351960
rect 172480 351948 172486 351960
rect 227162 351948 227168 351960
rect 172480 351920 227168 351948
rect 172480 351908 172486 351920
rect 227162 351908 227168 351920
rect 227220 351908 227226 351960
rect 171686 350480 171692 350532
rect 171744 350520 171750 350532
rect 171870 350520 171876 350532
rect 171744 350492 171876 350520
rect 171744 350480 171750 350492
rect 171870 350480 171876 350492
rect 171928 350480 171934 350532
rect 171134 349120 171140 349172
rect 171192 349160 171198 349172
rect 171870 349160 171876 349172
rect 171192 349132 171876 349160
rect 171192 349120 171198 349132
rect 171870 349120 171876 349132
rect 171928 349160 171934 349172
rect 192478 349160 192484 349172
rect 171928 349132 192484 349160
rect 171928 349120 171934 349132
rect 192478 349120 192484 349132
rect 192536 349120 192542 349172
rect 172422 346400 172428 346452
rect 172480 346440 172486 346452
rect 220078 346440 220084 346452
rect 172480 346412 220084 346440
rect 172480 346400 172486 346412
rect 220078 346400 220084 346412
rect 220136 346400 220142 346452
rect 172422 342252 172428 342304
rect 172480 342292 172486 342304
rect 231670 342292 231676 342304
rect 172480 342264 231676 342292
rect 172480 342252 172486 342264
rect 231670 342252 231676 342264
rect 231728 342252 231734 342304
rect 172422 336744 172428 336796
rect 172480 336784 172486 336796
rect 230290 336784 230296 336796
rect 172480 336756 230296 336784
rect 172480 336744 172486 336756
rect 230290 336744 230296 336756
rect 230348 336744 230354 336796
rect 172422 333956 172428 334008
rect 172480 333996 172486 334008
rect 228818 333996 228824 334008
rect 172480 333968 228824 333996
rect 172480 333956 172486 333968
rect 228818 333956 228824 333968
rect 228876 333956 228882 334008
rect 172422 331236 172428 331288
rect 172480 331276 172486 331288
rect 230382 331276 230388 331288
rect 172480 331248 230388 331276
rect 172480 331236 172486 331248
rect 230382 331236 230388 331248
rect 230440 331236 230446 331288
rect 172422 328448 172428 328500
rect 172480 328488 172486 328500
rect 225782 328488 225788 328500
rect 172480 328460 225788 328488
rect 172480 328448 172486 328460
rect 225782 328448 225788 328460
rect 225840 328448 225846 328500
rect 171410 325660 171416 325712
rect 171468 325700 171474 325712
rect 232222 325700 232228 325712
rect 171468 325672 232228 325700
rect 171468 325660 171474 325672
rect 232222 325660 232228 325672
rect 232280 325660 232286 325712
rect 362310 325592 362316 325644
rect 362368 325632 362374 325644
rect 580074 325632 580080 325644
rect 362368 325604 580080 325632
rect 362368 325592 362374 325604
rect 580074 325592 580080 325604
rect 580132 325592 580138 325644
rect 172422 320152 172428 320204
rect 172480 320192 172486 320204
rect 231762 320192 231768 320204
rect 172480 320164 231768 320192
rect 172480 320152 172486 320164
rect 231762 320152 231768 320164
rect 231820 320152 231826 320204
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 95878 320124 95884 320136
rect 3384 320096 95884 320124
rect 3384 320084 3390 320096
rect 95878 320084 95884 320096
rect 95936 320084 95942 320136
rect 172422 317432 172428 317484
rect 172480 317472 172486 317484
rect 231854 317472 231860 317484
rect 172480 317444 231860 317472
rect 172480 317432 172486 317444
rect 231854 317432 231860 317444
rect 231912 317432 231918 317484
rect 172422 314644 172428 314696
rect 172480 314684 172486 314696
rect 231946 314684 231952 314696
rect 172480 314656 231952 314684
rect 172480 314644 172486 314656
rect 231946 314644 231952 314656
rect 232004 314644 232010 314696
rect 377398 313216 377404 313268
rect 377456 313256 377462 313268
rect 579982 313256 579988 313268
rect 377456 313228 579988 313256
rect 377456 313216 377462 313228
rect 579982 313216 579988 313228
rect 580040 313216 580046 313268
rect 230934 312944 230940 312996
rect 230992 312984 230998 312996
rect 231302 312984 231308 312996
rect 230992 312956 231308 312984
rect 230992 312944 230998 312956
rect 231302 312944 231308 312956
rect 231360 312944 231366 312996
rect 231394 312672 231400 312724
rect 231452 312712 231458 312724
rect 231670 312712 231676 312724
rect 231452 312684 231676 312712
rect 231452 312672 231458 312684
rect 231670 312672 231676 312684
rect 231728 312672 231734 312724
rect 172422 311856 172428 311908
rect 172480 311896 172486 311908
rect 231854 311896 231860 311908
rect 172480 311868 231860 311896
rect 172480 311856 172486 311868
rect 231854 311856 231860 311868
rect 231912 311856 231918 311908
rect 231762 311788 231768 311840
rect 231820 311828 231826 311840
rect 232038 311828 232044 311840
rect 231820 311800 232044 311828
rect 231820 311788 231826 311800
rect 232038 311788 232044 311800
rect 232096 311788 232102 311840
rect 172146 311312 172152 311364
rect 172204 311352 172210 311364
rect 231026 311352 231032 311364
rect 172204 311324 231032 311352
rect 172204 311312 172210 311324
rect 231026 311312 231032 311324
rect 231084 311312 231090 311364
rect 171778 311244 171784 311296
rect 171836 311284 171842 311296
rect 232130 311284 232136 311296
rect 171836 311256 232136 311284
rect 171836 311244 171842 311256
rect 232130 311244 232136 311256
rect 232188 311244 232194 311296
rect 171962 311176 171968 311228
rect 172020 311216 172026 311228
rect 231762 311216 231768 311228
rect 172020 311188 231768 311216
rect 172020 311176 172026 311188
rect 231762 311176 231768 311188
rect 231820 311176 231826 311228
rect 192478 311108 192484 311160
rect 192536 311148 192542 311160
rect 232222 311148 232228 311160
rect 192536 311120 232228 311148
rect 192536 311108 192542 311120
rect 232222 311108 232228 311120
rect 232280 311108 232286 311160
rect 219406 310712 232084 310740
rect 171870 310564 171876 310616
rect 171928 310604 171934 310616
rect 219406 310604 219434 310712
rect 228818 310632 228824 310684
rect 228876 310672 228882 310684
rect 228876 310644 231992 310672
rect 228876 310632 228882 310644
rect 171928 310576 219434 310604
rect 171928 310564 171934 310576
rect 226978 310496 226984 310548
rect 227036 310536 227042 310548
rect 231964 310536 231992 310644
rect 232056 310604 232084 310712
rect 233142 310604 233148 310616
rect 232056 310576 233148 310604
rect 233142 310564 233148 310576
rect 233200 310564 233206 310616
rect 227036 310508 231808 310536
rect 231964 310508 232084 310536
rect 227036 310496 227042 310508
rect 231780 310400 231808 310508
rect 232056 310468 232084 310508
rect 232130 310496 232136 310548
rect 232188 310536 232194 310548
rect 232774 310536 232780 310548
rect 232188 310508 232780 310536
rect 232188 310496 232194 310508
rect 232774 310496 232780 310508
rect 232832 310496 232838 310548
rect 233694 310536 233700 310548
rect 232884 310508 233700 310536
rect 232884 310468 232912 310508
rect 233694 310496 233700 310508
rect 233752 310496 233758 310548
rect 255406 310496 255412 310548
rect 255464 310536 255470 310548
rect 255590 310536 255596 310548
rect 255464 310508 255596 310536
rect 255464 310496 255470 310508
rect 255590 310496 255596 310508
rect 255648 310496 255654 310548
rect 273530 310496 273536 310548
rect 273588 310536 273594 310548
rect 273714 310536 273720 310548
rect 273588 310508 273720 310536
rect 273588 310496 273594 310508
rect 273714 310496 273720 310508
rect 273772 310496 273778 310548
rect 232056 310440 232912 310468
rect 232590 310400 232596 310412
rect 231780 310372 232596 310400
rect 232590 310360 232596 310372
rect 232648 310360 232654 310412
rect 231946 310292 231952 310344
rect 232004 310332 232010 310344
rect 235534 310332 235540 310344
rect 232004 310304 235540 310332
rect 232004 310292 232010 310304
rect 235534 310292 235540 310304
rect 235592 310292 235598 310344
rect 231854 310224 231860 310276
rect 231912 310264 231918 310276
rect 236270 310264 236276 310276
rect 231912 310236 236276 310264
rect 231912 310224 231918 310236
rect 236270 310224 236276 310236
rect 236328 310224 236334 310276
rect 230290 310156 230296 310208
rect 230348 310196 230354 310208
rect 238938 310196 238944 310208
rect 230348 310168 238944 310196
rect 230348 310156 230354 310168
rect 238938 310156 238944 310168
rect 238996 310156 239002 310208
rect 235902 310128 235908 310140
rect 219406 310100 235908 310128
rect 172422 310020 172428 310072
rect 172480 310060 172486 310072
rect 219406 310060 219434 310100
rect 235902 310088 235908 310100
rect 235960 310088 235966 310140
rect 172480 310032 219434 310060
rect 172480 310020 172486 310032
rect 231026 310020 231032 310072
rect 231084 310060 231090 310072
rect 231946 310060 231952 310072
rect 231084 310032 231952 310060
rect 231084 310020 231090 310032
rect 231946 310020 231952 310032
rect 232004 310020 232010 310072
rect 172238 309952 172244 310004
rect 172296 309992 172302 310004
rect 239490 309992 239496 310004
rect 172296 309964 239496 309992
rect 172296 309952 172302 309964
rect 239490 309952 239496 309964
rect 239548 309952 239554 310004
rect 232958 309884 232964 309936
rect 233016 309924 233022 309936
rect 244458 309924 244464 309936
rect 233016 309896 244464 309924
rect 233016 309884 233022 309896
rect 244458 309884 244464 309896
rect 244516 309884 244522 309936
rect 230198 309816 230204 309868
rect 230256 309856 230262 309868
rect 238754 309856 238760 309868
rect 230256 309828 238760 309856
rect 230256 309816 230262 309828
rect 238754 309816 238760 309828
rect 238812 309816 238818 309868
rect 230382 309612 230388 309664
rect 230440 309652 230446 309664
rect 241790 309652 241796 309664
rect 230440 309624 241796 309652
rect 230440 309612 230446 309624
rect 241790 309612 241796 309624
rect 241848 309612 241854 309664
rect 228726 309476 228732 309528
rect 228784 309516 228790 309528
rect 242986 309516 242992 309528
rect 228784 309488 242992 309516
rect 228784 309476 228790 309488
rect 242986 309476 242992 309488
rect 243044 309476 243050 309528
rect 231578 309408 231584 309460
rect 231636 309448 231642 309460
rect 247494 309448 247500 309460
rect 231636 309420 247500 309448
rect 231636 309408 231642 309420
rect 247494 309408 247500 309420
rect 247552 309408 247558 309460
rect 315942 309408 315948 309460
rect 316000 309448 316006 309460
rect 316402 309448 316408 309460
rect 316000 309420 316408 309448
rect 316000 309408 316006 309420
rect 316402 309408 316408 309420
rect 316460 309408 316466 309460
rect 232038 309340 232044 309392
rect 232096 309380 232102 309392
rect 249610 309380 249616 309392
rect 232096 309352 249616 309380
rect 232096 309340 232102 309352
rect 249610 309340 249616 309352
rect 249668 309340 249674 309392
rect 231670 309272 231676 309324
rect 231728 309312 231734 309324
rect 236546 309312 236552 309324
rect 231728 309284 236552 309312
rect 231728 309272 231734 309284
rect 236546 309272 236552 309284
rect 236604 309272 236610 309324
rect 236656 309284 241514 309312
rect 231394 309204 231400 309256
rect 231452 309244 231458 309256
rect 236656 309244 236684 309284
rect 231452 309216 236684 309244
rect 241486 309244 241514 309284
rect 252830 309244 252836 309256
rect 241486 309216 252836 309244
rect 231452 309204 231458 309216
rect 252830 309204 252836 309216
rect 252888 309204 252894 309256
rect 170674 309136 170680 309188
rect 170732 309176 170738 309188
rect 234154 309176 234160 309188
rect 170732 309148 234160 309176
rect 170732 309136 170738 309148
rect 234154 309136 234160 309148
rect 234212 309136 234218 309188
rect 236546 309136 236552 309188
rect 236604 309176 236610 309188
rect 249794 309176 249800 309188
rect 236604 309148 249800 309176
rect 236604 309136 236610 309148
rect 249794 309136 249800 309148
rect 249852 309136 249858 309188
rect 354214 309136 354220 309188
rect 354272 309176 354278 309188
rect 354272 309148 355640 309176
rect 354272 309136 354278 309148
rect 229922 309068 229928 309120
rect 229980 309108 229986 309120
rect 233602 309108 233608 309120
rect 229980 309080 233608 309108
rect 229980 309068 229986 309080
rect 233602 309068 233608 309080
rect 233660 309068 233666 309120
rect 235810 309068 235816 309120
rect 235868 309108 235874 309120
rect 238570 309108 238576 309120
rect 235868 309080 238576 309108
rect 235868 309068 235874 309080
rect 238570 309068 238576 309080
rect 238628 309068 238634 309120
rect 347682 309068 347688 309120
rect 347740 309108 347746 309120
rect 347740 309080 355548 309108
rect 347740 309068 347746 309080
rect 231486 309000 231492 309052
rect 231544 309040 231550 309052
rect 235350 309040 235356 309052
rect 231544 309012 235356 309040
rect 231544 309000 231550 309012
rect 235350 309000 235356 309012
rect 235408 309000 235414 309052
rect 348694 309000 348700 309052
rect 348752 309040 348758 309052
rect 348752 309012 355364 309040
rect 348752 309000 348758 309012
rect 231210 308932 231216 308984
rect 231268 308972 231274 308984
rect 235718 308972 235724 308984
rect 231268 308944 235724 308972
rect 231268 308932 231274 308944
rect 235718 308932 235724 308944
rect 235776 308932 235782 308984
rect 262398 308972 262404 308984
rect 258184 308944 262404 308972
rect 230014 308864 230020 308916
rect 230072 308904 230078 308916
rect 238202 308904 238208 308916
rect 230072 308876 238208 308904
rect 230072 308864 230078 308876
rect 238202 308864 238208 308876
rect 238260 308864 238266 308916
rect 241606 308904 241612 308916
rect 238312 308876 241612 308904
rect 231854 308796 231860 308848
rect 231912 308836 231918 308848
rect 238312 308836 238340 308876
rect 241606 308864 241612 308876
rect 241664 308864 241670 308916
rect 245838 308836 245844 308848
rect 231912 308808 238340 308836
rect 239416 308808 245844 308836
rect 231912 308796 231918 308808
rect 231946 308728 231952 308780
rect 232004 308768 232010 308780
rect 239416 308768 239444 308808
rect 245838 308796 245844 308808
rect 245896 308796 245902 308848
rect 248138 308768 248144 308780
rect 232004 308740 239444 308768
rect 244246 308740 248144 308768
rect 232004 308728 232010 308740
rect 173158 308660 173164 308712
rect 173216 308700 173222 308712
rect 244246 308700 244274 308740
rect 248138 308728 248144 308740
rect 248196 308728 248202 308780
rect 173216 308672 244274 308700
rect 173216 308660 173222 308672
rect 247954 308660 247960 308712
rect 248012 308700 248018 308712
rect 254394 308700 254400 308712
rect 248012 308672 254400 308700
rect 248012 308660 248018 308672
rect 254394 308660 254400 308672
rect 254452 308660 254458 308712
rect 230934 308592 230940 308644
rect 230992 308632 230998 308644
rect 240318 308632 240324 308644
rect 230992 308604 240324 308632
rect 230992 308592 230998 308604
rect 240318 308592 240324 308604
rect 240376 308592 240382 308644
rect 253198 308592 253204 308644
rect 253256 308632 253262 308644
rect 258184 308632 258212 308944
rect 262398 308932 262404 308944
rect 262456 308932 262462 308984
rect 314838 308932 314844 308984
rect 314896 308972 314902 308984
rect 315022 308972 315028 308984
rect 314896 308944 315028 308972
rect 314896 308932 314902 308944
rect 315022 308932 315028 308944
rect 315080 308932 315086 308984
rect 326706 308932 326712 308984
rect 326764 308972 326770 308984
rect 338850 308972 338856 308984
rect 326764 308944 338856 308972
rect 326764 308932 326770 308944
rect 338850 308932 338856 308944
rect 338908 308932 338914 308984
rect 348510 308932 348516 308984
rect 348568 308972 348574 308984
rect 352098 308972 352104 308984
rect 348568 308944 352104 308972
rect 348568 308932 348574 308944
rect 352098 308932 352104 308944
rect 352156 308932 352162 308984
rect 355336 308972 355364 309012
rect 355520 308972 355548 309080
rect 355612 309040 355640 309148
rect 355686 309068 355692 309120
rect 355744 309108 355750 309120
rect 367738 309108 367744 309120
rect 355744 309080 367744 309108
rect 355744 309068 355750 309080
rect 367738 309068 367744 309080
rect 367796 309068 367802 309120
rect 366266 309040 366272 309052
rect 355612 309012 366272 309040
rect 366266 309000 366272 309012
rect 366324 309000 366330 309052
rect 367646 308972 367652 308984
rect 355336 308944 355456 308972
rect 355520 308944 367652 308972
rect 266998 308904 267004 308916
rect 253256 308604 258212 308632
rect 259104 308876 267004 308904
rect 253256 308592 253262 308604
rect 170582 308524 170588 308576
rect 170640 308564 170646 308576
rect 242342 308564 242348 308576
rect 170640 308536 242348 308564
rect 170640 308524 170646 308536
rect 242342 308524 242348 308536
rect 242400 308524 242406 308576
rect 250438 308524 250444 308576
rect 250496 308564 250502 308576
rect 258994 308564 259000 308576
rect 250496 308536 259000 308564
rect 250496 308524 250502 308536
rect 258994 308524 259000 308536
rect 259052 308524 259058 308576
rect 253290 308456 253296 308508
rect 253348 308496 253354 308508
rect 259104 308496 259132 308876
rect 266998 308864 267004 308876
rect 267056 308864 267062 308916
rect 310330 308864 310336 308916
rect 310388 308904 310394 308916
rect 310388 308876 316034 308904
rect 310388 308864 310394 308876
rect 260374 308796 260380 308848
rect 260432 308836 260438 308848
rect 268746 308836 268752 308848
rect 260432 308808 268752 308836
rect 260432 308796 260438 308808
rect 268746 308796 268752 308808
rect 268804 308796 268810 308848
rect 314654 308796 314660 308848
rect 314712 308836 314718 308848
rect 315390 308836 315396 308848
rect 314712 308808 315396 308836
rect 314712 308796 314718 308808
rect 315390 308796 315396 308808
rect 315448 308796 315454 308848
rect 316006 308836 316034 308876
rect 317414 308864 317420 308916
rect 317472 308904 317478 308916
rect 317966 308904 317972 308916
rect 317472 308876 317972 308904
rect 317472 308864 317478 308876
rect 317966 308864 317972 308876
rect 318024 308864 318030 308916
rect 319070 308864 319076 308916
rect 319128 308904 319134 308916
rect 319346 308904 319352 308916
rect 319128 308876 319352 308904
rect 319128 308864 319134 308876
rect 319346 308864 319352 308876
rect 319404 308864 319410 308916
rect 355428 308904 355456 308944
rect 367646 308932 367652 308944
rect 367704 308932 367710 308984
rect 371418 308904 371424 308916
rect 350506 308876 355364 308904
rect 355428 308876 371424 308904
rect 350506 308836 350534 308876
rect 316006 308808 350534 308836
rect 303798 308728 303804 308780
rect 303856 308768 303862 308780
rect 355226 308768 355232 308780
rect 303856 308740 355232 308768
rect 303856 308728 303862 308740
rect 355226 308728 355232 308740
rect 355284 308728 355290 308780
rect 355336 308768 355364 308876
rect 371418 308864 371424 308876
rect 371476 308864 371482 308916
rect 356514 308796 356520 308848
rect 356572 308836 356578 308848
rect 356572 308808 364334 308836
rect 356572 308796 356578 308808
rect 357158 308768 357164 308780
rect 355336 308740 357164 308768
rect 357158 308728 357164 308740
rect 357216 308728 357222 308780
rect 304534 308660 304540 308712
rect 304592 308700 304598 308712
rect 355502 308700 355508 308712
rect 304592 308672 355508 308700
rect 304592 308660 304598 308672
rect 355502 308660 355508 308672
rect 355560 308660 355566 308712
rect 364306 308700 364334 308808
rect 367370 308700 367376 308712
rect 364306 308672 367376 308700
rect 367370 308660 367376 308672
rect 367428 308660 367434 308712
rect 260098 308592 260104 308644
rect 260156 308632 260162 308644
rect 271598 308632 271604 308644
rect 260156 308604 271604 308632
rect 260156 308592 260162 308604
rect 271598 308592 271604 308604
rect 271656 308592 271662 308644
rect 302510 308592 302516 308644
rect 302568 308632 302574 308644
rect 355686 308632 355692 308644
rect 302568 308604 355692 308632
rect 302568 308592 302574 308604
rect 355686 308592 355692 308604
rect 355744 308592 355750 308644
rect 356054 308592 356060 308644
rect 356112 308632 356118 308644
rect 367554 308632 367560 308644
rect 356112 308604 367560 308632
rect 356112 308592 356118 308604
rect 367554 308592 367560 308604
rect 367612 308592 367618 308644
rect 271230 308524 271236 308576
rect 271288 308564 271294 308576
rect 273438 308564 273444 308576
rect 271288 308536 273444 308564
rect 271288 308524 271294 308536
rect 273438 308524 273444 308536
rect 273496 308524 273502 308576
rect 302326 308524 302332 308576
rect 302384 308564 302390 308576
rect 355594 308564 355600 308576
rect 302384 308536 355600 308564
rect 302384 308524 302390 308536
rect 355594 308524 355600 308536
rect 355652 308524 355658 308576
rect 357250 308524 357256 308576
rect 357308 308564 357314 308576
rect 368566 308564 368572 308576
rect 357308 308536 368572 308564
rect 357308 308524 357314 308536
rect 368566 308524 368572 308536
rect 368624 308524 368630 308576
rect 253348 308468 259132 308496
rect 253348 308456 253354 308468
rect 266998 308456 267004 308508
rect 267056 308496 267062 308508
rect 281258 308496 281264 308508
rect 267056 308468 281264 308496
rect 267056 308456 267062 308468
rect 281258 308456 281264 308468
rect 281316 308456 281322 308508
rect 301498 308456 301504 308508
rect 301556 308496 301562 308508
rect 355410 308496 355416 308508
rect 301556 308468 355416 308496
rect 301556 308456 301562 308468
rect 355410 308456 355416 308468
rect 355468 308456 355474 308508
rect 360194 308456 360200 308508
rect 360252 308496 360258 308508
rect 360838 308496 360844 308508
rect 360252 308468 360844 308496
rect 360252 308456 360258 308468
rect 360838 308456 360844 308468
rect 360896 308456 360902 308508
rect 370038 308496 370044 308508
rect 364306 308468 370044 308496
rect 224218 308388 224224 308440
rect 224276 308428 224282 308440
rect 237006 308428 237012 308440
rect 224276 308400 237012 308428
rect 224276 308388 224282 308400
rect 237006 308388 237012 308400
rect 237064 308388 237070 308440
rect 272702 308428 272708 308440
rect 253906 308400 272708 308428
rect 174538 308320 174544 308372
rect 174596 308360 174602 308372
rect 250346 308360 250352 308372
rect 174596 308332 250352 308360
rect 174596 308320 174602 308332
rect 250346 308320 250352 308332
rect 250404 308320 250410 308372
rect 228542 308252 228548 308304
rect 228600 308292 228606 308304
rect 228600 308264 244274 308292
rect 228600 308252 228606 308264
rect 230106 308184 230112 308236
rect 230164 308224 230170 308236
rect 242158 308224 242164 308236
rect 230164 308196 242164 308224
rect 230164 308184 230170 308196
rect 242158 308184 242164 308196
rect 242216 308184 242222 308236
rect 244246 308224 244274 308264
rect 246758 308224 246764 308236
rect 244246 308196 246764 308224
rect 246758 308184 246764 308196
rect 246816 308184 246822 308236
rect 246298 308116 246304 308168
rect 246356 308156 246362 308168
rect 253474 308156 253480 308168
rect 246356 308128 253480 308156
rect 246356 308116 246362 308128
rect 253474 308116 253480 308128
rect 253532 308116 253538 308168
rect 252186 308048 252192 308100
rect 252244 308088 252250 308100
rect 253906 308088 253934 308400
rect 272702 308388 272708 308400
rect 272760 308388 272766 308440
rect 301314 308388 301320 308440
rect 301372 308428 301378 308440
rect 356514 308428 356520 308440
rect 301372 308400 356520 308428
rect 301372 308388 301378 308400
rect 356514 308388 356520 308400
rect 356572 308388 356578 308440
rect 356882 308388 356888 308440
rect 356940 308428 356946 308440
rect 364306 308428 364334 308468
rect 370038 308456 370044 308468
rect 370096 308456 370102 308508
rect 356940 308400 364334 308428
rect 356940 308388 356946 308400
rect 312262 308320 312268 308372
rect 312320 308360 312326 308372
rect 312998 308360 313004 308372
rect 312320 308332 313004 308360
rect 312320 308320 312326 308332
rect 312998 308320 313004 308332
rect 313056 308320 313062 308372
rect 313918 308360 313924 308372
rect 313384 308332 313924 308360
rect 313384 308304 313412 308332
rect 313918 308320 313924 308332
rect 313976 308320 313982 308372
rect 314930 308320 314936 308372
rect 314988 308360 314994 308372
rect 315850 308360 315856 308372
rect 314988 308332 315856 308360
rect 314988 308320 314994 308332
rect 315850 308320 315856 308332
rect 315908 308320 315914 308372
rect 316126 308320 316132 308372
rect 316184 308360 316190 308372
rect 316954 308360 316960 308372
rect 316184 308332 316960 308360
rect 316184 308320 316190 308332
rect 316954 308320 316960 308332
rect 317012 308320 317018 308372
rect 317598 308320 317604 308372
rect 317656 308360 317662 308372
rect 318334 308360 318340 308372
rect 317656 308332 318340 308360
rect 317656 308320 317662 308332
rect 318334 308320 318340 308332
rect 318392 308320 318398 308372
rect 319162 308320 319168 308372
rect 319220 308360 319226 308372
rect 319806 308360 319812 308372
rect 319220 308332 319812 308360
rect 319220 308320 319226 308332
rect 319806 308320 319812 308332
rect 319864 308320 319870 308372
rect 320174 308320 320180 308372
rect 320232 308360 320238 308372
rect 321186 308360 321192 308372
rect 320232 308332 321192 308360
rect 320232 308320 320238 308332
rect 321186 308320 321192 308332
rect 321244 308320 321250 308372
rect 355318 308320 355324 308372
rect 355376 308360 355382 308372
rect 367462 308360 367468 308372
rect 355376 308332 367468 308360
rect 355376 308320 355382 308332
rect 367462 308320 367468 308332
rect 367520 308320 367526 308372
rect 312170 308252 312176 308304
rect 312228 308292 312234 308304
rect 312446 308292 312452 308304
rect 312228 308264 312452 308292
rect 312228 308252 312234 308264
rect 312446 308252 312452 308264
rect 312504 308252 312510 308304
rect 313366 308252 313372 308304
rect 313424 308252 313430 308304
rect 314746 308252 314752 308304
rect 314804 308292 314810 308304
rect 315666 308292 315672 308304
rect 314804 308264 315672 308292
rect 314804 308252 314810 308264
rect 315666 308252 315672 308264
rect 315724 308252 315730 308304
rect 316586 308252 316592 308304
rect 316644 308252 316650 308304
rect 317690 308252 317696 308304
rect 317748 308292 317754 308304
rect 317874 308292 317880 308304
rect 317748 308264 317880 308292
rect 317748 308252 317754 308264
rect 317874 308252 317880 308264
rect 317932 308252 317938 308304
rect 318978 308252 318984 308304
rect 319036 308292 319042 308304
rect 319622 308292 319628 308304
rect 319036 308264 319628 308292
rect 319036 308252 319042 308264
rect 319622 308252 319628 308264
rect 319680 308252 319686 308304
rect 320358 308252 320364 308304
rect 320416 308292 320422 308304
rect 320634 308292 320640 308304
rect 320416 308264 320640 308292
rect 320416 308252 320422 308264
rect 320634 308252 320640 308264
rect 320692 308252 320698 308304
rect 353846 308252 353852 308304
rect 353904 308292 353910 308304
rect 366174 308292 366180 308304
rect 353904 308264 366180 308292
rect 353904 308252 353910 308264
rect 366174 308252 366180 308264
rect 366232 308252 366238 308304
rect 311894 308184 311900 308236
rect 311952 308224 311958 308236
rect 313182 308224 313188 308236
rect 311952 308196 313188 308224
rect 311952 308184 311958 308196
rect 313182 308184 313188 308196
rect 313240 308184 313246 308236
rect 313274 308184 313280 308236
rect 313332 308224 313338 308236
rect 314286 308224 314292 308236
rect 313332 308196 314292 308224
rect 313332 308184 313338 308196
rect 314286 308184 314292 308196
rect 314344 308184 314350 308236
rect 314654 308184 314660 308236
rect 314712 308224 314718 308236
rect 315482 308224 315488 308236
rect 314712 308196 315488 308224
rect 314712 308184 314718 308196
rect 315482 308184 315488 308196
rect 315540 308184 315546 308236
rect 311986 308116 311992 308168
rect 312044 308156 312050 308168
rect 312446 308156 312452 308168
rect 312044 308128 312452 308156
rect 312044 308116 312050 308128
rect 312446 308116 312452 308128
rect 312504 308116 312510 308168
rect 315022 308116 315028 308168
rect 315080 308156 315086 308168
rect 315298 308156 315304 308168
rect 315080 308128 315304 308156
rect 315080 308116 315086 308128
rect 315298 308116 315304 308128
rect 315356 308116 315362 308168
rect 316218 308116 316224 308168
rect 316276 308156 316282 308168
rect 316604 308156 316632 308252
rect 317322 308184 317328 308236
rect 317380 308224 317386 308236
rect 318058 308224 318064 308236
rect 317380 308196 318064 308224
rect 317380 308184 317386 308196
rect 318058 308184 318064 308196
rect 318116 308184 318122 308236
rect 318794 308184 318800 308236
rect 318852 308224 318858 308236
rect 319438 308224 319444 308236
rect 318852 308196 319444 308224
rect 318852 308184 318858 308196
rect 319438 308184 319444 308196
rect 319496 308184 319502 308236
rect 354950 308184 354956 308236
rect 355008 308224 355014 308236
rect 367278 308224 367284 308236
rect 355008 308196 367284 308224
rect 355008 308184 355014 308196
rect 367278 308184 367284 308196
rect 367336 308184 367342 308236
rect 316276 308128 316632 308156
rect 316276 308116 316282 308128
rect 317690 308116 317696 308168
rect 317748 308156 317754 308168
rect 318702 308156 318708 308168
rect 317748 308128 318708 308156
rect 317748 308116 317754 308128
rect 318702 308116 318708 308128
rect 318760 308116 318766 308168
rect 318886 308116 318892 308168
rect 318944 308156 318950 308168
rect 319990 308156 319996 308168
rect 318944 308128 319996 308156
rect 318944 308116 318950 308128
rect 319990 308116 319996 308128
rect 320048 308116 320054 308168
rect 320266 308116 320272 308168
rect 320324 308156 320330 308168
rect 320634 308156 320640 308168
rect 320324 308128 320640 308156
rect 320324 308116 320330 308128
rect 320634 308116 320640 308128
rect 320692 308116 320698 308168
rect 354582 308116 354588 308168
rect 354640 308156 354646 308168
rect 364794 308156 364800 308168
rect 354640 308128 364800 308156
rect 354640 308116 354646 308128
rect 364794 308116 364800 308128
rect 364852 308116 364858 308168
rect 252244 308060 253934 308088
rect 252244 308048 252250 308060
rect 259730 308048 259736 308100
rect 259788 308088 259794 308100
rect 260006 308088 260012 308100
rect 259788 308060 260012 308088
rect 259788 308048 259794 308060
rect 260006 308048 260012 308060
rect 260064 308048 260070 308100
rect 317506 308048 317512 308100
rect 317564 308088 317570 308100
rect 318518 308088 318524 308100
rect 317564 308060 318524 308088
rect 317564 308048 317570 308060
rect 318518 308048 318524 308060
rect 318576 308048 318582 308100
rect 245746 307980 245752 308032
rect 245804 308020 245810 308032
rect 251910 308020 251916 308032
rect 245804 307992 251916 308020
rect 245804 307980 245810 307992
rect 251910 307980 251916 307992
rect 251968 307980 251974 308032
rect 269482 307980 269488 308032
rect 269540 308020 269546 308032
rect 269758 308020 269764 308032
rect 269540 307992 269764 308020
rect 269540 307980 269546 307992
rect 269758 307980 269764 307992
rect 269816 307980 269822 308032
rect 285674 307980 285680 308032
rect 285732 308020 285738 308032
rect 285950 308020 285956 308032
rect 285732 307992 285956 308020
rect 285732 307980 285738 307992
rect 285950 307980 285956 307992
rect 286008 307980 286014 308032
rect 311986 307980 311992 308032
rect 312044 308020 312050 308032
rect 312814 308020 312820 308032
rect 312044 307992 312820 308020
rect 312044 307980 312050 307992
rect 312814 307980 312820 307992
rect 312872 307980 312878 308032
rect 316494 307980 316500 308032
rect 316552 308020 316558 308032
rect 316770 308020 316776 308032
rect 316552 307992 316776 308020
rect 316552 307980 316558 307992
rect 316770 307980 316776 307992
rect 316828 307980 316834 308032
rect 320266 307980 320272 308032
rect 320324 308020 320330 308032
rect 321370 308020 321376 308032
rect 320324 307992 321376 308020
rect 320324 307980 320330 307992
rect 321370 307980 321376 307992
rect 321428 307980 321434 308032
rect 360286 307980 360292 308032
rect 360344 308020 360350 308032
rect 360654 308020 360660 308032
rect 360344 307992 360660 308020
rect 360344 307980 360350 307992
rect 360654 307980 360660 307992
rect 360712 307980 360718 308032
rect 251818 307912 251824 307964
rect 251876 307952 251882 307964
rect 256510 307952 256516 307964
rect 251876 307924 256516 307952
rect 251876 307912 251882 307924
rect 256510 307912 256516 307924
rect 256568 307912 256574 307964
rect 317782 307912 317788 307964
rect 317840 307952 317846 307964
rect 318150 307952 318156 307964
rect 317840 307924 318156 307952
rect 317840 307912 317846 307924
rect 318150 307912 318156 307924
rect 318208 307912 318214 307964
rect 320450 307912 320456 307964
rect 320508 307952 320514 307964
rect 321002 307952 321008 307964
rect 320508 307924 321008 307952
rect 320508 307912 320514 307924
rect 321002 307912 321008 307924
rect 321060 307912 321066 307964
rect 360470 307912 360476 307964
rect 360528 307952 360534 307964
rect 361206 307952 361212 307964
rect 360528 307924 361212 307952
rect 360528 307912 360534 307924
rect 361206 307912 361212 307924
rect 361264 307912 361270 307964
rect 243998 307844 244004 307896
rect 244056 307884 244062 307896
rect 249242 307884 249248 307896
rect 244056 307856 249248 307884
rect 244056 307844 244062 307856
rect 249242 307844 249248 307856
rect 249300 307844 249306 307896
rect 250530 307844 250536 307896
rect 250588 307884 250594 307896
rect 250588 307856 251496 307884
rect 250588 307844 250594 307856
rect 242802 307776 242808 307828
rect 242860 307816 242866 307828
rect 243538 307816 243544 307828
rect 242860 307788 243544 307816
rect 242860 307776 242866 307788
rect 243538 307776 243544 307788
rect 243596 307776 243602 307828
rect 247770 307776 247776 307828
rect 247828 307816 247834 307828
rect 248506 307816 248512 307828
rect 247828 307788 248512 307816
rect 247828 307776 247834 307788
rect 248506 307776 248512 307788
rect 248564 307776 248570 307828
rect 250898 307776 250904 307828
rect 250956 307816 250962 307828
rect 251358 307816 251364 307828
rect 250956 307788 251364 307816
rect 250956 307776 250962 307788
rect 251358 307776 251364 307788
rect 251416 307776 251422 307828
rect 251468 307816 251496 307856
rect 253382 307844 253388 307896
rect 253440 307884 253446 307896
rect 259546 307884 259552 307896
rect 253440 307856 259552 307884
rect 253440 307844 253446 307856
rect 259546 307844 259552 307856
rect 259604 307844 259610 307896
rect 261754 307844 261760 307896
rect 261812 307884 261818 307896
rect 269850 307884 269856 307896
rect 261812 307856 269856 307884
rect 261812 307844 261818 307856
rect 269850 307844 269856 307856
rect 269908 307844 269914 307896
rect 337010 307844 337016 307896
rect 337068 307884 337074 307896
rect 337286 307884 337292 307896
rect 337068 307856 337292 307884
rect 337068 307844 337074 307856
rect 337286 307844 337292 307856
rect 337344 307844 337350 307896
rect 353386 307844 353392 307896
rect 353444 307884 353450 307896
rect 360930 307884 360936 307896
rect 353444 307856 360936 307884
rect 353444 307844 353450 307856
rect 360930 307844 360936 307856
rect 360988 307844 360994 307896
rect 257798 307816 257804 307828
rect 251468 307788 257804 307816
rect 257798 307776 257804 307788
rect 257856 307776 257862 307828
rect 348418 307776 348424 307828
rect 348476 307816 348482 307828
rect 350350 307816 350356 307828
rect 348476 307788 350356 307816
rect 348476 307776 348482 307788
rect 350350 307776 350356 307788
rect 350408 307776 350414 307828
rect 353018 307776 353024 307828
rect 353076 307816 353082 307828
rect 363506 307816 363512 307828
rect 353076 307788 363512 307816
rect 353076 307776 353082 307788
rect 363506 307776 363512 307788
rect 363564 307776 363570 307828
rect 227162 307708 227168 307760
rect 227220 307748 227226 307760
rect 243722 307748 243728 307760
rect 227220 307720 243728 307748
rect 227220 307708 227226 307720
rect 243722 307708 243728 307720
rect 243780 307708 243786 307760
rect 225782 307640 225788 307692
rect 225840 307680 225846 307692
rect 241974 307680 241980 307692
rect 225840 307652 241980 307680
rect 225840 307640 225846 307652
rect 241974 307640 241980 307652
rect 242032 307640 242038 307692
rect 229830 307572 229836 307624
rect 229888 307612 229894 307624
rect 252278 307612 252284 307624
rect 229888 307584 252284 307612
rect 229888 307572 229894 307584
rect 252278 307572 252284 307584
rect 252336 307572 252342 307624
rect 175918 307504 175924 307556
rect 175976 307544 175982 307556
rect 244826 307544 244832 307556
rect 175976 307516 244832 307544
rect 175976 307504 175982 307516
rect 244826 307504 244832 307516
rect 244884 307504 244890 307556
rect 220078 307436 220084 307488
rect 220136 307476 220142 307488
rect 242526 307476 242532 307488
rect 220136 307448 242532 307476
rect 220136 307436 220142 307448
rect 242526 307436 242532 307448
rect 242584 307436 242590 307488
rect 229738 307368 229744 307420
rect 229796 307408 229802 307420
rect 251726 307408 251732 307420
rect 229796 307380 251732 307408
rect 229796 307368 229802 307380
rect 251726 307368 251732 307380
rect 251784 307368 251790 307420
rect 228450 307300 228456 307352
rect 228508 307340 228514 307352
rect 247126 307340 247132 307352
rect 228508 307312 247132 307340
rect 228508 307300 228514 307312
rect 247126 307300 247132 307312
rect 247184 307300 247190 307352
rect 315390 307300 315396 307352
rect 315448 307340 315454 307352
rect 373258 307340 373264 307352
rect 315448 307312 373264 307340
rect 315448 307300 315454 307312
rect 373258 307300 373264 307312
rect 373316 307300 373322 307352
rect 172422 307232 172428 307284
rect 172480 307272 172486 307284
rect 246942 307272 246948 307284
rect 172480 307244 246948 307272
rect 172480 307232 172486 307244
rect 246942 307232 246948 307244
rect 247000 307232 247006 307284
rect 313550 307232 313556 307284
rect 313608 307272 313614 307284
rect 313826 307272 313832 307284
rect 313608 307244 313832 307272
rect 313608 307232 313614 307244
rect 313826 307232 313832 307244
rect 313884 307232 313890 307284
rect 317966 307232 317972 307284
rect 318024 307272 318030 307284
rect 402974 307272 402980 307284
rect 318024 307244 402980 307272
rect 318024 307232 318030 307244
rect 402974 307232 402980 307244
rect 403032 307232 403038 307284
rect 170490 307164 170496 307216
rect 170548 307204 170554 307216
rect 249978 307204 249984 307216
rect 170548 307176 249984 307204
rect 170548 307164 170554 307176
rect 249978 307164 249984 307176
rect 250036 307164 250042 307216
rect 295610 307164 295616 307216
rect 295668 307204 295674 307216
rect 295886 307204 295892 307216
rect 295668 307176 295892 307204
rect 295668 307164 295674 307176
rect 295886 307164 295892 307176
rect 295944 307164 295950 307216
rect 323670 307164 323676 307216
rect 323728 307204 323734 307216
rect 427078 307204 427084 307216
rect 323728 307176 427084 307204
rect 323728 307164 323734 307176
rect 427078 307164 427084 307176
rect 427136 307164 427142 307216
rect 170582 307096 170588 307148
rect 170640 307136 170646 307148
rect 238386 307136 238392 307148
rect 170640 307108 238392 307136
rect 170640 307096 170646 307108
rect 238386 307096 238392 307108
rect 238444 307096 238450 307148
rect 313550 307096 313556 307148
rect 313608 307136 313614 307148
rect 314470 307136 314476 307148
rect 313608 307108 314476 307136
rect 313608 307096 313614 307108
rect 314470 307096 314476 307108
rect 314528 307096 314534 307148
rect 330110 307096 330116 307148
rect 330168 307136 330174 307148
rect 480254 307136 480260 307148
rect 330168 307108 480260 307136
rect 330168 307096 330174 307108
rect 480254 307096 480260 307108
rect 480312 307096 480318 307148
rect 200114 307028 200120 307080
rect 200172 307068 200178 307080
rect 284938 307068 284944 307080
rect 200172 307040 284944 307068
rect 200172 307028 200178 307040
rect 284938 307028 284944 307040
rect 284996 307028 285002 307080
rect 316402 307028 316408 307080
rect 316460 307068 316466 307080
rect 317138 307068 317144 307080
rect 316460 307040 317144 307068
rect 316460 307028 316466 307040
rect 317138 307028 317144 307040
rect 317196 307028 317202 307080
rect 340414 307028 340420 307080
rect 340472 307068 340478 307080
rect 543734 307068 543740 307080
rect 340472 307040 543740 307068
rect 340472 307028 340478 307040
rect 543734 307028 543740 307040
rect 543792 307028 543798 307080
rect 170398 306960 170404 307012
rect 170456 307000 170462 307012
rect 239674 307000 239680 307012
rect 170456 306972 239680 307000
rect 170456 306960 170462 306972
rect 239674 306960 239680 306972
rect 239732 306960 239738 307012
rect 262582 306960 262588 307012
rect 262640 306960 262646 307012
rect 267918 306960 267924 307012
rect 267976 306960 267982 307012
rect 276382 306960 276388 307012
rect 276440 306960 276446 307012
rect 292758 306960 292764 307012
rect 292816 307000 292822 307012
rect 293402 307000 293408 307012
rect 292816 306972 293408 307000
rect 292816 306960 292822 306972
rect 293402 306960 293408 306972
rect 293460 306960 293466 307012
rect 321830 306960 321836 307012
rect 321888 307000 321894 307012
rect 322106 307000 322112 307012
rect 321888 306972 322112 307000
rect 321888 306960 321894 306972
rect 322106 306960 322112 306972
rect 322164 306960 322170 307012
rect 262600 306796 262628 306960
rect 262674 306796 262680 306808
rect 262600 306768 262680 306796
rect 262674 306756 262680 306768
rect 262732 306756 262738 306808
rect 267936 306796 267964 306960
rect 268010 306796 268016 306808
rect 267936 306768 268016 306796
rect 268010 306756 268016 306768
rect 268068 306756 268074 306808
rect 276400 306796 276428 306960
rect 287054 306824 287060 306876
rect 287112 306864 287118 306876
rect 287330 306864 287336 306876
rect 287112 306836 287336 306864
rect 287112 306824 287118 306836
rect 287330 306824 287336 306836
rect 287388 306824 287394 306876
rect 276474 306796 276480 306808
rect 276400 306768 276480 306796
rect 276474 306756 276480 306768
rect 276532 306756 276538 306808
rect 277670 306688 277676 306740
rect 277728 306688 277734 306740
rect 324406 306688 324412 306740
rect 324464 306728 324470 306740
rect 325050 306728 325056 306740
rect 324464 306700 325056 306728
rect 324464 306688 324470 306700
rect 325050 306688 325056 306700
rect 325108 306688 325114 306740
rect 260834 306552 260840 306604
rect 260892 306592 260898 306604
rect 261294 306592 261300 306604
rect 260892 306564 261300 306592
rect 260892 306552 260898 306564
rect 261294 306552 261300 306564
rect 261352 306552 261358 306604
rect 238938 306484 238944 306536
rect 238996 306524 239002 306536
rect 239858 306524 239864 306536
rect 238996 306496 239864 306524
rect 238996 306484 239002 306496
rect 239858 306484 239864 306496
rect 239916 306484 239922 306536
rect 255314 306484 255320 306536
rect 255372 306524 255378 306536
rect 255866 306524 255872 306536
rect 255372 306496 255872 306524
rect 255372 306484 255378 306496
rect 255866 306484 255872 306496
rect 255924 306484 255930 306536
rect 267826 306484 267832 306536
rect 267884 306524 267890 306536
rect 268102 306524 268108 306536
rect 267884 306496 268108 306524
rect 267884 306484 267890 306496
rect 268102 306484 268108 306496
rect 268160 306484 268166 306536
rect 277688 306468 277716 306688
rect 295794 306552 295800 306604
rect 295852 306552 295858 306604
rect 327166 306552 327172 306604
rect 327224 306592 327230 306604
rect 327626 306592 327632 306604
rect 327224 306564 327632 306592
rect 327224 306552 327230 306564
rect 327626 306552 327632 306564
rect 327684 306552 327690 306604
rect 357526 306552 357532 306604
rect 357584 306592 357590 306604
rect 357986 306592 357992 306604
rect 357584 306564 357992 306592
rect 357584 306552 357590 306564
rect 357986 306552 357992 306564
rect 358044 306552 358050 306604
rect 278774 306484 278780 306536
rect 278832 306524 278838 306536
rect 279786 306524 279792 306536
rect 278832 306496 279792 306524
rect 278832 306484 278838 306496
rect 279786 306484 279792 306496
rect 279844 306484 279850 306536
rect 282730 306484 282736 306536
rect 282788 306524 282794 306536
rect 288526 306524 288532 306536
rect 282788 306496 288532 306524
rect 282788 306484 282794 306496
rect 288526 306484 288532 306496
rect 288584 306484 288590 306536
rect 294230 306484 294236 306536
rect 294288 306484 294294 306536
rect 239030 306416 239036 306468
rect 239088 306456 239094 306468
rect 240042 306456 240048 306468
rect 239088 306428 240048 306456
rect 239088 306416 239094 306428
rect 240042 306416 240048 306428
rect 240100 306416 240106 306468
rect 255498 306416 255504 306468
rect 255556 306456 255562 306468
rect 255958 306456 255964 306468
rect 255556 306428 255964 306456
rect 255556 306416 255562 306428
rect 255958 306416 255964 306428
rect 256016 306416 256022 306468
rect 259546 306416 259552 306468
rect 259604 306456 259610 306468
rect 260650 306456 260656 306468
rect 259604 306428 260656 306456
rect 259604 306416 259610 306428
rect 260650 306416 260656 306428
rect 260708 306416 260714 306468
rect 260926 306416 260932 306468
rect 260984 306456 260990 306468
rect 261202 306456 261208 306468
rect 260984 306428 261208 306456
rect 260984 306416 260990 306428
rect 261202 306416 261208 306428
rect 261260 306416 261266 306468
rect 263594 306416 263600 306468
rect 263652 306456 263658 306468
rect 263870 306456 263876 306468
rect 263652 306428 263876 306456
rect 263652 306416 263658 306428
rect 263870 306416 263876 306428
rect 263928 306416 263934 306468
rect 264146 306416 264152 306468
rect 264204 306456 264210 306468
rect 264422 306456 264428 306468
rect 264204 306428 264428 306456
rect 264204 306416 264210 306428
rect 264422 306416 264428 306428
rect 264480 306416 264486 306468
rect 266630 306416 266636 306468
rect 266688 306456 266694 306468
rect 266906 306456 266912 306468
rect 266688 306428 266912 306456
rect 266688 306416 266694 306428
rect 266906 306416 266912 306428
rect 266964 306416 266970 306468
rect 270678 306416 270684 306468
rect 270736 306456 270742 306468
rect 270954 306456 270960 306468
rect 270736 306428 270960 306456
rect 270736 306416 270742 306428
rect 270954 306416 270960 306428
rect 271012 306416 271018 306468
rect 273714 306416 273720 306468
rect 273772 306456 273778 306468
rect 274450 306456 274456 306468
rect 273772 306428 274456 306456
rect 273772 306416 273778 306428
rect 274450 306416 274456 306428
rect 274508 306416 274514 306468
rect 277670 306416 277676 306468
rect 277728 306416 277734 306468
rect 279050 306416 279056 306468
rect 279108 306456 279114 306468
rect 279418 306456 279424 306468
rect 279108 306428 279424 306456
rect 279108 306416 279114 306428
rect 279418 306416 279424 306428
rect 279476 306416 279482 306468
rect 280338 306416 280344 306468
rect 280396 306456 280402 306468
rect 280798 306456 280804 306468
rect 280396 306428 280804 306456
rect 280396 306416 280402 306428
rect 280798 306416 280804 306428
rect 280856 306416 280862 306468
rect 286042 306416 286048 306468
rect 286100 306416 286106 306468
rect 286226 306416 286232 306468
rect 286284 306416 286290 306468
rect 237374 306348 237380 306400
rect 237432 306388 237438 306400
rect 237926 306388 237932 306400
rect 237432 306360 237932 306388
rect 237432 306348 237438 306360
rect 237926 306348 237932 306360
rect 237984 306348 237990 306400
rect 238846 306348 238852 306400
rect 238904 306388 238910 306400
rect 239306 306388 239312 306400
rect 238904 306360 239312 306388
rect 238904 306348 238910 306360
rect 239306 306348 239312 306360
rect 239364 306348 239370 306400
rect 240226 306348 240232 306400
rect 240284 306388 240290 306400
rect 241422 306388 241428 306400
rect 240284 306360 241428 306388
rect 240284 306348 240290 306360
rect 241422 306348 241428 306360
rect 241480 306348 241486 306400
rect 243078 306348 243084 306400
rect 243136 306388 243142 306400
rect 244090 306388 244096 306400
rect 243136 306360 244096 306388
rect 243136 306348 243142 306360
rect 244090 306348 244096 306360
rect 244148 306348 244154 306400
rect 248506 306348 248512 306400
rect 248564 306388 248570 306400
rect 248874 306388 248880 306400
rect 248564 306360 248880 306388
rect 248564 306348 248570 306360
rect 248874 306348 248880 306360
rect 248932 306348 248938 306400
rect 249886 306348 249892 306400
rect 249944 306388 249950 306400
rect 250990 306388 250996 306400
rect 249944 306360 250996 306388
rect 249944 306348 249950 306360
rect 250990 306348 250996 306360
rect 251048 306348 251054 306400
rect 251726 306348 251732 306400
rect 251784 306388 251790 306400
rect 252094 306388 252100 306400
rect 251784 306360 252100 306388
rect 251784 306348 251790 306360
rect 252094 306348 252100 306360
rect 252152 306348 252158 306400
rect 252646 306348 252652 306400
rect 252704 306388 252710 306400
rect 253658 306388 253664 306400
rect 252704 306360 253664 306388
rect 252704 306348 252710 306360
rect 253658 306348 253664 306360
rect 253716 306348 253722 306400
rect 255590 306348 255596 306400
rect 255648 306388 255654 306400
rect 256142 306388 256148 306400
rect 255648 306360 256148 306388
rect 255648 306348 255654 306360
rect 256142 306348 256148 306360
rect 256200 306348 256206 306400
rect 256786 306348 256792 306400
rect 256844 306388 256850 306400
rect 257982 306388 257988 306400
rect 256844 306360 257988 306388
rect 256844 306348 256850 306360
rect 257982 306348 257988 306360
rect 258040 306348 258046 306400
rect 259638 306348 259644 306400
rect 259696 306388 259702 306400
rect 260466 306388 260472 306400
rect 259696 306360 260472 306388
rect 259696 306348 259702 306360
rect 260466 306348 260472 306360
rect 260524 306348 260530 306400
rect 261294 306348 261300 306400
rect 261352 306388 261358 306400
rect 261846 306388 261852 306400
rect 261352 306360 261852 306388
rect 261352 306348 261358 306360
rect 261846 306348 261852 306360
rect 261904 306348 261910 306400
rect 264054 306348 264060 306400
rect 264112 306388 264118 306400
rect 264882 306388 264888 306400
rect 264112 306360 264888 306388
rect 264112 306348 264118 306360
rect 264882 306348 264888 306360
rect 264940 306348 264946 306400
rect 265066 306348 265072 306400
rect 265124 306388 265130 306400
rect 265250 306388 265256 306400
rect 265124 306360 265256 306388
rect 265124 306348 265130 306360
rect 265250 306348 265256 306360
rect 265308 306348 265314 306400
rect 265342 306348 265348 306400
rect 265400 306388 265406 306400
rect 265618 306388 265624 306400
rect 265400 306360 265624 306388
rect 265400 306348 265406 306360
rect 265618 306348 265624 306360
rect 265676 306348 265682 306400
rect 267734 306348 267740 306400
rect 267792 306388 267798 306400
rect 268102 306388 268108 306400
rect 267792 306360 268108 306388
rect 267792 306348 267798 306360
rect 268102 306348 268108 306360
rect 268160 306348 268166 306400
rect 269206 306348 269212 306400
rect 269264 306388 269270 306400
rect 270218 306388 270224 306400
rect 269264 306360 270224 306388
rect 269264 306348 269270 306360
rect 270218 306348 270224 306360
rect 270276 306348 270282 306400
rect 272242 306348 272248 306400
rect 272300 306388 272306 306400
rect 273070 306388 273076 306400
rect 272300 306360 273076 306388
rect 272300 306348 272306 306360
rect 273070 306348 273076 306360
rect 273128 306348 273134 306400
rect 273622 306348 273628 306400
rect 273680 306388 273686 306400
rect 274082 306388 274088 306400
rect 273680 306360 274088 306388
rect 273680 306348 273686 306360
rect 274082 306348 274088 306360
rect 274140 306348 274146 306400
rect 274910 306348 274916 306400
rect 274968 306388 274974 306400
rect 275554 306388 275560 306400
rect 274968 306360 275560 306388
rect 274968 306348 274974 306360
rect 275554 306348 275560 306360
rect 275612 306348 275618 306400
rect 276106 306348 276112 306400
rect 276164 306388 276170 306400
rect 277302 306388 277308 306400
rect 276164 306360 277308 306388
rect 276164 306348 276170 306360
rect 277302 306348 277308 306360
rect 277360 306348 277366 306400
rect 277394 306348 277400 306400
rect 277452 306388 277458 306400
rect 278406 306388 278412 306400
rect 277452 306360 278412 306388
rect 277452 306348 277458 306360
rect 278406 306348 278412 306360
rect 278464 306348 278470 306400
rect 278866 306348 278872 306400
rect 278924 306388 278930 306400
rect 279142 306388 279148 306400
rect 278924 306360 279148 306388
rect 278924 306348 278930 306360
rect 279142 306348 279148 306360
rect 279200 306348 279206 306400
rect 282914 306348 282920 306400
rect 282972 306388 282978 306400
rect 283742 306388 283748 306400
rect 282972 306360 283748 306388
rect 282972 306348 282978 306360
rect 283742 306348 283748 306360
rect 283800 306348 283806 306400
rect 284386 306348 284392 306400
rect 284444 306388 284450 306400
rect 285122 306388 285128 306400
rect 284444 306360 285128 306388
rect 284444 306348 284450 306360
rect 285122 306348 285128 306360
rect 285180 306348 285186 306400
rect 285674 306348 285680 306400
rect 285732 306388 285738 306400
rect 286060 306388 286088 306416
rect 285732 306360 286088 306388
rect 285732 306348 285738 306360
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 94498 306320 94504 306332
rect 3384 306292 94504 306320
rect 3384 306280 3390 306292
rect 94498 306280 94504 306292
rect 94556 306280 94562 306332
rect 219066 306280 219072 306332
rect 219124 306320 219130 306332
rect 284202 306320 284208 306332
rect 219124 306292 284208 306320
rect 219124 306280 219130 306292
rect 284202 306280 284208 306292
rect 284260 306280 284266 306332
rect 284662 306280 284668 306332
rect 284720 306320 284726 306332
rect 285490 306320 285496 306332
rect 284720 306292 285496 306320
rect 284720 306280 284726 306292
rect 285490 306280 285496 306292
rect 285548 306280 285554 306332
rect 286244 306320 286272 306416
rect 287422 306320 287428 306332
rect 285876 306292 286272 306320
rect 287164 306292 287428 306320
rect 285876 306264 285904 306292
rect 287164 306264 287192 306292
rect 287422 306280 287428 306292
rect 287480 306280 287486 306332
rect 291562 306280 291568 306332
rect 291620 306320 291626 306332
rect 292206 306320 292212 306332
rect 291620 306292 292212 306320
rect 291620 306280 291626 306292
rect 292206 306280 292212 306292
rect 292264 306280 292270 306332
rect 293126 306280 293132 306332
rect 293184 306320 293190 306332
rect 293678 306320 293684 306332
rect 293184 306292 293684 306320
rect 293184 306280 293190 306292
rect 293678 306280 293684 306292
rect 293736 306280 293742 306332
rect 294248 306264 294276 306484
rect 295812 306400 295840 306552
rect 296714 306484 296720 306536
rect 296772 306524 296778 306536
rect 297174 306524 297180 306536
rect 296772 306496 297180 306524
rect 296772 306484 296778 306496
rect 297174 306484 297180 306496
rect 297232 306484 297238 306536
rect 362310 306524 362316 306536
rect 357406 306496 362316 306524
rect 296898 306416 296904 306468
rect 296956 306456 296962 306468
rect 297358 306456 297364 306468
rect 296956 306428 297364 306456
rect 296956 306416 296962 306428
rect 297358 306416 297364 306428
rect 297416 306416 297422 306468
rect 306834 306416 306840 306468
rect 306892 306416 306898 306468
rect 310606 306416 310612 306468
rect 310664 306456 310670 306468
rect 310882 306456 310888 306468
rect 310664 306428 310888 306456
rect 310664 306416 310670 306428
rect 310882 306416 310888 306428
rect 310940 306416 310946 306468
rect 325786 306416 325792 306468
rect 325844 306456 325850 306468
rect 326430 306456 326436 306468
rect 325844 306428 326436 306456
rect 325844 306416 325850 306428
rect 326430 306416 326436 306428
rect 326488 306416 326494 306468
rect 328546 306416 328552 306468
rect 328604 306456 328610 306468
rect 329374 306456 329380 306468
rect 328604 306428 329380 306456
rect 328604 306416 328610 306428
rect 329374 306416 329380 306428
rect 329432 306416 329438 306468
rect 331306 306416 331312 306468
rect 331364 306456 331370 306468
rect 331766 306456 331772 306468
rect 331364 306428 331772 306456
rect 331364 306416 331370 306428
rect 331766 306416 331772 306428
rect 331824 306416 331830 306468
rect 336826 306416 336832 306468
rect 336884 306456 336890 306468
rect 337194 306456 337200 306468
rect 336884 306428 337200 306456
rect 336884 306416 336890 306428
rect 337194 306416 337200 306428
rect 337252 306416 337258 306468
rect 339678 306416 339684 306468
rect 339736 306456 339742 306468
rect 339954 306456 339960 306468
rect 339736 306428 339960 306456
rect 339736 306416 339742 306428
rect 339954 306416 339960 306428
rect 340012 306416 340018 306468
rect 340874 306416 340880 306468
rect 340932 306456 340938 306468
rect 341426 306456 341432 306468
rect 340932 306428 341432 306456
rect 340932 306416 340938 306428
rect 341426 306416 341432 306428
rect 341484 306416 341490 306468
rect 345014 306416 345020 306468
rect 345072 306456 345078 306468
rect 345474 306456 345480 306468
rect 345072 306428 345480 306456
rect 345072 306416 345078 306428
rect 345474 306416 345480 306428
rect 345532 306416 345538 306468
rect 295794 306348 295800 306400
rect 295852 306348 295858 306400
rect 299658 306348 299664 306400
rect 299716 306388 299722 306400
rect 300394 306388 300400 306400
rect 299716 306360 300400 306388
rect 299716 306348 299722 306360
rect 300394 306348 300400 306360
rect 300452 306348 300458 306400
rect 300854 306348 300860 306400
rect 300912 306388 300918 306400
rect 301682 306388 301688 306400
rect 300912 306360 301688 306388
rect 300912 306348 300918 306360
rect 301682 306348 301688 306360
rect 301740 306348 301746 306400
rect 302418 306348 302424 306400
rect 302476 306388 302482 306400
rect 303246 306388 303252 306400
rect 302476 306360 303252 306388
rect 302476 306348 302482 306360
rect 303246 306348 303252 306360
rect 303304 306348 303310 306400
rect 303798 306348 303804 306400
rect 303856 306388 303862 306400
rect 304626 306388 304632 306400
rect 303856 306360 304632 306388
rect 303856 306348 303862 306360
rect 304626 306348 304632 306360
rect 304684 306348 304690 306400
rect 295518 306280 295524 306332
rect 295576 306320 295582 306332
rect 295978 306320 295984 306332
rect 295576 306292 295984 306320
rect 295576 306280 295582 306292
rect 295978 306280 295984 306292
rect 296036 306280 296042 306332
rect 298094 306280 298100 306332
rect 298152 306320 298158 306332
rect 298646 306320 298652 306332
rect 298152 306292 298652 306320
rect 298152 306280 298158 306292
rect 298646 306280 298652 306292
rect 298704 306280 298710 306332
rect 299566 306280 299572 306332
rect 299624 306320 299630 306332
rect 300210 306320 300216 306332
rect 299624 306292 300216 306320
rect 299624 306280 299630 306292
rect 300210 306280 300216 306292
rect 300268 306280 300274 306332
rect 302510 306280 302516 306332
rect 302568 306320 302574 306332
rect 303062 306320 303068 306332
rect 302568 306292 303068 306320
rect 302568 306280 302574 306292
rect 303062 306280 303068 306292
rect 303120 306280 303126 306332
rect 303706 306280 303712 306332
rect 303764 306320 303770 306332
rect 304350 306320 304356 306332
rect 303764 306292 304356 306320
rect 303764 306280 303770 306292
rect 304350 306280 304356 306292
rect 304408 306280 304414 306332
rect 216490 306212 216496 306264
rect 216548 306252 216554 306264
rect 216548 306224 283144 306252
rect 216548 306212 216554 306224
rect 171686 306144 171692 306196
rect 171744 306184 171750 306196
rect 245470 306184 245476 306196
rect 171744 306156 245476 306184
rect 171744 306144 171750 306156
rect 245470 306144 245476 306156
rect 245528 306144 245534 306196
rect 247218 306144 247224 306196
rect 247276 306184 247282 306196
rect 247862 306184 247868 306196
rect 247276 306156 247868 306184
rect 247276 306144 247282 306156
rect 247862 306144 247868 306156
rect 247920 306144 247926 306196
rect 251358 306144 251364 306196
rect 251416 306184 251422 306196
rect 252462 306184 252468 306196
rect 251416 306156 252468 306184
rect 251416 306144 251422 306156
rect 252462 306144 252468 306156
rect 252520 306144 252526 306196
rect 254026 306144 254032 306196
rect 254084 306184 254090 306196
rect 254762 306184 254768 306196
rect 254084 306156 254768 306184
rect 254084 306144 254090 306156
rect 254762 306144 254768 306156
rect 254820 306144 254826 306196
rect 255682 306144 255688 306196
rect 255740 306184 255746 306196
rect 256326 306184 256332 306196
rect 255740 306156 256332 306184
rect 255740 306144 255746 306156
rect 256326 306144 256332 306156
rect 256384 306144 256390 306196
rect 258074 306144 258080 306196
rect 258132 306184 258138 306196
rect 258534 306184 258540 306196
rect 258132 306156 258540 306184
rect 258132 306144 258138 306156
rect 258534 306144 258540 306156
rect 258592 306144 258598 306196
rect 259730 306144 259736 306196
rect 259788 306184 259794 306196
rect 260282 306184 260288 306196
rect 259788 306156 260288 306184
rect 259788 306144 259794 306156
rect 260282 306144 260288 306156
rect 260340 306144 260346 306196
rect 262582 306144 262588 306196
rect 262640 306184 262646 306196
rect 263318 306184 263324 306196
rect 262640 306156 263324 306184
rect 262640 306144 262646 306156
rect 263318 306144 263324 306156
rect 263376 306144 263382 306196
rect 263686 306144 263692 306196
rect 263744 306184 263750 306196
rect 264514 306184 264520 306196
rect 263744 306156 264520 306184
rect 263744 306144 263750 306156
rect 264514 306144 264520 306156
rect 264572 306144 264578 306196
rect 266722 306144 266728 306196
rect 266780 306184 266786 306196
rect 267366 306184 267372 306196
rect 266780 306156 267372 306184
rect 266780 306144 266786 306156
rect 267366 306144 267372 306156
rect 267424 306144 267430 306196
rect 267918 306144 267924 306196
rect 267976 306184 267982 306196
rect 268286 306184 268292 306196
rect 267976 306156 268292 306184
rect 267976 306144 267982 306156
rect 268286 306144 268292 306156
rect 268344 306144 268350 306196
rect 269114 306144 269120 306196
rect 269172 306184 269178 306196
rect 269482 306184 269488 306196
rect 269172 306156 269488 306184
rect 269172 306144 269178 306156
rect 269482 306144 269488 306156
rect 269540 306144 269546 306196
rect 270862 306144 270868 306196
rect 270920 306184 270926 306196
rect 271046 306184 271052 306196
rect 270920 306156 271052 306184
rect 270920 306144 270926 306156
rect 271046 306144 271052 306156
rect 271104 306144 271110 306196
rect 271966 306144 271972 306196
rect 272024 306184 272030 306196
rect 272518 306184 272524 306196
rect 272024 306156 272524 306184
rect 272024 306144 272030 306156
rect 272518 306144 272524 306156
rect 272576 306144 272582 306196
rect 273346 306144 273352 306196
rect 273404 306184 273410 306196
rect 274266 306184 274272 306196
rect 273404 306156 274272 306184
rect 273404 306144 273410 306156
rect 274266 306144 274272 306156
rect 274324 306144 274330 306196
rect 277486 306144 277492 306196
rect 277544 306184 277550 306196
rect 277854 306184 277860 306196
rect 277544 306156 277860 306184
rect 277544 306144 277550 306156
rect 277854 306144 277860 306156
rect 277912 306144 277918 306196
rect 279234 306144 279240 306196
rect 279292 306184 279298 306196
rect 279970 306184 279976 306196
rect 279292 306156 279976 306184
rect 279292 306144 279298 306156
rect 279970 306144 279976 306156
rect 280028 306144 280034 306196
rect 280062 306144 280068 306196
rect 280120 306184 280126 306196
rect 281534 306184 281540 306196
rect 280120 306156 281540 306184
rect 280120 306144 280126 306156
rect 281534 306144 281540 306156
rect 281592 306144 281598 306196
rect 283116 306184 283144 306224
rect 283374 306212 283380 306264
rect 283432 306252 283438 306264
rect 284018 306252 284024 306264
rect 283432 306224 284024 306252
rect 283432 306212 283438 306224
rect 284018 306212 284024 306224
rect 284076 306212 284082 306264
rect 284570 306212 284576 306264
rect 284628 306252 284634 306264
rect 285306 306252 285312 306264
rect 284628 306224 285312 306252
rect 284628 306212 284634 306224
rect 285306 306212 285312 306224
rect 285364 306212 285370 306264
rect 285858 306212 285864 306264
rect 285916 306212 285922 306264
rect 286134 306212 286140 306264
rect 286192 306252 286198 306264
rect 286870 306252 286876 306264
rect 286192 306224 286876 306252
rect 286192 306212 286198 306224
rect 286870 306212 286876 306224
rect 286928 306212 286934 306264
rect 287146 306212 287152 306264
rect 287204 306212 287210 306264
rect 287238 306212 287244 306264
rect 287296 306252 287302 306264
rect 287974 306252 287980 306264
rect 287296 306224 287980 306252
rect 287296 306212 287302 306224
rect 287974 306212 287980 306224
rect 288032 306212 288038 306264
rect 294230 306212 294236 306264
rect 294288 306212 294294 306264
rect 297174 306212 297180 306264
rect 297232 306252 297238 306264
rect 297910 306252 297916 306264
rect 297232 306224 297916 306252
rect 297232 306212 297238 306224
rect 297910 306212 297916 306224
rect 297968 306212 297974 306264
rect 300946 306212 300952 306264
rect 301004 306252 301010 306264
rect 302050 306252 302056 306264
rect 301004 306224 302056 306252
rect 301004 306212 301010 306224
rect 302050 306212 302056 306224
rect 302108 306212 302114 306264
rect 302326 306212 302332 306264
rect 302384 306252 302390 306264
rect 303430 306252 303436 306264
rect 302384 306224 303436 306252
rect 302384 306212 302390 306224
rect 303430 306212 303436 306224
rect 303488 306212 303494 306264
rect 305454 306212 305460 306264
rect 305512 306252 305518 306264
rect 305914 306252 305920 306264
rect 305512 306224 305920 306252
rect 305512 306212 305518 306224
rect 305914 306212 305920 306224
rect 305972 306212 305978 306264
rect 306650 306212 306656 306264
rect 306708 306252 306714 306264
rect 306852 306252 306880 306416
rect 328730 306348 328736 306400
rect 328788 306388 328794 306400
rect 329558 306388 329564 306400
rect 328788 306360 329564 306388
rect 328788 306348 328794 306360
rect 329558 306348 329564 306360
rect 329616 306348 329622 306400
rect 329834 306348 329840 306400
rect 329892 306388 329898 306400
rect 331122 306388 331128 306400
rect 329892 306360 331128 306388
rect 329892 306348 329898 306360
rect 331122 306348 331128 306360
rect 331180 306348 331186 306400
rect 331214 306348 331220 306400
rect 331272 306388 331278 306400
rect 332226 306388 332232 306400
rect 331272 306360 332232 306388
rect 331272 306348 331278 306360
rect 332226 306348 332232 306360
rect 332284 306348 332290 306400
rect 332594 306348 332600 306400
rect 332652 306388 332658 306400
rect 332870 306388 332876 306400
rect 332652 306360 332876 306388
rect 332652 306348 332658 306360
rect 332870 306348 332876 306360
rect 332928 306348 332934 306400
rect 333054 306348 333060 306400
rect 333112 306388 333118 306400
rect 333606 306388 333612 306400
rect 333112 306360 333612 306388
rect 333112 306348 333118 306360
rect 333606 306348 333612 306360
rect 333664 306348 333670 306400
rect 335354 306348 335360 306400
rect 335412 306388 335418 306400
rect 336090 306388 336096 306400
rect 335412 306360 336096 306388
rect 335412 306348 335418 306360
rect 336090 306348 336096 306360
rect 336148 306348 336154 306400
rect 336734 306348 336740 306400
rect 336792 306388 336798 306400
rect 337378 306388 337384 306400
rect 336792 306360 337384 306388
rect 336792 306348 336798 306360
rect 337378 306348 337384 306360
rect 337436 306348 337442 306400
rect 345106 306348 345112 306400
rect 345164 306388 345170 306400
rect 346210 306388 346216 306400
rect 345164 306360 346216 306388
rect 345164 306348 345170 306360
rect 346210 306348 346216 306360
rect 346268 306348 346274 306400
rect 347774 306348 347780 306400
rect 347832 306388 347838 306400
rect 349062 306388 349068 306400
rect 347832 306360 349068 306388
rect 347832 306348 347838 306360
rect 349062 306348 349068 306360
rect 349120 306348 349126 306400
rect 307938 306280 307944 306332
rect 307996 306320 308002 306332
rect 308950 306320 308956 306332
rect 307996 306292 308956 306320
rect 307996 306280 308002 306292
rect 308950 306280 308956 306292
rect 309008 306280 309014 306332
rect 310974 306280 310980 306332
rect 311032 306320 311038 306332
rect 311434 306320 311440 306332
rect 311032 306292 311440 306320
rect 311032 306280 311038 306292
rect 311434 306280 311440 306292
rect 311492 306280 311498 306332
rect 321830 306280 321836 306332
rect 321888 306320 321894 306332
rect 322658 306320 322664 306332
rect 321888 306292 322664 306320
rect 321888 306280 321894 306292
rect 322658 306280 322664 306292
rect 322716 306280 322722 306332
rect 325694 306280 325700 306332
rect 325752 306320 325758 306332
rect 326154 306320 326160 306332
rect 325752 306292 326160 306320
rect 325752 306280 325758 306292
rect 326154 306280 326160 306292
rect 326212 306280 326218 306332
rect 327534 306280 327540 306332
rect 327592 306320 327598 306332
rect 327810 306320 327816 306332
rect 327592 306292 327816 306320
rect 327592 306280 327598 306292
rect 327810 306280 327816 306292
rect 327868 306280 327874 306332
rect 328638 306280 328644 306332
rect 328696 306320 328702 306332
rect 329098 306320 329104 306332
rect 328696 306292 329104 306320
rect 328696 306280 328702 306292
rect 329098 306280 329104 306292
rect 329156 306280 329162 306332
rect 329926 306280 329932 306332
rect 329984 306320 329990 306332
rect 330938 306320 330944 306332
rect 329984 306292 330944 306320
rect 329984 306280 329990 306292
rect 330938 306280 330944 306292
rect 330996 306280 331002 306332
rect 331306 306280 331312 306332
rect 331364 306320 331370 306332
rect 332042 306320 332048 306332
rect 331364 306292 332048 306320
rect 331364 306280 331370 306292
rect 332042 306280 332048 306292
rect 332100 306280 332106 306332
rect 332962 306280 332968 306332
rect 333020 306320 333026 306332
rect 333238 306320 333244 306332
rect 333020 306292 333244 306320
rect 333020 306280 333026 306292
rect 333238 306280 333244 306292
rect 333296 306280 333302 306332
rect 335538 306280 335544 306332
rect 335596 306320 335602 306332
rect 336274 306320 336280 306332
rect 335596 306292 336280 306320
rect 335596 306280 335602 306292
rect 336274 306280 336280 306292
rect 336332 306280 336338 306332
rect 336918 306280 336924 306332
rect 336976 306320 336982 306332
rect 337746 306320 337752 306332
rect 336976 306292 337752 306320
rect 336976 306280 336982 306292
rect 337746 306280 337752 306292
rect 337804 306280 337810 306332
rect 338114 306280 338120 306332
rect 338172 306320 338178 306332
rect 338942 306320 338948 306332
rect 338172 306292 338948 306320
rect 338172 306280 338178 306292
rect 338942 306280 338948 306292
rect 339000 306280 339006 306332
rect 342254 306280 342260 306332
rect 342312 306320 342318 306332
rect 342898 306320 342904 306332
rect 342312 306292 342904 306320
rect 342312 306280 342318 306292
rect 342898 306280 342904 306292
rect 342956 306280 342962 306332
rect 343818 306280 343824 306332
rect 343876 306320 343882 306332
rect 344278 306320 344284 306332
rect 343876 306292 344284 306320
rect 343876 306280 343882 306292
rect 344278 306280 344284 306292
rect 344336 306280 344342 306332
rect 345014 306280 345020 306332
rect 345072 306320 345078 306332
rect 345750 306320 345756 306332
rect 345072 306292 345756 306320
rect 345072 306280 345078 306292
rect 345750 306280 345756 306292
rect 345808 306280 345814 306332
rect 347866 306280 347872 306332
rect 347924 306320 347930 306332
rect 348234 306320 348240 306332
rect 347924 306292 348240 306320
rect 347924 306280 347930 306292
rect 348234 306280 348240 306292
rect 348292 306280 348298 306332
rect 350534 306280 350540 306332
rect 350592 306320 350598 306332
rect 351546 306320 351552 306332
rect 350592 306292 351552 306320
rect 350592 306280 350598 306292
rect 351546 306280 351552 306292
rect 351604 306280 351610 306332
rect 353202 306280 353208 306332
rect 353260 306320 353266 306332
rect 357406 306320 357434 306496
rect 362310 306484 362316 306496
rect 362368 306484 362374 306536
rect 357618 306416 357624 306468
rect 357676 306416 357682 306468
rect 353260 306292 357434 306320
rect 353260 306280 353266 306292
rect 306708 306224 306880 306252
rect 306708 306212 306714 306224
rect 308030 306212 308036 306264
rect 308088 306252 308094 306264
rect 308582 306252 308588 306264
rect 308088 306224 308588 306252
rect 308088 306212 308094 306224
rect 308582 306212 308588 306224
rect 308640 306212 308646 306264
rect 311066 306212 311072 306264
rect 311124 306252 311130 306264
rect 311618 306252 311624 306264
rect 311124 306224 311624 306252
rect 311124 306212 311130 306224
rect 311618 306212 311624 306224
rect 311676 306212 311682 306264
rect 321554 306212 321560 306264
rect 321612 306252 321618 306264
rect 322014 306252 322020 306264
rect 321612 306224 322020 306252
rect 321612 306212 321618 306224
rect 322014 306212 322020 306224
rect 322072 306212 322078 306264
rect 322934 306212 322940 306264
rect 322992 306252 322998 306264
rect 323486 306252 323492 306264
rect 322992 306224 323492 306252
rect 322992 306212 322998 306224
rect 323486 306212 323492 306224
rect 323544 306212 323550 306264
rect 325878 306212 325884 306264
rect 325936 306252 325942 306264
rect 326890 306252 326896 306264
rect 325936 306224 326896 306252
rect 325936 306212 325942 306224
rect 326890 306212 326896 306224
rect 326948 306212 326954 306264
rect 328822 306212 328828 306264
rect 328880 306252 328886 306264
rect 329006 306252 329012 306264
rect 328880 306224 329012 306252
rect 328880 306212 328886 306224
rect 329006 306212 329012 306224
rect 329064 306212 329070 306264
rect 332594 306212 332600 306264
rect 332652 306252 332658 306264
rect 333790 306252 333796 306264
rect 332652 306224 333796 306252
rect 332652 306212 332658 306224
rect 333790 306212 333796 306224
rect 333848 306212 333854 306264
rect 335446 306212 335452 306264
rect 335504 306252 335510 306264
rect 336642 306252 336648 306264
rect 335504 306224 336648 306252
rect 335504 306212 335510 306224
rect 336642 306212 336648 306224
rect 336700 306212 336706 306264
rect 336826 306212 336832 306264
rect 336884 306252 336890 306264
rect 337930 306252 337936 306264
rect 336884 306224 337936 306252
rect 336884 306212 336890 306224
rect 337930 306212 337936 306224
rect 337988 306212 337994 306264
rect 338482 306212 338488 306264
rect 338540 306252 338546 306264
rect 339310 306252 339316 306264
rect 338540 306224 339316 306252
rect 338540 306212 338546 306224
rect 339310 306212 339316 306224
rect 339368 306212 339374 306264
rect 339678 306212 339684 306264
rect 339736 306252 339742 306264
rect 340046 306252 340052 306264
rect 339736 306224 340052 306252
rect 339736 306212 339742 306224
rect 340046 306212 340052 306224
rect 340104 306212 340110 306264
rect 341058 306212 341064 306264
rect 341116 306252 341122 306264
rect 341426 306252 341432 306264
rect 341116 306224 341432 306252
rect 341116 306212 341122 306224
rect 341426 306212 341432 306224
rect 341484 306212 341490 306264
rect 342714 306212 342720 306264
rect 342772 306252 342778 306264
rect 343266 306252 343272 306264
rect 342772 306224 343272 306252
rect 342772 306212 342778 306224
rect 343266 306212 343272 306224
rect 343324 306212 343330 306264
rect 345290 306252 345296 306264
rect 345216 306224 345296 306252
rect 289078 306184 289084 306196
rect 283116 306156 289084 306184
rect 289078 306144 289084 306156
rect 289136 306144 289142 306196
rect 295702 306144 295708 306196
rect 295760 306184 295766 306196
rect 296530 306184 296536 306196
rect 295760 306156 296536 306184
rect 295760 306144 295766 306156
rect 296530 306144 296536 306156
rect 296588 306144 296594 306196
rect 301038 306144 301044 306196
rect 301096 306184 301102 306196
rect 301866 306184 301872 306196
rect 301096 306156 301872 306184
rect 301096 306144 301102 306156
rect 301866 306144 301872 306156
rect 301924 306144 301930 306196
rect 303982 306144 303988 306196
rect 304040 306144 304046 306196
rect 305362 306144 305368 306196
rect 305420 306184 305426 306196
rect 305730 306184 305736 306196
rect 305420 306156 305736 306184
rect 305420 306144 305426 306156
rect 305730 306144 305736 306156
rect 305788 306144 305794 306196
rect 306374 306144 306380 306196
rect 306432 306184 306438 306196
rect 306834 306184 306840 306196
rect 306432 306156 306840 306184
rect 306432 306144 306438 306156
rect 306834 306144 306840 306156
rect 306892 306144 306898 306196
rect 307846 306144 307852 306196
rect 307904 306184 307910 306196
rect 308398 306184 308404 306196
rect 307904 306156 308404 306184
rect 307904 306144 307910 306156
rect 308398 306144 308404 306156
rect 308456 306144 308462 306196
rect 310698 306144 310704 306196
rect 310756 306184 310762 306196
rect 311342 306184 311348 306196
rect 310756 306156 311348 306184
rect 310756 306144 310762 306156
rect 311342 306144 311348 306156
rect 311400 306144 311406 306196
rect 321738 306144 321744 306196
rect 321796 306184 321802 306196
rect 322474 306184 322480 306196
rect 321796 306156 322480 306184
rect 321796 306144 321802 306156
rect 322474 306144 322480 306156
rect 322532 306144 322538 306196
rect 324590 306144 324596 306196
rect 324648 306184 324654 306196
rect 325602 306184 325608 306196
rect 324648 306156 325608 306184
rect 324648 306144 324654 306156
rect 325602 306144 325608 306156
rect 325660 306144 325666 306196
rect 328638 306144 328644 306196
rect 328696 306184 328702 306196
rect 329190 306184 329196 306196
rect 328696 306156 329196 306184
rect 328696 306144 328702 306156
rect 329190 306144 329196 306156
rect 329248 306144 329254 306196
rect 332778 306144 332784 306196
rect 332836 306184 332842 306196
rect 333422 306184 333428 306196
rect 332836 306156 333428 306184
rect 332836 306144 332842 306156
rect 333422 306144 333428 306156
rect 333480 306144 333486 306196
rect 333974 306144 333980 306196
rect 334032 306184 334038 306196
rect 334434 306184 334440 306196
rect 334032 306156 334440 306184
rect 334032 306144 334038 306156
rect 334434 306144 334440 306156
rect 334492 306144 334498 306196
rect 334526 306144 334532 306196
rect 334584 306184 334590 306196
rect 334894 306184 334900 306196
rect 334584 306156 334900 306184
rect 334584 306144 334590 306156
rect 334894 306144 334900 306156
rect 334952 306144 334958 306196
rect 338206 306144 338212 306196
rect 338264 306184 338270 306196
rect 338666 306184 338672 306196
rect 338264 306156 338672 306184
rect 338264 306144 338270 306156
rect 338666 306144 338672 306156
rect 338724 306144 338730 306196
rect 339494 306144 339500 306196
rect 339552 306184 339558 306196
rect 340230 306184 340236 306196
rect 339552 306156 340236 306184
rect 339552 306144 339558 306156
rect 340230 306144 340236 306156
rect 340288 306144 340294 306196
rect 340966 306144 340972 306196
rect 341024 306184 341030 306196
rect 341518 306184 341524 306196
rect 341024 306156 341524 306184
rect 341024 306144 341030 306156
rect 341518 306144 341524 306156
rect 341576 306144 341582 306196
rect 215202 306076 215208 306128
rect 215260 306116 215266 306128
rect 282730 306116 282736 306128
rect 215260 306088 282736 306116
rect 215260 306076 215266 306088
rect 282730 306076 282736 306088
rect 282788 306076 282794 306128
rect 295610 306076 295616 306128
rect 295668 306116 295674 306128
rect 296346 306116 296352 306128
rect 295668 306088 296352 306116
rect 295668 306076 295674 306088
rect 296346 306076 296352 306088
rect 296404 306076 296410 306128
rect 219158 306008 219164 306060
rect 219216 306048 219222 306060
rect 282546 306048 282552 306060
rect 219216 306020 282552 306048
rect 219216 306008 219222 306020
rect 282546 306008 282552 306020
rect 282604 306008 282610 306060
rect 283650 306008 283656 306060
rect 283708 306048 283714 306060
rect 293494 306048 293500 306060
rect 283708 306020 293500 306048
rect 283708 306008 283714 306020
rect 293494 306008 293500 306020
rect 293552 306008 293558 306060
rect 304000 305992 304028 306144
rect 304994 306076 305000 306128
rect 305052 306116 305058 306128
rect 305638 306116 305644 306128
rect 305052 306088 305644 306116
rect 305052 306076 305058 306088
rect 305638 306076 305644 306088
rect 305696 306076 305702 306128
rect 306558 306076 306564 306128
rect 306616 306116 306622 306128
rect 307294 306116 307300 306128
rect 306616 306088 307300 306116
rect 306616 306076 306622 306088
rect 307294 306076 307300 306088
rect 307352 306076 307358 306128
rect 309226 306076 309232 306128
rect 309284 306116 309290 306128
rect 309686 306116 309692 306128
rect 309284 306088 309692 306116
rect 309284 306076 309290 306088
rect 309686 306076 309692 306088
rect 309744 306076 309750 306128
rect 310790 306076 310796 306128
rect 310848 306116 310854 306128
rect 311802 306116 311808 306128
rect 310848 306088 311808 306116
rect 310848 306076 310854 306088
rect 311802 306076 311808 306088
rect 311860 306076 311866 306128
rect 321554 306076 321560 306128
rect 321612 306116 321618 306128
rect 322290 306116 322296 306128
rect 321612 306088 322296 306116
rect 321612 306076 321618 306088
rect 322290 306076 322296 306088
rect 322348 306076 322354 306128
rect 323210 306076 323216 306128
rect 323268 306116 323274 306128
rect 324038 306116 324044 306128
rect 323268 306088 324044 306116
rect 323268 306076 323274 306088
rect 324038 306076 324044 306088
rect 324096 306076 324102 306128
rect 324498 306076 324504 306128
rect 324556 306116 324562 306128
rect 325234 306116 325240 306128
rect 324556 306088 325240 306116
rect 324556 306076 324562 306088
rect 325234 306076 325240 306088
rect 325292 306076 325298 306128
rect 327166 306076 327172 306128
rect 327224 306116 327230 306128
rect 327902 306116 327908 306128
rect 327224 306088 327908 306116
rect 327224 306076 327230 306088
rect 327902 306076 327908 306088
rect 327960 306076 327966 306128
rect 328454 306076 328460 306128
rect 328512 306116 328518 306128
rect 329006 306116 329012 306128
rect 328512 306088 329012 306116
rect 328512 306076 328518 306088
rect 329006 306076 329012 306088
rect 329064 306076 329070 306128
rect 334158 306076 334164 306128
rect 334216 306116 334222 306128
rect 335078 306116 335084 306128
rect 334216 306088 335084 306116
rect 334216 306076 334222 306088
rect 335078 306076 335084 306088
rect 335136 306076 335142 306128
rect 339586 306076 339592 306128
rect 339644 306116 339650 306128
rect 340598 306116 340604 306128
rect 339644 306088 340604 306116
rect 339644 306076 339650 306088
rect 340598 306076 340604 306088
rect 340656 306076 340662 306128
rect 341058 306076 341064 306128
rect 341116 306116 341122 306128
rect 341794 306116 341800 306128
rect 341116 306088 341800 306116
rect 341116 306076 341122 306088
rect 341794 306076 341800 306088
rect 341852 306076 341858 306128
rect 342438 306076 342444 306128
rect 342496 306116 342502 306128
rect 343082 306116 343088 306128
rect 342496 306088 343088 306116
rect 342496 306076 342502 306088
rect 343082 306076 343088 306088
rect 343140 306076 343146 306128
rect 305086 306008 305092 306060
rect 305144 306048 305150 306060
rect 306282 306048 306288 306060
rect 305144 306020 306288 306048
rect 305144 306008 305150 306020
rect 306282 306008 306288 306020
rect 306340 306008 306346 306060
rect 306374 306008 306380 306060
rect 306432 306048 306438 306060
rect 307202 306048 307208 306060
rect 306432 306020 307208 306048
rect 306432 306008 306438 306020
rect 307202 306008 307208 306020
rect 307260 306008 307266 306060
rect 309134 306008 309140 306060
rect 309192 306048 309198 306060
rect 309594 306048 309600 306060
rect 309192 306020 309600 306048
rect 309192 306008 309198 306020
rect 309594 306008 309600 306020
rect 309652 306008 309658 306060
rect 323118 306008 323124 306060
rect 323176 306048 323182 306060
rect 323854 306048 323860 306060
rect 323176 306020 323860 306048
rect 323176 306008 323182 306020
rect 323854 306008 323860 306020
rect 323912 306008 323918 306060
rect 327258 306008 327264 306060
rect 327316 306048 327322 306060
rect 328270 306048 328276 306060
rect 327316 306020 328276 306048
rect 327316 306008 327322 306020
rect 328270 306008 328276 306020
rect 328328 306008 328334 306060
rect 334434 306008 334440 306060
rect 334492 306048 334498 306060
rect 335262 306048 335268 306060
rect 334492 306020 335268 306048
rect 334492 306008 334498 306020
rect 335262 306008 335268 306020
rect 335320 306008 335326 306060
rect 338206 306008 338212 306060
rect 338264 306048 338270 306060
rect 339126 306048 339132 306060
rect 338264 306020 339132 306048
rect 338264 306008 338270 306020
rect 339126 306008 339132 306020
rect 339184 306008 339190 306060
rect 340966 306008 340972 306060
rect 341024 306048 341030 306060
rect 341978 306048 341984 306060
rect 341024 306020 341984 306048
rect 341024 306008 341030 306020
rect 341978 306008 341984 306020
rect 342036 306008 342042 306060
rect 342346 306008 342352 306060
rect 342404 306048 342410 306060
rect 343358 306048 343364 306060
rect 342404 306020 343364 306048
rect 342404 306008 342410 306020
rect 343358 306008 343364 306020
rect 343416 306008 343422 306060
rect 345216 305992 345244 306224
rect 345290 306212 345296 306224
rect 345348 306212 345354 306264
rect 356514 306212 356520 306264
rect 356572 306252 356578 306264
rect 356790 306252 356796 306264
rect 356572 306224 356796 306252
rect 356572 306212 356578 306224
rect 356790 306212 356796 306224
rect 356848 306212 356854 306264
rect 357636 306252 357664 306416
rect 357802 306348 357808 306400
rect 357860 306388 357866 306400
rect 357986 306388 357992 306400
rect 357860 306360 357992 306388
rect 357860 306348 357866 306360
rect 357986 306348 357992 306360
rect 358044 306348 358050 306400
rect 359642 306348 359648 306400
rect 359700 306388 359706 306400
rect 359700 306360 360148 306388
rect 359700 306348 359706 306360
rect 360120 306320 360148 306360
rect 366358 306320 366364 306332
rect 360120 306292 366364 306320
rect 366358 306280 366364 306292
rect 366416 306280 366422 306332
rect 357710 306252 357716 306264
rect 357636 306224 357716 306252
rect 357710 306212 357716 306224
rect 357768 306212 357774 306264
rect 371602 306252 371608 306264
rect 358464 306224 371608 306252
rect 356330 306144 356336 306196
rect 356388 306184 356394 306196
rect 358464 306184 358492 306224
rect 371602 306212 371608 306224
rect 371660 306212 371666 306264
rect 368934 306184 368940 306196
rect 356388 306156 358492 306184
rect 358556 306156 368940 306184
rect 356388 306144 356394 306156
rect 357434 306076 357440 306128
rect 357492 306116 357498 306128
rect 357894 306116 357900 306128
rect 357492 306088 357900 306116
rect 357492 306076 357498 306088
rect 357894 306076 357900 306088
rect 357952 306076 357958 306128
rect 354030 306008 354036 306060
rect 354088 306048 354094 306060
rect 358556 306048 358584 306156
rect 368934 306144 368940 306156
rect 368992 306144 368998 306196
rect 359274 306076 359280 306128
rect 359332 306116 359338 306128
rect 359734 306116 359740 306128
rect 359332 306088 359740 306116
rect 359332 306076 359338 306088
rect 359734 306076 359740 306088
rect 359792 306076 359798 306128
rect 359826 306076 359832 306128
rect 359884 306116 359890 306128
rect 369026 306116 369032 306128
rect 359884 306088 369032 306116
rect 359884 306076 359890 306088
rect 369026 306076 369032 306088
rect 369084 306076 369090 306128
rect 354088 306020 358584 306048
rect 354088 306008 354094 306020
rect 359366 306008 359372 306060
rect 359424 306048 359430 306060
rect 359918 306048 359924 306060
rect 359424 306020 359924 306048
rect 359424 306008 359430 306020
rect 359918 306008 359924 306020
rect 359976 306008 359982 306060
rect 362310 306008 362316 306060
rect 362368 306048 362374 306060
rect 368750 306048 368756 306060
rect 362368 306020 368756 306048
rect 362368 306008 362374 306020
rect 368750 306008 368756 306020
rect 368808 306008 368814 306060
rect 214926 305940 214932 305992
rect 214984 305980 214990 305992
rect 282362 305980 282368 305992
rect 214984 305952 282368 305980
rect 214984 305940 214990 305952
rect 282362 305940 282368 305952
rect 282420 305940 282426 305992
rect 284202 305940 284208 305992
rect 284260 305980 284266 305992
rect 291838 305980 291844 305992
rect 284260 305952 291844 305980
rect 284260 305940 284266 305952
rect 291838 305940 291844 305952
rect 291896 305940 291902 305992
rect 303982 305940 303988 305992
rect 304040 305940 304046 305992
rect 328454 305940 328460 305992
rect 328512 305980 328518 305992
rect 329742 305980 329748 305992
rect 328512 305952 329748 305980
rect 328512 305940 328518 305952
rect 329742 305940 329748 305952
rect 329800 305940 329806 305992
rect 343910 305940 343916 305992
rect 343968 305980 343974 305992
rect 344186 305980 344192 305992
rect 343968 305952 344192 305980
rect 343968 305940 343974 305952
rect 344186 305940 344192 305952
rect 344244 305940 344250 305992
rect 345198 305940 345204 305992
rect 345256 305940 345262 305992
rect 345290 305940 345296 305992
rect 345348 305980 345354 305992
rect 345842 305980 345848 305992
rect 345348 305952 345848 305980
rect 345348 305940 345354 305952
rect 345842 305940 345848 305952
rect 345900 305940 345906 305992
rect 354766 305940 354772 305992
rect 354824 305980 354830 305992
rect 371510 305980 371516 305992
rect 354824 305952 371516 305980
rect 354824 305940 354830 305952
rect 371510 305940 371516 305952
rect 371568 305940 371574 305992
rect 216306 305872 216312 305924
rect 216364 305912 216370 305924
rect 282730 305912 282736 305924
rect 216364 305884 282736 305912
rect 216364 305872 216370 305884
rect 282730 305872 282736 305884
rect 282788 305872 282794 305924
rect 284938 305872 284944 305924
rect 284996 305912 285002 305924
rect 292666 305912 292672 305924
rect 284996 305884 292672 305912
rect 284996 305872 285002 305884
rect 292666 305872 292672 305884
rect 292724 305872 292730 305924
rect 355134 305872 355140 305924
rect 355192 305912 355198 305924
rect 371786 305912 371792 305924
rect 355192 305884 371792 305912
rect 355192 305872 355198 305884
rect 371786 305872 371792 305884
rect 371844 305872 371850 305924
rect 213822 305804 213828 305856
rect 213880 305844 213886 305856
rect 213880 305816 273254 305844
rect 213880 305804 213886 305816
rect 170398 305736 170404 305788
rect 170456 305776 170462 305788
rect 255130 305776 255136 305788
rect 170456 305748 255136 305776
rect 170456 305736 170462 305748
rect 255130 305736 255136 305748
rect 255188 305736 255194 305788
rect 256970 305736 256976 305788
rect 257028 305776 257034 305788
rect 257614 305776 257620 305788
rect 257028 305748 257620 305776
rect 257028 305736 257034 305748
rect 257614 305736 257620 305748
rect 257672 305736 257678 305788
rect 258258 305736 258264 305788
rect 258316 305776 258322 305788
rect 258810 305776 258816 305788
rect 258316 305748 258816 305776
rect 258316 305736 258322 305748
rect 258810 305736 258816 305748
rect 258868 305736 258874 305788
rect 261018 305736 261024 305788
rect 261076 305776 261082 305788
rect 261478 305776 261484 305788
rect 261076 305748 261484 305776
rect 261076 305736 261082 305748
rect 261478 305736 261484 305748
rect 261536 305736 261542 305788
rect 262306 305736 262312 305788
rect 262364 305776 262370 305788
rect 263134 305776 263140 305788
rect 262364 305748 263140 305776
rect 262364 305736 262370 305748
rect 263134 305736 263140 305748
rect 263192 305736 263198 305788
rect 263962 305736 263968 305788
rect 264020 305776 264026 305788
rect 264698 305776 264704 305788
rect 264020 305748 264704 305776
rect 264020 305736 264026 305748
rect 264698 305736 264704 305748
rect 264756 305736 264762 305788
rect 266814 305736 266820 305788
rect 266872 305776 266878 305788
rect 267550 305776 267556 305788
rect 266872 305748 267556 305776
rect 266872 305736 266878 305748
rect 267550 305736 267556 305748
rect 267608 305736 267614 305788
rect 270770 305736 270776 305788
rect 270828 305776 270834 305788
rect 271414 305776 271420 305788
rect 270828 305748 271420 305776
rect 270828 305736 270834 305748
rect 271414 305736 271420 305748
rect 271472 305736 271478 305788
rect 273226 305776 273254 305816
rect 277578 305804 277584 305856
rect 277636 305844 277642 305856
rect 278222 305844 278228 305856
rect 277636 305816 278228 305844
rect 277636 305804 277642 305816
rect 278222 305804 278228 305816
rect 278280 305804 278286 305856
rect 278866 305804 278872 305856
rect 278924 305844 278930 305856
rect 279602 305844 279608 305856
rect 278924 305816 279608 305844
rect 278924 305804 278930 305816
rect 279602 305804 279608 305816
rect 279660 305804 279666 305856
rect 280430 305804 280436 305856
rect 280488 305844 280494 305856
rect 281074 305844 281080 305856
rect 280488 305816 281080 305844
rect 280488 305804 280494 305816
rect 281074 305804 281080 305816
rect 281132 305804 281138 305856
rect 281810 305804 281816 305856
rect 281868 305844 281874 305856
rect 282270 305844 282276 305856
rect 281868 305816 282276 305844
rect 281868 305804 281874 305816
rect 282270 305804 282276 305816
rect 282328 305804 282334 305856
rect 294690 305844 294696 305856
rect 283116 305816 294696 305844
rect 283116 305776 283144 305816
rect 294690 305804 294696 305816
rect 294748 305804 294754 305856
rect 343910 305804 343916 305856
rect 343968 305844 343974 305856
rect 344646 305844 344652 305856
rect 343968 305816 344652 305844
rect 343968 305804 343974 305816
rect 344646 305804 344652 305816
rect 344704 305804 344710 305856
rect 353570 305804 353576 305856
rect 353628 305844 353634 305856
rect 359826 305844 359832 305856
rect 353628 305816 359832 305844
rect 353628 305804 353634 305816
rect 359826 305804 359832 305816
rect 359884 305804 359890 305856
rect 359918 305804 359924 305856
rect 359976 305844 359982 305856
rect 369118 305844 369124 305856
rect 359976 305816 369124 305844
rect 359976 305804 359982 305816
rect 369118 305804 369124 305816
rect 369176 305804 369182 305856
rect 273226 305748 283144 305776
rect 284846 305736 284852 305788
rect 284904 305776 284910 305788
rect 292390 305776 292396 305788
rect 284904 305748 292396 305776
rect 284904 305736 284910 305748
rect 292390 305736 292396 305748
rect 292448 305736 292454 305788
rect 354398 305736 354404 305788
rect 354456 305776 354462 305788
rect 371694 305776 371700 305788
rect 354456 305748 371700 305776
rect 354456 305736 354462 305748
rect 371694 305736 371700 305748
rect 371752 305736 371758 305788
rect 195974 305668 195980 305720
rect 196032 305708 196038 305720
rect 284294 305708 284300 305720
rect 196032 305680 284300 305708
rect 196032 305668 196038 305680
rect 284294 305668 284300 305680
rect 284352 305668 284358 305720
rect 287422 305668 287428 305720
rect 287480 305708 287486 305720
rect 287790 305708 287796 305720
rect 287480 305680 287796 305708
rect 287480 305668 287486 305680
rect 287790 305668 287796 305680
rect 287848 305668 287854 305720
rect 293034 305668 293040 305720
rect 293092 305708 293098 305720
rect 293862 305708 293868 305720
rect 293092 305680 293868 305708
rect 293092 305668 293098 305680
rect 293862 305668 293868 305680
rect 293920 305668 293926 305720
rect 351178 305668 351184 305720
rect 351236 305708 351242 305720
rect 359642 305708 359648 305720
rect 351236 305680 359648 305708
rect 351236 305668 351242 305680
rect 359642 305668 359648 305680
rect 359700 305668 359706 305720
rect 359734 305668 359740 305720
rect 359792 305708 359798 305720
rect 370222 305708 370228 305720
rect 359792 305680 370228 305708
rect 359792 305668 359798 305680
rect 370222 305668 370228 305680
rect 370280 305668 370286 305720
rect 178034 305600 178040 305652
rect 178092 305640 178098 305652
rect 280062 305640 280068 305652
rect 178092 305612 280068 305640
rect 178092 305600 178098 305612
rect 280062 305600 280068 305612
rect 280120 305600 280126 305652
rect 280246 305600 280252 305652
rect 280304 305640 280310 305652
rect 280890 305640 280896 305652
rect 280304 305612 280896 305640
rect 280304 305600 280310 305612
rect 280890 305600 280896 305612
rect 280948 305600 280954 305652
rect 281718 305600 281724 305652
rect 281776 305640 281782 305652
rect 282822 305640 282828 305652
rect 281776 305612 282828 305640
rect 281776 305600 281782 305612
rect 282822 305600 282828 305612
rect 282880 305600 282886 305652
rect 283190 305600 283196 305652
rect 283248 305640 283254 305652
rect 283926 305640 283932 305652
rect 283248 305612 283932 305640
rect 283248 305600 283254 305612
rect 283926 305600 283932 305612
rect 283984 305600 283990 305652
rect 298186 305600 298192 305652
rect 298244 305640 298250 305652
rect 299198 305640 299204 305652
rect 298244 305612 299204 305640
rect 298244 305600 298250 305612
rect 299198 305600 299204 305612
rect 299256 305600 299262 305652
rect 347130 305600 347136 305652
rect 347188 305640 347194 305652
rect 370406 305640 370412 305652
rect 347188 305612 370412 305640
rect 347188 305600 347194 305612
rect 370406 305600 370412 305612
rect 370464 305600 370470 305652
rect 218974 305532 218980 305584
rect 219032 305572 219038 305584
rect 290642 305572 290648 305584
rect 219032 305544 290648 305572
rect 219032 305532 219038 305544
rect 290642 305532 290648 305544
rect 290700 305532 290706 305584
rect 352282 305532 352288 305584
rect 352340 305572 352346 305584
rect 359918 305572 359924 305584
rect 352340 305544 359924 305572
rect 352340 305532 352346 305544
rect 359918 305532 359924 305544
rect 359976 305532 359982 305584
rect 360010 305532 360016 305584
rect 360068 305572 360074 305584
rect 363598 305572 363604 305584
rect 360068 305544 363604 305572
rect 360068 305532 360074 305544
rect 363598 305532 363604 305544
rect 363656 305532 363662 305584
rect 218882 305464 218888 305516
rect 218940 305504 218946 305516
rect 289538 305504 289544 305516
rect 218940 305476 289544 305504
rect 218940 305464 218946 305476
rect 289538 305464 289544 305476
rect 289596 305464 289602 305516
rect 309318 305464 309324 305516
rect 309376 305504 309382 305516
rect 310146 305504 310152 305516
rect 309376 305476 310152 305504
rect 309376 305464 309382 305476
rect 310146 305464 310152 305476
rect 310204 305464 310210 305516
rect 355778 305464 355784 305516
rect 355836 305504 355842 305516
rect 365070 305504 365076 305516
rect 355836 305476 365076 305504
rect 355836 305464 355842 305476
rect 365070 305464 365076 305476
rect 365128 305464 365134 305516
rect 172146 305396 172152 305448
rect 172204 305436 172210 305448
rect 235166 305436 235172 305448
rect 172204 305408 235172 305436
rect 172204 305396 172210 305408
rect 235166 305396 235172 305408
rect 235224 305396 235230 305448
rect 235902 305396 235908 305448
rect 235960 305436 235966 305448
rect 236638 305436 236644 305448
rect 235960 305408 236644 305436
rect 235960 305396 235966 305408
rect 236638 305396 236644 305408
rect 236696 305396 236702 305448
rect 247678 305396 247684 305448
rect 247736 305436 247742 305448
rect 247954 305436 247960 305448
rect 247736 305408 247960 305436
rect 247736 305396 247742 305408
rect 247954 305396 247960 305408
rect 248012 305396 248018 305448
rect 256878 305396 256884 305448
rect 256936 305436 256942 305448
rect 257430 305436 257436 305448
rect 256936 305408 257436 305436
rect 256936 305396 256942 305408
rect 257430 305396 257436 305408
rect 257488 305396 257494 305448
rect 261110 305396 261116 305448
rect 261168 305436 261174 305448
rect 262030 305436 262036 305448
rect 261168 305408 262036 305436
rect 261168 305396 261174 305408
rect 262030 305396 262036 305408
rect 262088 305396 262094 305448
rect 266446 305396 266452 305448
rect 266504 305436 266510 305448
rect 267182 305436 267188 305448
rect 266504 305408 267188 305436
rect 266504 305396 266510 305408
rect 267182 305396 267188 305408
rect 267240 305396 267246 305448
rect 271046 305396 271052 305448
rect 271104 305436 271110 305448
rect 271782 305436 271788 305448
rect 271104 305408 271788 305436
rect 271104 305396 271110 305408
rect 271782 305396 271788 305408
rect 271840 305396 271846 305448
rect 276382 305396 276388 305448
rect 276440 305436 276446 305448
rect 276934 305436 276940 305448
rect 276440 305408 276940 305436
rect 276440 305396 276446 305408
rect 276934 305396 276940 305408
rect 276992 305396 276998 305448
rect 280154 305396 280160 305448
rect 280212 305436 280218 305448
rect 280522 305436 280528 305448
rect 280212 305408 280528 305436
rect 280212 305396 280218 305408
rect 280522 305396 280528 305408
rect 280580 305396 280586 305448
rect 282730 305396 282736 305448
rect 282788 305436 282794 305448
rect 284938 305436 284944 305448
rect 282788 305408 284944 305436
rect 282788 305396 282794 305408
rect 284938 305396 284944 305408
rect 284996 305396 285002 305448
rect 349430 305396 349436 305448
rect 349488 305436 349494 305448
rect 349488 305408 350534 305436
rect 349488 305396 349494 305408
rect 97442 305328 97448 305380
rect 97500 305328 97506 305380
rect 256694 305328 256700 305380
rect 256752 305368 256758 305380
rect 257338 305368 257344 305380
rect 256752 305340 257344 305368
rect 256752 305328 256758 305340
rect 257338 305328 257344 305340
rect 257396 305328 257402 305380
rect 282362 305328 282368 305380
rect 282420 305368 282426 305380
rect 284846 305368 284852 305380
rect 282420 305340 284852 305368
rect 282420 305328 282426 305340
rect 284846 305328 284852 305340
rect 284904 305328 284910 305380
rect 350506 305368 350534 305408
rect 359182 305396 359188 305448
rect 359240 305436 359246 305448
rect 360102 305436 360108 305448
rect 359240 305408 360108 305436
rect 359240 305396 359246 305408
rect 360102 305396 360108 305408
rect 360160 305396 360166 305448
rect 359550 305368 359556 305380
rect 350506 305340 359556 305368
rect 359550 305328 359556 305340
rect 359608 305328 359614 305380
rect 97460 305176 97488 305328
rect 352650 305260 352656 305312
rect 352708 305300 352714 305312
rect 360010 305300 360016 305312
rect 352708 305272 360016 305300
rect 352708 305260 352714 305272
rect 360010 305260 360016 305272
rect 360068 305260 360074 305312
rect 343634 305192 343640 305244
rect 343692 305232 343698 305244
rect 344830 305232 344836 305244
rect 343692 305204 344836 305232
rect 343692 305192 343698 305204
rect 344830 305192 344836 305204
rect 344888 305192 344894 305244
rect 351730 305192 351736 305244
rect 351788 305232 351794 305244
rect 359734 305232 359740 305244
rect 351788 305204 359740 305232
rect 351788 305192 351794 305204
rect 359734 305192 359740 305204
rect 359792 305192 359798 305244
rect 97442 305124 97448 305176
rect 97500 305124 97506 305176
rect 276014 305056 276020 305108
rect 276072 305096 276078 305108
rect 277118 305096 277124 305108
rect 276072 305068 277124 305096
rect 276072 305056 276078 305068
rect 277118 305056 277124 305068
rect 277176 305056 277182 305108
rect 97626 304920 97632 304972
rect 97684 304960 97690 304972
rect 97902 304960 97908 304972
rect 97684 304932 97908 304960
rect 97684 304920 97690 304932
rect 97902 304920 97908 304932
rect 97960 304920 97966 304972
rect 172330 304920 172336 304972
rect 172388 304960 172394 304972
rect 245194 304960 245200 304972
rect 172388 304932 245200 304960
rect 172388 304920 172394 304932
rect 245194 304920 245200 304932
rect 245252 304920 245258 304972
rect 294138 304852 294144 304904
rect 294196 304892 294202 304904
rect 294322 304892 294328 304904
rect 294196 304864 294328 304892
rect 294196 304852 294202 304864
rect 294322 304852 294328 304864
rect 294380 304852 294386 304904
rect 294322 304716 294328 304768
rect 294380 304756 294386 304768
rect 295058 304756 295064 304768
rect 294380 304728 295064 304756
rect 294380 304716 294386 304728
rect 295058 304716 295064 304728
rect 295116 304716 295122 304768
rect 258350 304648 258356 304700
rect 258408 304688 258414 304700
rect 259178 304688 259184 304700
rect 258408 304660 259184 304688
rect 258408 304648 258414 304660
rect 259178 304648 259184 304660
rect 259236 304648 259242 304700
rect 264974 304648 264980 304700
rect 265032 304688 265038 304700
rect 265894 304688 265900 304700
rect 265032 304660 265900 304688
rect 265032 304648 265038 304660
rect 265894 304648 265900 304660
rect 265952 304648 265958 304700
rect 169938 304580 169944 304632
rect 169996 304620 170002 304632
rect 237190 304620 237196 304632
rect 169996 304592 237196 304620
rect 169996 304580 170002 304592
rect 237190 304580 237196 304592
rect 237248 304580 237254 304632
rect 274634 304580 274640 304632
rect 274692 304620 274698 304632
rect 275738 304620 275744 304632
rect 274692 304592 275744 304620
rect 274692 304580 274698 304592
rect 275738 304580 275744 304592
rect 275796 304580 275802 304632
rect 169846 304512 169852 304564
rect 169904 304552 169910 304564
rect 243170 304552 243176 304564
rect 169904 304524 243176 304552
rect 169904 304512 169910 304524
rect 243170 304512 243176 304524
rect 243228 304512 243234 304564
rect 290182 304512 290188 304564
rect 290240 304552 290246 304564
rect 291010 304552 291016 304564
rect 290240 304524 291016 304552
rect 290240 304512 290246 304524
rect 291010 304512 291016 304524
rect 291068 304512 291074 304564
rect 172238 304444 172244 304496
rect 172296 304484 172302 304496
rect 246022 304484 246028 304496
rect 172296 304456 246028 304484
rect 172296 304444 172302 304456
rect 246022 304444 246028 304456
rect 246080 304444 246086 304496
rect 324222 304444 324228 304496
rect 324280 304484 324286 304496
rect 440878 304484 440884 304496
rect 324280 304456 440884 304484
rect 324280 304444 324286 304456
rect 440878 304444 440884 304456
rect 440936 304444 440942 304496
rect 171410 304376 171416 304428
rect 171468 304416 171474 304428
rect 249426 304416 249432 304428
rect 171468 304388 249432 304416
rect 171468 304376 171474 304388
rect 249426 304376 249432 304388
rect 249484 304376 249490 304428
rect 250346 304376 250352 304428
rect 250404 304416 250410 304428
rect 250806 304416 250812 304428
rect 250404 304388 250812 304416
rect 250404 304376 250410 304388
rect 250806 304376 250812 304388
rect 250864 304376 250870 304428
rect 299934 304376 299940 304428
rect 299992 304416 299998 304428
rect 300762 304416 300768 304428
rect 299992 304388 300768 304416
rect 299992 304376 299998 304388
rect 300762 304376 300768 304388
rect 300820 304376 300826 304428
rect 326430 304376 326436 304428
rect 326488 304416 326494 304428
rect 452654 304416 452660 304428
rect 326488 304388 452660 304416
rect 326488 304376 326494 304388
rect 452654 304376 452660 304388
rect 452712 304376 452718 304428
rect 207014 304308 207020 304360
rect 207072 304348 207078 304360
rect 285674 304348 285680 304360
rect 207072 304320 285680 304348
rect 207072 304308 207078 304320
rect 285674 304308 285680 304320
rect 285732 304308 285738 304360
rect 331766 304308 331772 304360
rect 331824 304348 331830 304360
rect 485038 304348 485044 304360
rect 331824 304320 485044 304348
rect 331824 304308 331830 304320
rect 485038 304308 485044 304320
rect 485096 304308 485102 304360
rect 189074 304240 189080 304292
rect 189132 304280 189138 304292
rect 283098 304280 283104 304292
rect 189132 304252 283104 304280
rect 189132 304240 189138 304252
rect 283098 304240 283104 304252
rect 283156 304240 283162 304292
rect 303890 304240 303896 304292
rect 303948 304280 303954 304292
rect 304166 304280 304172 304292
rect 303948 304252 304172 304280
rect 303948 304240 303954 304252
rect 304166 304240 304172 304252
rect 304224 304240 304230 304292
rect 335906 304240 335912 304292
rect 335964 304280 335970 304292
rect 514018 304280 514024 304292
rect 335964 304252 514024 304280
rect 335964 304240 335970 304252
rect 514018 304240 514024 304252
rect 514076 304240 514082 304292
rect 252738 304172 252744 304224
rect 252796 304212 252802 304224
rect 253106 304212 253112 304224
rect 252796 304184 253112 304212
rect 252796 304172 252802 304184
rect 253106 304172 253112 304184
rect 253164 304172 253170 304224
rect 262490 304172 262496 304224
rect 262548 304212 262554 304224
rect 262766 304212 262772 304224
rect 262548 304184 262772 304212
rect 262548 304172 262554 304184
rect 262766 304172 262772 304184
rect 262824 304172 262830 304224
rect 295334 304172 295340 304224
rect 295392 304212 295398 304224
rect 296162 304212 296168 304224
rect 295392 304184 296168 304212
rect 295392 304172 295398 304184
rect 296162 304172 296168 304184
rect 296220 304172 296226 304224
rect 252922 303832 252928 303884
rect 252980 303872 252986 303884
rect 253842 303872 253848 303884
rect 252980 303844 253848 303872
rect 252980 303832 252986 303844
rect 253842 303832 253848 303844
rect 253900 303832 253906 303884
rect 269298 303696 269304 303748
rect 269356 303736 269362 303748
rect 270402 303736 270408 303748
rect 269356 303708 270408 303736
rect 269356 303696 269362 303708
rect 270402 303696 270408 303708
rect 270460 303696 270466 303748
rect 265158 303628 265164 303680
rect 265216 303668 265222 303680
rect 266262 303668 266268 303680
rect 265216 303640 266268 303668
rect 265216 303628 265222 303640
rect 266262 303628 266268 303640
rect 266320 303628 266326 303680
rect 217962 303560 217968 303612
rect 218020 303600 218026 303612
rect 292850 303600 292856 303612
rect 218020 303572 292856 303600
rect 218020 303560 218026 303572
rect 292850 303560 292856 303572
rect 292908 303560 292914 303612
rect 355870 303560 355876 303612
rect 355928 303600 355934 303612
rect 372062 303600 372068 303612
rect 355928 303572 372068 303600
rect 355928 303560 355934 303572
rect 372062 303560 372068 303572
rect 372120 303560 372126 303612
rect 216398 303492 216404 303544
rect 216456 303532 216462 303544
rect 291378 303532 291384 303544
rect 216456 303504 291384 303532
rect 216456 303492 216462 303504
rect 291378 303492 291384 303504
rect 291436 303492 291442 303544
rect 347958 303492 347964 303544
rect 348016 303532 348022 303544
rect 367922 303532 367928 303544
rect 348016 303504 367928 303532
rect 348016 303492 348022 303504
rect 367922 303492 367928 303504
rect 367980 303492 367986 303544
rect 214834 303424 214840 303476
rect 214892 303464 214898 303476
rect 290826 303464 290832 303476
rect 214892 303436 290832 303464
rect 214892 303424 214898 303436
rect 290826 303424 290832 303436
rect 290884 303424 290890 303476
rect 352466 303424 352472 303476
rect 352524 303464 352530 303476
rect 372798 303464 372804 303476
rect 352524 303436 372804 303464
rect 352524 303424 352530 303436
rect 372798 303424 372804 303436
rect 372856 303424 372862 303476
rect 212442 303356 212448 303408
rect 212500 303396 212506 303408
rect 289354 303396 289360 303408
rect 212500 303368 289360 303396
rect 212500 303356 212506 303368
rect 289354 303356 289360 303368
rect 289412 303356 289418 303408
rect 350166 303356 350172 303408
rect 350224 303396 350230 303408
rect 370590 303396 370596 303408
rect 350224 303368 370596 303396
rect 350224 303356 350230 303368
rect 370590 303356 370596 303368
rect 370648 303356 370654 303408
rect 219250 303288 219256 303340
rect 219308 303328 219314 303340
rect 295426 303328 295432 303340
rect 219308 303300 295432 303328
rect 219308 303288 219314 303300
rect 295426 303288 295432 303300
rect 295484 303288 295490 303340
rect 352834 303288 352840 303340
rect 352892 303328 352898 303340
rect 374178 303328 374184 303340
rect 352892 303300 374184 303328
rect 352892 303288 352898 303300
rect 374178 303288 374184 303300
rect 374236 303288 374242 303340
rect 216214 303220 216220 303272
rect 216272 303260 216278 303272
rect 292574 303260 292580 303272
rect 216272 303232 292580 303260
rect 216272 303220 216278 303232
rect 292574 303220 292580 303232
rect 292632 303220 292638 303272
rect 351914 303220 351920 303272
rect 351972 303260 351978 303272
rect 374362 303260 374368 303272
rect 351972 303232 374368 303260
rect 351972 303220 351978 303232
rect 374362 303220 374368 303232
rect 374420 303220 374426 303272
rect 214558 303152 214564 303204
rect 214616 303192 214622 303204
rect 292022 303192 292028 303204
rect 214616 303164 292028 303192
rect 214616 303152 214622 303164
rect 292022 303152 292028 303164
rect 292080 303152 292086 303204
rect 299842 303152 299848 303204
rect 299900 303192 299906 303204
rect 300578 303192 300584 303204
rect 299900 303164 300584 303192
rect 299900 303152 299906 303164
rect 300578 303152 300584 303164
rect 300636 303152 300642 303204
rect 348878 303152 348884 303204
rect 348936 303192 348942 303204
rect 372982 303192 372988 303204
rect 348936 303164 372988 303192
rect 348936 303152 348942 303164
rect 372982 303152 372988 303164
rect 373040 303152 373046 303204
rect 212074 303084 212080 303136
rect 212132 303124 212138 303136
rect 289906 303124 289912 303136
rect 212132 303096 289912 303124
rect 212132 303084 212138 303096
rect 289906 303084 289912 303096
rect 289964 303084 289970 303136
rect 349614 303084 349620 303136
rect 349672 303124 349678 303136
rect 374270 303124 374276 303136
rect 349672 303096 374276 303124
rect 349672 303084 349678 303096
rect 374270 303084 374276 303096
rect 374328 303084 374334 303136
rect 169754 303016 169760 303068
rect 169812 303056 169818 303068
rect 251542 303056 251548 303068
rect 169812 303028 251548 303056
rect 169812 303016 169818 303028
rect 251542 303016 251548 303028
rect 251600 303016 251606 303068
rect 301130 303016 301136 303068
rect 301188 303056 301194 303068
rect 363690 303056 363696 303068
rect 301188 303028 363696 303056
rect 301188 303016 301194 303028
rect 363690 303016 363696 303028
rect 363748 303016 363754 303068
rect 213638 302948 213644 303000
rect 213696 302988 213702 303000
rect 294046 302988 294052 303000
rect 213696 302960 294052 302988
rect 213696 302948 213702 302960
rect 294046 302948 294052 302960
rect 294104 302948 294110 303000
rect 298370 302948 298376 303000
rect 298428 302988 298434 303000
rect 367094 302988 367100 303000
rect 298428 302960 367100 302988
rect 298428 302948 298434 302960
rect 367094 302948 367100 302960
rect 367152 302948 367158 303000
rect 184934 302880 184940 302932
rect 184992 302920 184998 302932
rect 282638 302920 282644 302932
rect 184992 302892 282644 302920
rect 184992 302880 184998 302892
rect 282638 302880 282644 302892
rect 282696 302880 282702 302932
rect 298830 302880 298836 302932
rect 298888 302920 298894 302932
rect 367830 302920 367836 302932
rect 298888 302892 367836 302920
rect 298888 302880 298894 302892
rect 367830 302880 367836 302892
rect 367888 302880 367894 302932
rect 214650 302812 214656 302864
rect 214708 302852 214714 302864
rect 289722 302852 289728 302864
rect 214708 302824 289728 302852
rect 214708 302812 214714 302824
rect 289722 302812 289728 302824
rect 289780 302812 289786 302864
rect 350718 302812 350724 302864
rect 350776 302852 350782 302864
rect 366450 302852 366456 302864
rect 350776 302824 366456 302852
rect 350776 302812 350782 302824
rect 366450 302812 366456 302824
rect 366508 302812 366514 302864
rect 216122 302744 216128 302796
rect 216180 302784 216186 302796
rect 290274 302784 290280 302796
rect 216180 302756 290280 302784
rect 216180 302744 216186 302756
rect 290274 302744 290280 302756
rect 290332 302744 290338 302796
rect 341150 302744 341156 302796
rect 341208 302784 341214 302796
rect 342162 302784 342168 302796
rect 341208 302756 342168 302784
rect 341208 302744 341214 302756
rect 342162 302744 342168 302756
rect 342220 302744 342226 302796
rect 356606 302744 356612 302796
rect 356664 302784 356670 302796
rect 370682 302784 370688 302796
rect 356664 302756 370688 302784
rect 356664 302744 356670 302756
rect 370682 302744 370688 302756
rect 370740 302744 370746 302796
rect 214742 302676 214748 302728
rect 214800 302716 214806 302728
rect 288158 302716 288164 302728
rect 214800 302688 288164 302716
rect 214800 302676 214806 302688
rect 288158 302676 288164 302688
rect 288216 302676 288222 302728
rect 351362 302676 351368 302728
rect 351420 302716 351426 302728
rect 362310 302716 362316 302728
rect 351420 302688 362316 302716
rect 351420 302676 351426 302688
rect 362310 302676 362316 302688
rect 362368 302676 362374 302728
rect 269574 302472 269580 302524
rect 269632 302512 269638 302524
rect 270034 302512 270040 302524
rect 269632 302484 270040 302512
rect 269632 302472 269638 302484
rect 270034 302472 270040 302484
rect 270092 302472 270098 302524
rect 334250 302472 334256 302524
rect 334308 302512 334314 302524
rect 334710 302512 334716 302524
rect 334308 302484 334716 302512
rect 334308 302472 334314 302484
rect 334710 302472 334716 302484
rect 334768 302472 334774 302524
rect 236454 302308 236460 302320
rect 236196 302280 236460 302308
rect 236196 302252 236224 302280
rect 236454 302268 236460 302280
rect 236512 302268 236518 302320
rect 236178 302200 236184 302252
rect 236236 302200 236242 302252
rect 172422 302132 172428 302184
rect 172480 302172 172486 302184
rect 240134 302172 240140 302184
rect 172480 302144 240140 302172
rect 172480 302132 172486 302144
rect 240134 302132 240140 302144
rect 240192 302132 240198 302184
rect 210970 301724 210976 301776
rect 211028 301764 211034 301776
rect 295334 301764 295340 301776
rect 211028 301736 295340 301764
rect 211028 301724 211034 301736
rect 295334 301724 295340 301736
rect 295392 301724 295398 301776
rect 212166 301656 212172 301708
rect 212224 301696 212230 301708
rect 296806 301696 296812 301708
rect 212224 301668 296812 301696
rect 212224 301656 212230 301668
rect 296806 301656 296812 301668
rect 296864 301656 296870 301708
rect 312262 301656 312268 301708
rect 312320 301696 312326 301708
rect 373994 301696 374000 301708
rect 312320 301668 374000 301696
rect 312320 301656 312326 301668
rect 373994 301656 374000 301668
rect 374052 301656 374058 301708
rect 211890 301588 211896 301640
rect 211948 301628 211954 301640
rect 347958 301628 347964 301640
rect 211948 301600 347964 301628
rect 211948 301588 211954 301600
rect 347958 301588 347964 301600
rect 348016 301588 348022 301640
rect 358814 301588 358820 301640
rect 358872 301628 358878 301640
rect 358998 301628 359004 301640
rect 358872 301600 359004 301628
rect 358872 301588 358878 301600
rect 358998 301588 359004 301600
rect 359056 301588 359062 301640
rect 171778 301520 171784 301572
rect 171836 301560 171842 301572
rect 257338 301560 257344 301572
rect 171836 301532 257344 301560
rect 171836 301520 171842 301532
rect 257338 301520 257344 301532
rect 257396 301520 257402 301572
rect 331582 301520 331588 301572
rect 331640 301560 331646 301572
rect 494054 301560 494060 301572
rect 331640 301532 494060 301560
rect 331640 301520 331646 301532
rect 494054 301520 494060 301532
rect 494112 301520 494118 301572
rect 193214 301452 193220 301504
rect 193272 301492 193278 301504
rect 282914 301492 282920 301504
rect 193272 301464 282920 301492
rect 193272 301452 193278 301464
rect 282914 301452 282920 301464
rect 282972 301452 282978 301504
rect 338666 301452 338672 301504
rect 338724 301492 338730 301504
rect 529934 301492 529940 301504
rect 338724 301464 529940 301492
rect 338724 301452 338730 301464
rect 529934 301452 529940 301464
rect 529992 301452 529998 301504
rect 276290 300840 276296 300892
rect 276348 300880 276354 300892
rect 276566 300880 276572 300892
rect 276348 300852 276572 300880
rect 276348 300840 276354 300852
rect 276566 300840 276572 300852
rect 276624 300840 276630 300892
rect 97442 300772 97448 300824
rect 97500 300812 97506 300824
rect 249978 300812 249984 300824
rect 97500 300784 249984 300812
rect 97500 300772 97506 300784
rect 249978 300772 249984 300784
rect 250036 300772 250042 300824
rect 99098 300704 99104 300756
rect 99156 300744 99162 300756
rect 251358 300744 251364 300756
rect 99156 300716 251364 300744
rect 99156 300704 99162 300716
rect 251358 300704 251364 300716
rect 251416 300704 251422 300756
rect 97074 300636 97080 300688
rect 97132 300676 97138 300688
rect 245746 300676 245752 300688
rect 97132 300648 245752 300676
rect 97132 300636 97138 300648
rect 245746 300636 245752 300648
rect 245804 300636 245810 300688
rect 313826 300636 313832 300688
rect 313884 300676 313890 300688
rect 376754 300676 376760 300688
rect 313884 300648 376760 300676
rect 313884 300636 313890 300648
rect 376754 300636 376760 300648
rect 376812 300636 376818 300688
rect 97810 300568 97816 300620
rect 97868 300608 97874 300620
rect 246206 300608 246212 300620
rect 97868 300580 246212 300608
rect 97868 300568 97874 300580
rect 246206 300568 246212 300580
rect 246264 300568 246270 300620
rect 298278 300568 298284 300620
rect 298336 300608 298342 300620
rect 365162 300608 365168 300620
rect 298336 300580 365168 300608
rect 298336 300568 298342 300580
rect 365162 300568 365168 300580
rect 365220 300568 365226 300620
rect 99374 300500 99380 300552
rect 99432 300540 99438 300552
rect 247126 300540 247132 300552
rect 99432 300512 247132 300540
rect 99432 300500 99438 300512
rect 247126 300500 247132 300512
rect 247184 300500 247190 300552
rect 299842 300500 299848 300552
rect 299900 300540 299906 300552
rect 369210 300540 369216 300552
rect 299900 300512 369216 300540
rect 299900 300500 299906 300512
rect 369210 300500 369216 300512
rect 369268 300500 369274 300552
rect 97902 300432 97908 300484
rect 97960 300472 97966 300484
rect 242802 300472 242808 300484
rect 97960 300444 242808 300472
rect 97960 300432 97966 300444
rect 242802 300432 242808 300444
rect 242860 300432 242866 300484
rect 301130 300432 301136 300484
rect 301188 300472 301194 300484
rect 370498 300472 370504 300484
rect 301188 300444 370504 300472
rect 301188 300432 301194 300444
rect 370498 300432 370504 300444
rect 370556 300432 370562 300484
rect 98914 300364 98920 300416
rect 98972 300404 98978 300416
rect 243354 300404 243360 300416
rect 98972 300376 243360 300404
rect 98972 300364 98978 300376
rect 243354 300364 243360 300376
rect 243412 300364 243418 300416
rect 299934 300364 299940 300416
rect 299992 300404 299998 300416
rect 372890 300404 372896 300416
rect 299992 300376 372896 300404
rect 299992 300364 299998 300376
rect 372890 300364 372896 300376
rect 372948 300364 372954 300416
rect 97718 300296 97724 300348
rect 97776 300336 97782 300348
rect 242710 300336 242716 300348
rect 97776 300308 242716 300336
rect 97776 300296 97782 300308
rect 242710 300296 242716 300308
rect 242768 300296 242774 300348
rect 320818 300296 320824 300348
rect 320876 300336 320882 300348
rect 422294 300336 422300 300348
rect 320876 300308 422300 300336
rect 320876 300296 320882 300308
rect 422294 300296 422300 300308
rect 422352 300296 422358 300348
rect 99834 300228 99840 300280
rect 99892 300268 99898 300280
rect 240410 300268 240416 300280
rect 99892 300240 240416 300268
rect 99892 300228 99898 300240
rect 240410 300228 240416 300240
rect 240468 300228 240474 300280
rect 333146 300228 333152 300280
rect 333204 300268 333210 300280
rect 498286 300268 498292 300280
rect 333204 300240 498292 300268
rect 333204 300228 333210 300240
rect 498286 300228 498292 300240
rect 498344 300228 498350 300280
rect 99466 300160 99472 300212
rect 99524 300200 99530 300212
rect 241054 300200 241060 300212
rect 99524 300172 241060 300200
rect 99524 300160 99530 300172
rect 241054 300160 241060 300172
rect 241112 300160 241118 300212
rect 339862 300160 339868 300212
rect 339920 300200 339926 300212
rect 538858 300200 538864 300212
rect 339920 300172 538864 300200
rect 339920 300160 339926 300172
rect 538858 300160 538864 300172
rect 538916 300160 538922 300212
rect 97626 300092 97632 300144
rect 97684 300132 97690 300144
rect 237558 300132 237564 300144
rect 97684 300104 237564 300132
rect 97684 300092 97690 300104
rect 237558 300092 237564 300104
rect 237616 300092 237622 300144
rect 341518 300092 341524 300144
rect 341576 300132 341582 300144
rect 545758 300132 545764 300144
rect 341576 300104 545764 300132
rect 341576 300092 341582 300104
rect 545758 300092 545764 300104
rect 545816 300092 545822 300144
rect 98822 300024 98828 300076
rect 98880 300064 98886 300076
rect 233326 300064 233332 300076
rect 98880 300036 233332 300064
rect 98880 300024 98886 300036
rect 233326 300024 233332 300036
rect 233384 300024 233390 300076
rect 205634 299956 205640 300008
rect 205692 299996 205698 300008
rect 285766 299996 285772 300008
rect 205692 299968 285772 299996
rect 205692 299956 205698 299968
rect 285766 299956 285772 299968
rect 285824 299956 285830 300008
rect 213362 299888 213368 299940
rect 213420 299928 213426 299940
rect 290274 299928 290280 299940
rect 213420 299900 290280 299928
rect 213420 299888 213426 299900
rect 290274 299888 290280 299900
rect 290332 299888 290338 299940
rect 99006 299412 99012 299464
rect 99064 299452 99070 299464
rect 240502 299452 240508 299464
rect 99064 299424 240508 299452
rect 99064 299412 99070 299424
rect 240502 299412 240508 299424
rect 240560 299412 240566 299464
rect 98638 299344 98644 299396
rect 98696 299384 98702 299396
rect 240226 299384 240232 299396
rect 98696 299356 240232 299384
rect 98696 299344 98702 299356
rect 240226 299344 240232 299356
rect 240284 299344 240290 299396
rect 98546 299276 98552 299328
rect 98604 299316 98610 299328
rect 238938 299316 238944 299328
rect 98604 299288 238944 299316
rect 98604 299276 98610 299288
rect 238938 299276 238944 299288
rect 238996 299276 239002 299328
rect 104526 299208 104532 299260
rect 104584 299248 104590 299260
rect 234982 299248 234988 299260
rect 104584 299220 234988 299248
rect 104584 299208 104590 299220
rect 234982 299208 234988 299220
rect 235040 299208 235046 299260
rect 114830 299140 114836 299192
rect 114888 299180 114894 299192
rect 244458 299180 244464 299192
rect 114888 299152 244464 299180
rect 114888 299140 114894 299152
rect 244458 299140 244464 299152
rect 244516 299140 244522 299192
rect 119982 299072 119988 299124
rect 120040 299112 120046 299124
rect 247218 299112 247224 299124
rect 120040 299084 247224 299112
rect 120040 299072 120046 299084
rect 247218 299072 247224 299084
rect 247276 299072 247282 299124
rect 117406 299004 117412 299056
rect 117464 299044 117470 299056
rect 243078 299044 243084 299056
rect 117464 299016 243084 299044
rect 117464 299004 117470 299016
rect 243078 299004 243084 299016
rect 243136 299004 243142 299056
rect 130286 298936 130292 298988
rect 130344 298976 130350 298988
rect 250346 298976 250352 298988
rect 130344 298948 250352 298976
rect 130344 298936 130350 298948
rect 250346 298936 250352 298948
rect 250404 298936 250410 298988
rect 319346 298936 319352 298988
rect 319404 298976 319410 298988
rect 377398 298976 377404 298988
rect 319404 298948 377404 298976
rect 319404 298936 319410 298948
rect 377398 298936 377404 298948
rect 377456 298936 377462 298988
rect 125134 298868 125140 298920
rect 125192 298908 125198 298920
rect 238846 298908 238852 298920
rect 125192 298880 238852 298908
rect 125192 298868 125198 298880
rect 238846 298868 238852 298880
rect 238904 298868 238910 298920
rect 315114 298868 315120 298920
rect 315172 298908 315178 298920
rect 385034 298908 385040 298920
rect 315172 298880 385040 298908
rect 315172 298868 315178 298880
rect 385034 298868 385040 298880
rect 385092 298868 385098 298920
rect 140590 298800 140596 298852
rect 140648 298840 140654 298852
rect 250622 298840 250628 298852
rect 140648 298812 250628 298840
rect 140648 298800 140654 298812
rect 250622 298800 250628 298812
rect 250680 298800 250686 298852
rect 333054 298800 333060 298852
rect 333112 298840 333118 298852
rect 500218 298840 500224 298852
rect 333112 298812 500224 298840
rect 333112 298800 333118 298812
rect 500218 298800 500224 298812
rect 500276 298800 500282 298852
rect 156046 298732 156052 298784
rect 156104 298772 156110 298784
rect 251726 298772 251732 298784
rect 156104 298744 251732 298772
rect 156104 298732 156110 298744
rect 251726 298732 251732 298744
rect 251784 298732 251790 298784
rect 341426 298732 341432 298784
rect 341484 298772 341490 298784
rect 547966 298772 547972 298784
rect 341484 298744 547972 298772
rect 341484 298732 341490 298744
rect 547966 298732 547972 298744
rect 548024 298732 548030 298784
rect 145742 298664 145748 298716
rect 145800 298704 145806 298716
rect 236178 298704 236184 298716
rect 145800 298676 236184 298704
rect 145800 298664 145806 298676
rect 236178 298664 236184 298676
rect 236236 298664 236242 298716
rect 161198 298596 161204 298648
rect 161256 298636 161262 298648
rect 247770 298636 247776 298648
rect 161256 298608 247776 298636
rect 161256 298596 161262 298608
rect 247770 298596 247776 298608
rect 247828 298596 247834 298648
rect 163774 298528 163780 298580
rect 163832 298568 163838 298580
rect 234706 298568 234712 298580
rect 163832 298540 234712 298568
rect 163832 298528 163838 298540
rect 234706 298528 234712 298540
rect 234764 298528 234770 298580
rect 158622 298052 158628 298104
rect 158680 298092 158686 298104
rect 158680 298064 161474 298092
rect 158680 298052 158686 298064
rect 161446 298024 161474 298064
rect 166350 298052 166356 298104
rect 166408 298092 166414 298104
rect 170582 298092 170588 298104
rect 166408 298064 170588 298092
rect 166408 298052 166414 298064
rect 170582 298052 170588 298064
rect 170640 298052 170646 298104
rect 169846 298024 169852 298036
rect 161446 297996 169852 298024
rect 169846 297984 169852 297996
rect 169904 297984 169910 298036
rect 132862 297916 132868 297968
rect 132920 297956 132926 297968
rect 251450 297956 251456 297968
rect 132920 297928 251456 297956
rect 132920 297916 132926 297928
rect 251450 297916 251456 297928
rect 251508 297916 251514 297968
rect 122558 297848 122564 297900
rect 122616 297888 122622 297900
rect 237926 297888 237932 297900
rect 122616 297860 237932 297888
rect 122616 297848 122622 297860
rect 237926 297848 237932 297860
rect 237984 297848 237990 297900
rect 138014 297780 138020 297832
rect 138072 297820 138078 297832
rect 239122 297820 239128 297832
rect 138072 297792 239128 297820
rect 138072 297780 138078 297792
rect 239122 297780 239128 297792
rect 239180 297780 239186 297832
rect 148318 297712 148324 297764
rect 148376 297752 148382 297764
rect 236270 297752 236276 297764
rect 148376 297724 236276 297752
rect 148376 297712 148382 297724
rect 236270 297712 236276 297724
rect 236328 297712 236334 297764
rect 100018 297644 100024 297696
rect 100076 297684 100082 297696
rect 172238 297684 172244 297696
rect 100076 297656 172244 297684
rect 100076 297644 100082 297656
rect 172238 297644 172244 297656
rect 172296 297644 172302 297696
rect 214466 297644 214472 297696
rect 214524 297684 214530 297696
rect 294414 297684 294420 297696
rect 214524 297656 294420 297684
rect 214524 297644 214530 297656
rect 294414 297644 294420 297656
rect 294472 297644 294478 297696
rect 322198 297644 322204 297696
rect 322256 297684 322262 297696
rect 381538 297684 381544 297696
rect 322256 297656 381544 297684
rect 322256 297644 322262 297656
rect 381538 297644 381544 297656
rect 381596 297644 381602 297696
rect 101950 297576 101956 297628
rect 102008 297616 102014 297628
rect 171410 297616 171416 297628
rect 102008 297588 171416 297616
rect 102008 297576 102014 297588
rect 171410 297576 171416 297588
rect 171468 297576 171474 297628
rect 213730 297576 213736 297628
rect 213788 297616 213794 297628
rect 294230 297616 294236 297628
rect 213788 297588 294236 297616
rect 213788 297576 213794 297588
rect 294230 297576 294236 297588
rect 294288 297576 294294 297628
rect 319254 297576 319260 297628
rect 319312 297616 319318 297628
rect 412634 297616 412640 297628
rect 319312 297588 412640 297616
rect 319312 297576 319318 297588
rect 412634 297576 412640 297588
rect 412692 297576 412698 297628
rect 107102 297508 107108 297560
rect 107160 297548 107166 297560
rect 169938 297548 169944 297560
rect 107160 297520 169944 297548
rect 107160 297508 107166 297520
rect 169938 297508 169944 297520
rect 169996 297508 170002 297560
rect 213270 297508 213276 297560
rect 213328 297548 213334 297560
rect 346578 297548 346584 297560
rect 213328 297520 346584 297548
rect 213328 297508 213334 297520
rect 346578 297508 346584 297520
rect 346636 297508 346642 297560
rect 135438 297440 135444 297492
rect 135496 297480 135502 297492
rect 171686 297480 171692 297492
rect 135496 297452 171692 297480
rect 135496 297440 135502 297452
rect 171686 297440 171692 297452
rect 171744 297440 171750 297492
rect 210878 297440 210884 297492
rect 210936 297480 210942 297492
rect 293034 297480 293040 297492
rect 210936 297452 293040 297480
rect 210936 297440 210942 297452
rect 293034 297440 293040 297452
rect 293092 297440 293098 297492
rect 327626 297440 327632 297492
rect 327684 297480 327690 297492
rect 463694 297480 463700 297492
rect 327684 297452 463700 297480
rect 327684 297440 327690 297452
rect 463694 297440 463700 297452
rect 463752 297440 463758 297492
rect 143166 297372 143172 297424
rect 143224 297412 143230 297424
rect 143224 297384 161474 297412
rect 143224 297372 143230 297384
rect 161446 297344 161474 297384
rect 211706 297372 211712 297424
rect 211764 297412 211770 297424
rect 294138 297412 294144 297424
rect 211764 297384 294144 297412
rect 211764 297372 211770 297384
rect 294138 297372 294144 297384
rect 294196 297372 294202 297424
rect 342806 297372 342812 297424
rect 342864 297412 342870 297424
rect 557534 297412 557540 297424
rect 342864 297384 557540 297412
rect 342864 297372 342870 297384
rect 557534 297372 557540 297384
rect 557592 297372 557598 297424
rect 172146 297344 172152 297356
rect 161446 297316 172152 297344
rect 172146 297304 172152 297316
rect 172204 297304 172210 297356
rect 213454 297304 213460 297356
rect 213512 297344 213518 297356
rect 293126 297344 293132 297356
rect 213512 297316 293132 297344
rect 213512 297304 213518 297316
rect 293126 297304 293132 297316
rect 293184 297304 293190 297356
rect 215846 297236 215852 297288
rect 215904 297276 215910 297288
rect 295242 297276 295248 297288
rect 215904 297248 295248 297276
rect 215904 297236 215910 297248
rect 295242 297236 295248 297248
rect 295300 297236 295306 297288
rect 216030 297168 216036 297220
rect 216088 297208 216094 297220
rect 293218 297208 293224 297220
rect 216088 297180 293224 297208
rect 216088 297168 216094 297180
rect 293218 297168 293224 297180
rect 293276 297168 293282 297220
rect 98730 297100 98736 297152
rect 98788 297140 98794 297152
rect 236362 297140 236368 297152
rect 98788 297112 236368 297140
rect 98788 297100 98794 297112
rect 236362 297100 236368 297112
rect 236420 297100 236426 297152
rect 112254 297032 112260 297084
rect 112312 297072 112318 297084
rect 235902 297072 235908 297084
rect 112312 297044 235908 297072
rect 112312 297032 112318 297044
rect 235902 297032 235908 297044
rect 235960 297032 235966 297084
rect 126974 296624 126980 296676
rect 127032 296664 127038 296676
rect 243538 296664 243544 296676
rect 127032 296636 243544 296664
rect 127032 296624 127038 296636
rect 243538 296624 243544 296636
rect 243596 296624 243602 296676
rect 153194 296556 153200 296608
rect 153252 296596 153258 296608
rect 248598 296596 248604 296608
rect 153252 296568 248604 296596
rect 153252 296556 153258 296568
rect 248598 296556 248604 296568
rect 248656 296556 248662 296608
rect 209774 296216 209780 296268
rect 209832 296256 209838 296268
rect 286226 296256 286232 296268
rect 209832 296228 286232 296256
rect 209832 296216 209838 296228
rect 286226 296216 286232 296228
rect 286284 296216 286290 296268
rect 129734 296148 129740 296200
rect 129792 296188 129798 296200
rect 273806 296188 273812 296200
rect 129792 296160 273812 296188
rect 129792 296148 129798 296160
rect 273806 296148 273812 296160
rect 273864 296148 273870 296200
rect 318058 296148 318064 296200
rect 318116 296188 318122 296200
rect 400214 296188 400220 296200
rect 318116 296160 400220 296188
rect 318116 296148 318122 296160
rect 400214 296148 400220 296160
rect 400272 296148 400278 296200
rect 125594 296080 125600 296132
rect 125652 296120 125658 296132
rect 272426 296120 272432 296132
rect 125652 296092 272432 296120
rect 125652 296080 125658 296092
rect 272426 296080 272432 296092
rect 272484 296080 272490 296132
rect 322014 296080 322020 296132
rect 322072 296120 322078 296132
rect 421558 296120 421564 296132
rect 322072 296092 421564 296120
rect 322072 296080 322078 296092
rect 421558 296080 421564 296092
rect 421616 296080 421622 296132
rect 63494 296012 63500 296064
rect 63552 296052 63558 296064
rect 262766 296052 262772 296064
rect 63552 296024 262772 296052
rect 63552 296012 63558 296024
rect 262766 296012 262772 296024
rect 262824 296012 262830 296064
rect 335814 296012 335820 296064
rect 335872 296052 335878 296064
rect 516778 296052 516784 296064
rect 335872 296024 516784 296052
rect 335872 296012 335878 296024
rect 516778 296012 516784 296024
rect 516836 296012 516842 296064
rect 16574 295944 16580 295996
rect 16632 295984 16638 295996
rect 255866 295984 255872 295996
rect 16632 295956 255872 295984
rect 16632 295944 16638 295956
rect 255866 295944 255872 295956
rect 255924 295944 255930 295996
rect 344186 295944 344192 295996
rect 344244 295984 344250 295996
rect 563698 295984 563704 295996
rect 344244 295956 563704 295984
rect 344244 295944 344250 295956
rect 563698 295944 563704 295956
rect 563756 295944 563762 295996
rect 217870 295264 217876 295316
rect 217928 295304 217934 295316
rect 296990 295304 296996 295316
rect 217928 295276 296996 295304
rect 217928 295264 217934 295276
rect 296990 295264 296996 295276
rect 297048 295264 297054 295316
rect 215754 295196 215760 295248
rect 215812 295236 215818 295248
rect 297082 295236 297088 295248
rect 215812 295208 297088 295236
rect 215812 295196 215818 295208
rect 297082 295196 297088 295208
rect 297140 295196 297146 295248
rect 215110 295128 215116 295180
rect 215168 295168 215174 295180
rect 296898 295168 296904 295180
rect 215168 295140 296904 295168
rect 215168 295128 215174 295140
rect 296898 295128 296904 295140
rect 296956 295128 296962 295180
rect 214374 295060 214380 295112
rect 214432 295100 214438 295112
rect 296714 295100 296720 295112
rect 214432 295072 296720 295100
rect 214432 295060 214438 295072
rect 296714 295060 296720 295072
rect 296772 295060 296778 295112
rect 212258 294992 212264 295044
rect 212316 295032 212322 295044
rect 295702 295032 295708 295044
rect 212316 295004 295708 295032
rect 212316 294992 212322 295004
rect 295702 294992 295708 295004
rect 295760 294992 295766 295044
rect 211062 294924 211068 294976
rect 211120 294964 211126 294976
rect 295518 294964 295524 294976
rect 211120 294936 295524 294964
rect 211120 294924 211126 294936
rect 295518 294924 295524 294936
rect 295576 294924 295582 294976
rect 210694 294856 210700 294908
rect 210752 294896 210758 294908
rect 295794 294896 295800 294908
rect 210752 294868 295800 294896
rect 210752 294856 210758 294868
rect 295794 294856 295800 294868
rect 295852 294856 295858 294908
rect 210786 294788 210792 294840
rect 210844 294828 210850 294840
rect 295610 294828 295616 294840
rect 210844 294800 295616 294828
rect 210844 294788 210850 294800
rect 295610 294788 295616 294800
rect 295668 294788 295674 294840
rect 168374 294720 168380 294772
rect 168432 294760 168438 294772
rect 278774 294760 278780 294772
rect 168432 294732 278780 294760
rect 168432 294720 168438 294732
rect 278774 294720 278780 294732
rect 278832 294720 278838 294772
rect 313734 294720 313740 294772
rect 313792 294760 313798 294772
rect 380894 294760 380900 294772
rect 313792 294732 380900 294760
rect 313792 294720 313798 294732
rect 380894 294720 380900 294732
rect 380952 294720 380958 294772
rect 135254 294652 135260 294704
rect 135312 294692 135318 294704
rect 274726 294692 274732 294704
rect 135312 294664 274732 294692
rect 135312 294652 135318 294664
rect 274726 294652 274732 294664
rect 274784 294652 274790 294704
rect 329098 294652 329104 294704
rect 329156 294692 329162 294704
rect 468478 294692 468484 294704
rect 329156 294664 468484 294692
rect 329156 294652 329162 294664
rect 468478 294652 468484 294664
rect 468536 294652 468542 294704
rect 43438 294584 43444 294636
rect 43496 294624 43502 294636
rect 258442 294624 258448 294636
rect 43496 294596 258448 294624
rect 43496 294584 43502 294596
rect 258442 294584 258448 294596
rect 258500 294584 258506 294636
rect 337194 294584 337200 294636
rect 337252 294624 337258 294636
rect 525794 294624 525800 294636
rect 337252 294596 525800 294624
rect 337252 294584 337258 294596
rect 525794 294584 525800 294596
rect 525852 294584 525858 294636
rect 215018 294516 215024 294568
rect 215076 294556 215082 294568
rect 294322 294556 294328 294568
rect 215076 294528 294328 294556
rect 215076 294516 215082 294528
rect 294322 294516 294328 294528
rect 294380 294516 294386 294568
rect 218790 294448 218796 294500
rect 218848 294488 218854 294500
rect 295886 294488 295892 294500
rect 218848 294460 295892 294488
rect 218848 294448 218854 294460
rect 295886 294448 295892 294460
rect 295944 294448 295950 294500
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 228358 293944 228364 293956
rect 3384 293916 228364 293944
rect 3384 293904 3390 293916
rect 228358 293904 228364 293916
rect 228416 293904 228422 293956
rect 317782 293496 317788 293548
rect 317840 293536 317846 293548
rect 405734 293536 405740 293548
rect 317840 293508 405740 293536
rect 317840 293496 317846 293508
rect 405734 293496 405740 293508
rect 405792 293496 405798 293548
rect 218698 293428 218704 293480
rect 218756 293468 218762 293480
rect 349706 293468 349712 293480
rect 218756 293440 349712 293468
rect 218756 293428 218762 293440
rect 349706 293428 349712 293440
rect 349764 293428 349770 293480
rect 202874 293360 202880 293412
rect 202932 293400 202938 293412
rect 284662 293400 284668 293412
rect 202932 293372 284668 293400
rect 202932 293360 202938 293372
rect 284662 293360 284668 293372
rect 284720 293360 284726 293412
rect 329006 293360 329012 293412
rect 329064 293400 329070 293412
rect 467098 293400 467104 293412
rect 329064 293372 467104 293400
rect 329064 293360 329070 293372
rect 467098 293360 467104 293372
rect 467156 293360 467162 293412
rect 71038 293292 71044 293344
rect 71096 293332 71102 293344
rect 263594 293332 263600 293344
rect 71096 293304 263600 293332
rect 71096 293292 71102 293304
rect 263594 293292 263600 293304
rect 263652 293292 263658 293344
rect 335722 293292 335728 293344
rect 335780 293332 335786 293344
rect 509878 293332 509884 293344
rect 335780 293304 509884 293332
rect 335780 293292 335786 293304
rect 509878 293292 509884 293304
rect 509936 293292 509942 293344
rect 52454 293224 52460 293276
rect 52512 293264 52518 293276
rect 260834 293264 260840 293276
rect 52512 293236 260840 293264
rect 52512 293224 52518 293236
rect 260834 293224 260840 293236
rect 260892 293224 260898 293276
rect 338574 293224 338580 293276
rect 338632 293264 338638 293276
rect 527818 293264 527824 293276
rect 338632 293236 527824 293264
rect 338632 293224 338638 293236
rect 527818 293224 527824 293236
rect 527876 293224 527882 293276
rect 315022 292000 315028 292052
rect 315080 292040 315086 292052
rect 387058 292040 387064 292052
rect 315080 292012 387064 292040
rect 315080 292000 315086 292012
rect 387058 292000 387064 292012
rect 387116 292000 387122 292052
rect 161474 291932 161480 291984
rect 161532 291972 161538 291984
rect 279142 291972 279148 291984
rect 161532 291944 279148 291972
rect 161532 291932 161538 291944
rect 279142 291932 279148 291944
rect 279200 291932 279206 291984
rect 327534 291932 327540 291984
rect 327592 291972 327598 291984
rect 464338 291972 464344 291984
rect 327592 291944 464344 291972
rect 327592 291932 327598 291944
rect 464338 291932 464344 291944
rect 464396 291932 464402 291984
rect 128354 291864 128360 291916
rect 128412 291904 128418 291916
rect 271138 291904 271144 291916
rect 128412 291876 271144 291904
rect 128412 291864 128418 291876
rect 271138 291864 271144 291876
rect 271196 291864 271202 291916
rect 330110 291864 330116 291916
rect 330168 291904 330174 291916
rect 478138 291904 478144 291916
rect 330168 291876 478144 291904
rect 330168 291864 330174 291876
rect 478138 291864 478144 291876
rect 478196 291864 478202 291916
rect 22094 291796 22100 291848
rect 22152 291836 22158 291848
rect 255682 291836 255688 291848
rect 22152 291808 255688 291836
rect 22152 291796 22158 291808
rect 255682 291796 255688 291808
rect 255740 291796 255746 291848
rect 338482 291796 338488 291848
rect 338540 291836 338546 291848
rect 534718 291836 534724 291848
rect 338540 291808 534724 291836
rect 338540 291796 338546 291808
rect 534718 291796 534724 291808
rect 534776 291796 534782 291848
rect 151814 290708 151820 290760
rect 151872 290748 151878 290760
rect 276014 290748 276020 290760
rect 151872 290720 276020 290748
rect 151872 290708 151878 290720
rect 276014 290708 276020 290720
rect 276072 290708 276078 290760
rect 317690 290708 317696 290760
rect 317748 290748 317754 290760
rect 408494 290748 408500 290760
rect 317748 290720 408500 290748
rect 317748 290708 317754 290720
rect 408494 290708 408500 290720
rect 408552 290708 408558 290760
rect 217686 290640 217692 290692
rect 217744 290680 217750 290692
rect 348510 290680 348516 290692
rect 217744 290652 348516 290680
rect 217744 290640 217750 290652
rect 348510 290640 348516 290652
rect 348568 290640 348574 290692
rect 143534 290572 143540 290624
rect 143592 290612 143598 290624
rect 274634 290612 274640 290624
rect 143592 290584 274640 290612
rect 143592 290572 143598 290584
rect 274634 290572 274640 290584
rect 274692 290572 274698 290624
rect 320634 290572 320640 290624
rect 320692 290612 320698 290624
rect 418154 290612 418160 290624
rect 320692 290584 418160 290612
rect 320692 290572 320698 290584
rect 418154 290572 418160 290584
rect 418212 290572 418218 290624
rect 44174 290504 44180 290556
rect 44232 290544 44238 290556
rect 259822 290544 259828 290556
rect 44232 290516 259828 290544
rect 44232 290504 44238 290516
rect 259822 290504 259828 290516
rect 259880 290504 259886 290556
rect 341242 290504 341248 290556
rect 341300 290544 341306 290556
rect 542998 290544 543004 290556
rect 341300 290516 543004 290544
rect 341300 290504 341306 290516
rect 542998 290504 543004 290516
rect 543056 290504 543062 290556
rect 13078 290436 13084 290488
rect 13136 290476 13142 290488
rect 254302 290476 254308 290488
rect 13136 290448 254308 290476
rect 13136 290436 13142 290448
rect 254302 290436 254308 290448
rect 254360 290436 254366 290488
rect 341334 290436 341340 290488
rect 341392 290476 341398 290488
rect 549898 290476 549904 290488
rect 341392 290448 549904 290476
rect 341392 290436 341398 290448
rect 549898 290436 549904 290448
rect 549956 290436 549962 290488
rect 201494 289280 201500 289332
rect 201552 289320 201558 289332
rect 284570 289320 284576 289332
rect 201552 289292 284576 289320
rect 201552 289280 201558 289292
rect 284570 289280 284576 289292
rect 284628 289280 284634 289332
rect 132494 289212 132500 289264
rect 132552 289252 132558 289264
rect 273622 289252 273628 289264
rect 132552 289224 273628 289252
rect 132552 289212 132558 289224
rect 273622 289212 273628 289224
rect 273680 289212 273686 289264
rect 321922 289212 321928 289264
rect 321980 289252 321986 289264
rect 430574 289252 430580 289264
rect 321980 289224 430580 289252
rect 321980 289212 321986 289224
rect 430574 289212 430580 289224
rect 430632 289212 430638 289264
rect 103514 289144 103520 289196
rect 103572 289184 103578 289196
rect 269758 289184 269764 289196
rect 103572 289156 269764 289184
rect 103572 289144 103578 289156
rect 269758 289144 269764 289156
rect 269816 289144 269822 289196
rect 331490 289144 331496 289196
rect 331548 289184 331554 289196
rect 490006 289184 490012 289196
rect 331548 289156 490012 289184
rect 331548 289144 331554 289156
rect 490006 289144 490012 289156
rect 490064 289144 490070 289196
rect 9674 289076 9680 289128
rect 9732 289116 9738 289128
rect 254210 289116 254216 289128
rect 9732 289088 254216 289116
rect 9732 289076 9738 289088
rect 254210 289076 254216 289088
rect 254268 289076 254274 289128
rect 341150 289076 341156 289128
rect 341208 289116 341214 289128
rect 552658 289116 552664 289128
rect 341208 289088 552664 289116
rect 341208 289076 341214 289088
rect 552658 289076 552664 289088
rect 552716 289076 552722 289128
rect 181438 287784 181444 287836
rect 181496 287824 181502 287836
rect 281902 287824 281908 287836
rect 181496 287796 281908 287824
rect 181496 287784 181502 287796
rect 281902 287784 281908 287796
rect 281960 287784 281966 287836
rect 327442 287784 327448 287836
rect 327500 287824 327506 287836
rect 460198 287824 460204 287836
rect 327500 287796 460204 287824
rect 327500 287784 327506 287796
rect 460198 287784 460204 287796
rect 460256 287784 460262 287836
rect 139394 287716 139400 287768
rect 139452 287756 139458 287768
rect 275094 287756 275100 287768
rect 139452 287728 275100 287756
rect 139452 287716 139458 287728
rect 275094 287716 275100 287728
rect 275152 287716 275158 287768
rect 342622 287716 342628 287768
rect 342680 287756 342686 287768
rect 554038 287756 554044 287768
rect 342680 287728 554044 287756
rect 342680 287716 342686 287728
rect 554038 287716 554044 287728
rect 554096 287716 554102 287768
rect 27614 287648 27620 287700
rect 27672 287688 27678 287700
rect 257154 287688 257160 287700
rect 27672 287660 257160 287688
rect 27672 287648 27678 287660
rect 257154 287648 257160 287660
rect 257212 287648 257218 287700
rect 342714 287648 342720 287700
rect 342772 287688 342778 287700
rect 561674 287688 561680 287700
rect 342772 287660 561680 287688
rect 342772 287648 342778 287660
rect 561674 287648 561680 287660
rect 561732 287648 561738 287700
rect 312170 286560 312176 286612
rect 312228 286600 312234 286612
rect 371234 286600 371240 286612
rect 312228 286572 371240 286600
rect 312228 286560 312234 286572
rect 371234 286560 371240 286572
rect 371292 286560 371298 286612
rect 199470 286492 199476 286544
rect 199528 286532 199534 286544
rect 283282 286532 283288 286544
rect 199528 286504 283288 286532
rect 199528 286492 199534 286504
rect 283282 286492 283288 286504
rect 283340 286492 283346 286544
rect 323394 286492 323400 286544
rect 323452 286532 323458 286544
rect 435358 286532 435364 286544
rect 323452 286504 435364 286532
rect 323452 286492 323458 286504
rect 435358 286492 435364 286504
rect 435416 286492 435422 286544
rect 146294 286424 146300 286476
rect 146352 286464 146358 286476
rect 276474 286464 276480 286476
rect 146352 286436 276480 286464
rect 146352 286424 146358 286436
rect 276474 286424 276480 286436
rect 276532 286424 276538 286476
rect 324866 286424 324872 286476
rect 324924 286464 324930 286476
rect 448514 286464 448520 286476
rect 324924 286436 448520 286464
rect 324924 286424 324930 286436
rect 448514 286424 448520 286436
rect 448572 286424 448578 286476
rect 46934 286356 46940 286408
rect 46992 286396 46998 286408
rect 259730 286396 259736 286408
rect 46992 286368 259736 286396
rect 46992 286356 46998 286368
rect 259730 286356 259736 286368
rect 259788 286356 259794 286408
rect 328914 286356 328920 286408
rect 328972 286396 328978 286408
rect 471974 286396 471980 286408
rect 328972 286368 471980 286396
rect 328972 286356 328978 286368
rect 471974 286356 471980 286368
rect 472032 286356 472038 286408
rect 8294 286288 8300 286340
rect 8352 286328 8358 286340
rect 254118 286328 254124 286340
rect 8352 286300 254124 286328
rect 8352 286288 8358 286300
rect 254118 286288 254124 286300
rect 254176 286288 254182 286340
rect 344094 286288 344100 286340
rect 344152 286328 344158 286340
rect 566458 286328 566464 286340
rect 344152 286300 566464 286328
rect 344152 286288 344158 286300
rect 566458 286288 566464 286300
rect 566516 286288 566522 286340
rect 150434 285132 150440 285184
rect 150492 285172 150498 285184
rect 276382 285172 276388 285184
rect 150492 285144 276388 285172
rect 150492 285132 150498 285144
rect 276382 285132 276388 285144
rect 276440 285132 276446 285184
rect 313642 285132 313648 285184
rect 313700 285172 313706 285184
rect 378134 285172 378140 285184
rect 313700 285144 378140 285172
rect 313700 285132 313706 285144
rect 378134 285132 378140 285144
rect 378192 285132 378198 285184
rect 81434 285064 81440 285116
rect 81492 285104 81498 285116
rect 265526 285104 265532 285116
rect 81492 285076 265532 285104
rect 81492 285064 81498 285076
rect 265526 285064 265532 285076
rect 265584 285064 265590 285116
rect 313550 285064 313556 285116
rect 313608 285104 313614 285116
rect 382274 285104 382280 285116
rect 313608 285076 382280 285104
rect 313608 285064 313614 285076
rect 382274 285064 382280 285076
rect 382332 285064 382338 285116
rect 40034 284996 40040 285048
rect 40092 285036 40098 285048
rect 258350 285036 258356 285048
rect 40092 285008 258356 285036
rect 40092 284996 40098 285008
rect 258350 284996 258356 285008
rect 258408 284996 258414 285048
rect 323302 284996 323308 285048
rect 323360 285036 323366 285048
rect 436094 285036 436100 285048
rect 323360 285008 436100 285036
rect 323360 284996 323366 285008
rect 436094 284996 436100 285008
rect 436152 284996 436158 285048
rect 2774 284928 2780 284980
rect 2832 284968 2838 284980
rect 252830 284968 252836 284980
rect 2832 284940 252836 284968
rect 2832 284928 2838 284940
rect 252830 284928 252836 284940
rect 252888 284928 252894 284980
rect 345474 284928 345480 284980
rect 345532 284968 345538 284980
rect 575474 284968 575480 284980
rect 345532 284940 575480 284968
rect 345532 284928 345538 284940
rect 575474 284928 575480 284940
rect 575532 284928 575538 284980
rect 153194 283840 153200 283892
rect 153252 283880 153258 283892
rect 277854 283880 277860 283892
rect 153252 283852 277860 283880
rect 153252 283840 153258 283852
rect 277854 283840 277860 283852
rect 277912 283840 277918 283892
rect 314930 283840 314936 283892
rect 314988 283880 314994 283892
rect 390554 283880 390560 283892
rect 314988 283852 390560 283880
rect 314988 283840 314994 283852
rect 390554 283840 390560 283852
rect 390612 283840 390618 283892
rect 217594 283772 217600 283824
rect 217652 283812 217658 283824
rect 350626 283812 350632 283824
rect 217652 283784 350632 283812
rect 217652 283772 217658 283784
rect 350626 283772 350632 283784
rect 350684 283772 350690 283824
rect 138014 283704 138020 283756
rect 138072 283744 138078 283756
rect 275002 283744 275008 283756
rect 138072 283716 275008 283744
rect 138072 283704 138078 283716
rect 275002 283704 275008 283716
rect 275060 283704 275066 283756
rect 324774 283704 324780 283756
rect 324832 283744 324838 283756
rect 442258 283744 442264 283756
rect 324832 283716 442264 283744
rect 324832 283704 324838 283716
rect 442258 283704 442264 283716
rect 442316 283704 442322 283756
rect 58618 283636 58624 283688
rect 58676 283676 58682 283688
rect 261294 283676 261300 283688
rect 58676 283648 261300 283676
rect 58676 283636 58682 283648
rect 261294 283636 261300 283648
rect 261352 283636 261358 283688
rect 337102 283636 337108 283688
rect 337160 283676 337166 283688
rect 521654 283676 521660 283688
rect 337160 283648 521660 283676
rect 337160 283636 337166 283648
rect 521654 283636 521660 283648
rect 521712 283636 521718 283688
rect 20714 283568 20720 283620
rect 20772 283608 20778 283620
rect 255590 283608 255596 283620
rect 20772 283580 255596 283608
rect 20772 283568 20778 283580
rect 255590 283568 255596 283580
rect 255648 283568 255654 283620
rect 339770 283568 339776 283620
rect 339828 283608 339834 283620
rect 536098 283608 536104 283620
rect 339828 283580 536104 283608
rect 339828 283568 339834 283580
rect 536098 283568 536104 283580
rect 536156 283568 536162 283620
rect 313458 282412 313464 282464
rect 313516 282452 313522 282464
rect 371878 282452 371884 282464
rect 313516 282424 371884 282452
rect 313516 282412 313522 282424
rect 371878 282412 371884 282424
rect 371936 282412 371942 282464
rect 157334 282344 157340 282396
rect 157392 282384 157398 282396
rect 277762 282384 277768 282396
rect 157392 282356 277768 282384
rect 157392 282344 157398 282356
rect 277762 282344 277768 282356
rect 277820 282344 277826 282396
rect 319162 282344 319168 282396
rect 319220 282384 319226 282396
rect 414658 282384 414664 282396
rect 319220 282356 414664 282384
rect 319220 282344 319226 282356
rect 414658 282344 414664 282356
rect 414716 282344 414722 282396
rect 131114 282276 131120 282328
rect 131172 282316 131178 282328
rect 273530 282316 273536 282328
rect 131172 282288 273536 282316
rect 131172 282276 131178 282288
rect 273530 282276 273536 282288
rect 273588 282276 273594 282328
rect 327350 282276 327356 282328
rect 327408 282316 327414 282328
rect 458818 282316 458824 282328
rect 327408 282288 458824 282316
rect 327408 282276 327414 282288
rect 458818 282276 458824 282288
rect 458876 282276 458882 282328
rect 107654 282208 107660 282260
rect 107712 282248 107718 282260
rect 269574 282248 269580 282260
rect 107712 282220 269580 282248
rect 107712 282208 107718 282220
rect 269574 282208 269580 282220
rect 269632 282208 269638 282260
rect 328822 282208 328828 282260
rect 328880 282248 328886 282260
rect 471238 282248 471244 282260
rect 328880 282220 471244 282248
rect 328880 282208 328886 282220
rect 471238 282208 471244 282220
rect 471296 282208 471302 282260
rect 39298 282140 39304 282192
rect 39356 282180 39362 282192
rect 258258 282180 258264 282192
rect 39356 282152 258264 282180
rect 39356 282140 39362 282152
rect 258258 282140 258264 282152
rect 258316 282140 258322 282192
rect 342530 282140 342536 282192
rect 342588 282180 342594 282192
rect 556246 282180 556252 282192
rect 342588 282152 556252 282180
rect 342588 282140 342594 282152
rect 556246 282140 556252 282152
rect 556304 282140 556310 282192
rect 320542 280984 320548 281036
rect 320600 281024 320606 281036
rect 417418 281024 417424 281036
rect 320600 280996 417424 281024
rect 320600 280984 320606 280996
rect 417418 280984 417424 280996
rect 417476 280984 417482 281036
rect 142154 280916 142160 280968
rect 142212 280956 142218 280968
rect 274910 280956 274916 280968
rect 142212 280928 274916 280956
rect 142212 280916 142218 280928
rect 274910 280916 274916 280928
rect 274968 280916 274974 280968
rect 326062 280916 326068 280968
rect 326120 280956 326126 280968
rect 445018 280956 445024 280968
rect 326120 280928 445024 280956
rect 326120 280916 326126 280928
rect 445018 280916 445024 280928
rect 445076 280916 445082 280968
rect 126974 280848 126980 280900
rect 127032 280888 127038 280900
rect 272242 280888 272248 280900
rect 127032 280860 272248 280888
rect 127032 280848 127038 280860
rect 272242 280848 272248 280860
rect 272300 280848 272306 280900
rect 330018 280848 330024 280900
rect 330076 280888 330082 280900
rect 481726 280888 481732 280900
rect 330076 280860 481732 280888
rect 330076 280848 330082 280860
rect 481726 280848 481732 280860
rect 481784 280848 481790 280900
rect 26234 280780 26240 280832
rect 26292 280820 26298 280832
rect 257062 280820 257068 280832
rect 26292 280792 257068 280820
rect 26292 280780 26298 280792
rect 257062 280780 257068 280792
rect 257120 280780 257126 280832
rect 345382 280780 345388 280832
rect 345440 280820 345446 280832
rect 571978 280820 571984 280832
rect 345440 280792 571984 280820
rect 345440 280780 345446 280792
rect 571978 280780 571984 280792
rect 572036 280780 572042 280832
rect 319070 279624 319076 279676
rect 319128 279664 319134 279676
rect 409874 279664 409880 279676
rect 319128 279636 409880 279664
rect 319128 279624 319134 279636
rect 409874 279624 409880 279636
rect 409932 279624 409938 279676
rect 165614 279556 165620 279608
rect 165672 279596 165678 279608
rect 279050 279596 279056 279608
rect 165672 279568 279056 279596
rect 165672 279556 165678 279568
rect 279050 279556 279056 279568
rect 279108 279556 279114 279608
rect 320450 279556 320456 279608
rect 320508 279596 320514 279608
rect 423674 279596 423680 279608
rect 320508 279568 423680 279596
rect 320508 279556 320514 279568
rect 423674 279556 423680 279568
rect 423732 279556 423738 279608
rect 57238 279488 57244 279540
rect 57296 279528 57302 279540
rect 261202 279528 261208 279540
rect 57296 279500 261208 279528
rect 57296 279488 57302 279500
rect 261202 279488 261208 279500
rect 261260 279488 261266 279540
rect 332962 279488 332968 279540
rect 333020 279528 333026 279540
rect 493318 279528 493324 279540
rect 333020 279500 493324 279528
rect 333020 279488 333026 279500
rect 493318 279488 493324 279500
rect 493376 279488 493382 279540
rect 21358 279420 21364 279472
rect 21416 279460 21422 279472
rect 255498 279460 255504 279472
rect 21416 279432 255504 279460
rect 21416 279420 21422 279432
rect 255498 279420 255504 279432
rect 255556 279420 255562 279472
rect 338390 279420 338396 279472
rect 338448 279460 338454 279472
rect 531314 279460 531320 279472
rect 338448 279432 531320 279460
rect 338448 279420 338454 279432
rect 531314 279420 531320 279432
rect 531372 279420 531378 279472
rect 188338 278264 188344 278316
rect 188396 278304 188402 278316
rect 281810 278304 281816 278316
rect 188396 278276 281816 278304
rect 188396 278264 188402 278276
rect 281810 278264 281816 278276
rect 281868 278264 281874 278316
rect 147674 278196 147680 278248
rect 147732 278236 147738 278248
rect 276290 278236 276296 278248
rect 147732 278208 276296 278236
rect 147732 278196 147738 278208
rect 276290 278196 276296 278208
rect 276348 278196 276354 278248
rect 321830 278196 321836 278248
rect 321888 278236 321894 278248
rect 428458 278236 428464 278248
rect 321888 278208 428464 278236
rect 321888 278196 321894 278208
rect 428458 278196 428464 278208
rect 428516 278196 428522 278248
rect 97994 278128 98000 278180
rect 98052 278168 98058 278180
rect 268194 278168 268200 278180
rect 98052 278140 268200 278168
rect 98052 278128 98058 278140
rect 268194 278128 268200 278140
rect 268252 278128 268258 278180
rect 323210 278128 323216 278180
rect 323268 278168 323274 278180
rect 441614 278168 441620 278180
rect 323268 278140 441620 278168
rect 323268 278128 323274 278140
rect 441614 278128 441620 278140
rect 441672 278128 441678 278180
rect 71774 278060 71780 278112
rect 71832 278100 71838 278112
rect 264146 278100 264152 278112
rect 71832 278072 264152 278100
rect 71832 278060 71838 278072
rect 264146 278060 264152 278072
rect 264204 278060 264210 278112
rect 335630 278060 335636 278112
rect 335688 278100 335694 278112
rect 511258 278100 511264 278112
rect 335688 278072 511264 278100
rect 335688 278060 335694 278072
rect 511258 278060 511264 278072
rect 511316 278060 511322 278112
rect 42794 277992 42800 278044
rect 42852 278032 42858 278044
rect 253382 278032 253388 278044
rect 42852 278004 253388 278032
rect 42852 277992 42858 278004
rect 253382 277992 253388 278004
rect 253440 277992 253446 278044
rect 345290 277992 345296 278044
rect 345348 278032 345354 278044
rect 578234 278032 578240 278044
rect 345348 278004 578240 278032
rect 345348 277992 345354 278004
rect 578234 277992 578240 278004
rect 578292 277992 578298 278044
rect 196618 276904 196624 276956
rect 196676 276944 196682 276956
rect 281718 276944 281724 276956
rect 196676 276916 281724 276944
rect 196676 276904 196682 276916
rect 281718 276904 281724 276916
rect 281776 276904 281782 276956
rect 136634 276836 136640 276888
rect 136692 276876 136698 276888
rect 274818 276876 274824 276888
rect 136692 276848 274824 276876
rect 136692 276836 136698 276848
rect 274818 276836 274824 276848
rect 274876 276836 274882 276888
rect 317598 276836 317604 276888
rect 317656 276876 317662 276888
rect 407206 276876 407212 276888
rect 317656 276848 407212 276876
rect 317656 276836 317662 276848
rect 407206 276836 407212 276848
rect 407264 276836 407270 276888
rect 102134 276768 102140 276820
rect 102192 276808 102198 276820
rect 269482 276808 269488 276820
rect 102192 276780 269488 276808
rect 102192 276768 102198 276780
rect 269482 276768 269488 276780
rect 269540 276768 269546 276820
rect 323118 276768 323124 276820
rect 323176 276808 323182 276820
rect 439498 276808 439504 276820
rect 323176 276780 439504 276808
rect 323176 276768 323182 276780
rect 439498 276768 439504 276780
rect 439556 276768 439562 276820
rect 78674 276700 78680 276752
rect 78732 276740 78738 276752
rect 265434 276740 265440 276752
rect 78732 276712 265440 276740
rect 78732 276700 78738 276712
rect 265434 276700 265440 276712
rect 265492 276700 265498 276752
rect 337010 276700 337016 276752
rect 337068 276740 337074 276752
rect 522298 276740 522304 276752
rect 337068 276712 522304 276740
rect 337068 276700 337074 276712
rect 522298 276700 522304 276712
rect 522356 276700 522362 276752
rect 35894 276632 35900 276684
rect 35952 276672 35958 276684
rect 258166 276672 258172 276684
rect 35952 276644 258172 276672
rect 35952 276632 35958 276644
rect 258166 276632 258172 276644
rect 258224 276632 258230 276684
rect 342438 276632 342444 276684
rect 342496 276672 342502 276684
rect 560294 276672 560300 276684
rect 342496 276644 560300 276672
rect 342496 276632 342502 276644
rect 560294 276632 560300 276644
rect 560352 276632 560358 276684
rect 193306 275544 193312 275596
rect 193364 275584 193370 275596
rect 283190 275584 283196 275596
rect 193364 275556 283196 275584
rect 193364 275544 193370 275556
rect 283190 275544 283196 275556
rect 283248 275544 283254 275596
rect 127066 275476 127072 275528
rect 127124 275516 127130 275528
rect 273438 275516 273444 275528
rect 127124 275488 273444 275516
rect 127124 275476 127130 275488
rect 273438 275476 273444 275488
rect 273496 275476 273502 275528
rect 317506 275476 317512 275528
rect 317564 275516 317570 275528
rect 404998 275516 405004 275528
rect 317564 275488 405004 275516
rect 317564 275476 317570 275488
rect 404998 275476 405004 275488
rect 405056 275476 405062 275528
rect 111794 275408 111800 275460
rect 111852 275448 111858 275460
rect 270954 275448 270960 275460
rect 111852 275420 270960 275448
rect 111852 275408 111858 275420
rect 270954 275408 270960 275420
rect 271012 275408 271018 275460
rect 324682 275408 324688 275460
rect 324740 275448 324746 275460
rect 448606 275448 448612 275460
rect 324740 275420 448612 275448
rect 324740 275408 324746 275420
rect 448606 275408 448612 275420
rect 448664 275408 448670 275460
rect 93854 275340 93860 275392
rect 93912 275380 93918 275392
rect 268102 275380 268108 275392
rect 93912 275352 268108 275380
rect 93912 275340 93918 275352
rect 268102 275340 268108 275352
rect 268160 275340 268166 275392
rect 325970 275340 325976 275392
rect 326028 275380 326034 275392
rect 454678 275380 454684 275392
rect 326028 275352 454684 275380
rect 326028 275340 326034 275352
rect 454678 275340 454684 275352
rect 454736 275340 454742 275392
rect 11054 275272 11060 275324
rect 11112 275312 11118 275324
rect 247678 275312 247684 275324
rect 11112 275284 247684 275312
rect 11112 275272 11118 275284
rect 247678 275272 247684 275284
rect 247736 275272 247742 275324
rect 336918 275272 336924 275324
rect 336976 275312 336982 275324
rect 525058 275312 525064 275324
rect 336976 275284 525064 275312
rect 336976 275272 336982 275284
rect 525058 275272 525064 275284
rect 525116 275272 525122 275324
rect 324590 274184 324596 274236
rect 324648 274224 324654 274236
rect 446398 274224 446404 274236
rect 324648 274196 446404 274224
rect 324648 274184 324654 274196
rect 446398 274184 446404 274196
rect 446456 274184 446462 274236
rect 197354 274116 197360 274168
rect 197412 274156 197418 274168
rect 284478 274156 284484 274168
rect 197412 274128 284484 274156
rect 197412 274116 197418 274128
rect 284478 274116 284484 274128
rect 284536 274116 284542 274168
rect 324498 274116 324504 274168
rect 324556 274156 324562 274168
rect 449894 274156 449900 274168
rect 324556 274128 449900 274156
rect 324556 274116 324562 274128
rect 449894 274116 449900 274128
rect 449952 274116 449958 274168
rect 162854 274048 162860 274100
rect 162912 274088 162918 274100
rect 278958 274088 278964 274100
rect 162912 274060 278964 274088
rect 162912 274048 162918 274060
rect 278958 274048 278964 274060
rect 279016 274048 279022 274100
rect 325878 274048 325884 274100
rect 325936 274088 325942 274100
rect 459554 274088 459560 274100
rect 325936 274060 459560 274088
rect 325936 274048 325942 274060
rect 459554 274048 459560 274060
rect 459612 274048 459618 274100
rect 120074 273980 120080 274032
rect 120132 274020 120138 274032
rect 272150 274020 272156 274032
rect 120132 273992 272156 274020
rect 120132 273980 120138 273992
rect 272150 273980 272156 273992
rect 272208 273980 272214 274032
rect 338298 273980 338304 274032
rect 338356 274020 338362 274032
rect 531406 274020 531412 274032
rect 338356 273992 531412 274020
rect 338356 273980 338362 273992
rect 531406 273980 531412 273992
rect 531464 273980 531470 274032
rect 93946 273912 93952 273964
rect 94004 273952 94010 273964
rect 268010 273952 268016 273964
rect 94004 273924 268016 273952
rect 94004 273912 94010 273924
rect 268010 273912 268016 273924
rect 268068 273912 268074 273964
rect 362218 273912 362224 273964
rect 362276 273952 362282 273964
rect 580166 273952 580172 273964
rect 362276 273924 580172 273952
rect 362276 273912 362282 273924
rect 580166 273912 580172 273924
rect 580224 273912 580230 273964
rect 201586 272756 201592 272808
rect 201644 272796 201650 272808
rect 284386 272796 284392 272808
rect 201644 272768 284392 272796
rect 201644 272756 201650 272768
rect 284386 272756 284392 272768
rect 284444 272756 284450 272808
rect 187694 272688 187700 272740
rect 187752 272728 187758 272740
rect 283098 272728 283104 272740
rect 187752 272700 283104 272728
rect 187752 272688 187758 272700
rect 283098 272688 283104 272700
rect 283156 272688 283162 272740
rect 102226 272620 102232 272672
rect 102284 272660 102290 272672
rect 269390 272660 269396 272672
rect 102284 272632 269396 272660
rect 102284 272620 102290 272632
rect 269390 272620 269396 272632
rect 269448 272620 269454 272672
rect 80054 272552 80060 272604
rect 80112 272592 80118 272604
rect 265342 272592 265348 272604
rect 80112 272564 265348 272592
rect 80112 272552 80118 272564
rect 265342 272552 265348 272564
rect 265400 272552 265406 272604
rect 328730 272552 328736 272604
rect 328788 272592 328794 272604
rect 475378 272592 475384 272604
rect 328788 272564 475384 272592
rect 328788 272552 328794 272564
rect 475378 272552 475384 272564
rect 475436 272552 475442 272604
rect 57974 272484 57980 272536
rect 58032 272524 58038 272536
rect 261110 272524 261116 272536
rect 58032 272496 261116 272524
rect 58032 272484 58038 272496
rect 261110 272484 261116 272496
rect 261168 272484 261174 272536
rect 339678 272484 339684 272536
rect 339736 272524 339742 272536
rect 540238 272524 540244 272536
rect 339736 272496 540244 272524
rect 339736 272484 339742 272496
rect 540238 272484 540244 272496
rect 540296 272484 540302 272536
rect 211798 271396 211804 271448
rect 211856 271436 211862 271448
rect 285858 271436 285864 271448
rect 211856 271408 285864 271436
rect 211856 271396 211862 271408
rect 285858 271396 285864 271408
rect 285916 271396 285922 271448
rect 180794 271328 180800 271380
rect 180852 271368 180858 271380
rect 282086 271368 282092 271380
rect 180852 271340 282092 271368
rect 180852 271328 180858 271340
rect 282086 271328 282092 271340
rect 282144 271328 282150 271380
rect 99374 271260 99380 271312
rect 99432 271300 99438 271312
rect 260190 271300 260196 271312
rect 99432 271272 260196 271300
rect 99432 271260 99438 271272
rect 260190 271260 260196 271272
rect 260248 271260 260254 271312
rect 314838 271260 314844 271312
rect 314896 271300 314902 271312
rect 386414 271300 386420 271312
rect 314896 271272 386420 271300
rect 314896 271260 314902 271272
rect 386414 271260 386420 271272
rect 386472 271260 386478 271312
rect 77294 271192 77300 271244
rect 77352 271232 77358 271244
rect 265250 271232 265256 271244
rect 77352 271204 265256 271232
rect 77352 271192 77358 271204
rect 265250 271192 265256 271204
rect 265308 271192 265314 271244
rect 329926 271192 329932 271244
rect 329984 271232 329990 271244
rect 484394 271232 484400 271244
rect 329984 271204 484400 271232
rect 329984 271192 329990 271204
rect 484394 271192 484400 271204
rect 484452 271192 484458 271244
rect 53834 271124 53840 271176
rect 53892 271164 53898 271176
rect 261018 271164 261024 271176
rect 53892 271136 261024 271164
rect 53892 271124 53898 271136
rect 261018 271124 261024 271136
rect 261076 271124 261082 271176
rect 339586 271124 339592 271176
rect 339644 271164 339650 271176
rect 545114 271164 545120 271176
rect 339644 271136 545120 271164
rect 339644 271124 339650 271136
rect 545114 271124 545120 271136
rect 545172 271124 545178 271176
rect 166994 269968 167000 270020
rect 167052 270008 167058 270020
rect 278866 270008 278872 270020
rect 167052 269980 278872 270008
rect 167052 269968 167058 269980
rect 278866 269968 278872 269980
rect 278924 269968 278930 270020
rect 314746 269968 314752 270020
rect 314804 270008 314810 270020
rect 390646 270008 390652 270020
rect 314804 269980 390652 270008
rect 314804 269968 314810 269980
rect 390646 269968 390652 269980
rect 390704 269968 390710 270020
rect 92474 269900 92480 269952
rect 92532 269940 92538 269952
rect 266814 269940 266820 269952
rect 92532 269912 266820 269940
rect 92532 269900 92538 269912
rect 266814 269900 266820 269912
rect 266872 269900 266878 269952
rect 331398 269900 331404 269952
rect 331456 269940 331462 269952
rect 486418 269940 486424 269952
rect 331456 269912 486424 269940
rect 331456 269900 331462 269912
rect 486418 269900 486424 269912
rect 486476 269900 486482 269952
rect 75914 269832 75920 269884
rect 75972 269872 75978 269884
rect 264054 269872 264060 269884
rect 75972 269844 264060 269872
rect 75972 269832 75978 269844
rect 264054 269832 264060 269844
rect 264112 269832 264118 269884
rect 335538 269832 335544 269884
rect 335596 269872 335602 269884
rect 517514 269872 517520 269884
rect 335596 269844 517520 269872
rect 335596 269832 335602 269844
rect 517514 269832 517520 269844
rect 517572 269832 517578 269884
rect 14458 269764 14464 269816
rect 14516 269804 14522 269816
rect 254026 269804 254032 269816
rect 14516 269776 254032 269804
rect 14516 269764 14522 269776
rect 254026 269764 254032 269776
rect 254084 269764 254090 269816
rect 341058 269764 341064 269816
rect 341116 269804 341122 269816
rect 552014 269804 552020 269816
rect 341116 269776 552020 269804
rect 341116 269764 341122 269776
rect 552014 269764 552020 269776
rect 552072 269764 552078 269816
rect 144914 268472 144920 268524
rect 144972 268512 144978 268524
rect 276198 268512 276204 268524
rect 144972 268484 276204 268512
rect 144972 268472 144978 268484
rect 276198 268472 276204 268484
rect 276256 268472 276262 268524
rect 74534 268404 74540 268456
rect 74592 268444 74598 268456
rect 263962 268444 263968 268456
rect 74592 268416 263968 268444
rect 74592 268404 74598 268416
rect 263962 268404 263968 268416
rect 264020 268404 264026 268456
rect 327258 268404 327264 268456
rect 327316 268444 327322 268456
rect 467834 268444 467840 268456
rect 327316 268416 467840 268444
rect 327316 268404 327322 268416
rect 467834 268404 467840 268416
rect 467892 268404 467898 268456
rect 7558 268336 7564 268388
rect 7616 268376 7622 268388
rect 252738 268376 252744 268388
rect 7616 268348 252744 268376
rect 7616 268336 7622 268348
rect 252738 268336 252744 268348
rect 252796 268336 252802 268388
rect 328638 268336 328644 268388
rect 328696 268376 328702 268388
rect 473446 268376 473452 268388
rect 328696 268348 473452 268376
rect 328696 268336 328702 268348
rect 473446 268336 473452 268348
rect 473504 268336 473510 268388
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 225598 267696 225604 267708
rect 3016 267668 225604 267696
rect 3016 267656 3022 267668
rect 225598 267656 225604 267668
rect 225656 267656 225662 267708
rect 218606 267180 218612 267232
rect 218664 267220 218670 267232
rect 347866 267220 347872 267232
rect 218664 267192 347872 267220
rect 218664 267180 218670 267192
rect 347866 267180 347872 267192
rect 347924 267180 347930 267232
rect 332870 267112 332876 267164
rect 332928 267152 332934 267164
rect 495434 267152 495440 267164
rect 332928 267124 495440 267152
rect 332928 267112 332934 267124
rect 495434 267112 495440 267124
rect 495492 267112 495498 267164
rect 67634 267044 67640 267096
rect 67692 267084 67698 267096
rect 263870 267084 263876 267096
rect 67692 267056 263876 267084
rect 67692 267044 67698 267056
rect 263870 267044 263876 267056
rect 263928 267044 263934 267096
rect 340966 267044 340972 267096
rect 341024 267084 341030 267096
rect 553394 267084 553400 267096
rect 341024 267056 553400 267084
rect 341024 267044 341030 267056
rect 553394 267044 553400 267056
rect 553452 267044 553458 267096
rect 48314 266976 48320 267028
rect 48372 267016 48378 267028
rect 259638 267016 259644 267028
rect 48372 266988 259644 267016
rect 48372 266976 48378 266988
rect 259638 266976 259644 266988
rect 259696 266976 259702 267028
rect 344002 266976 344008 267028
rect 344060 267016 344066 267028
rect 565814 267016 565820 267028
rect 344060 266988 565820 267016
rect 344060 266976 344066 266988
rect 565814 266976 565820 266988
rect 565872 266976 565878 267028
rect 191834 265888 191840 265940
rect 191892 265928 191898 265940
rect 283466 265928 283472 265940
rect 191892 265900 283472 265928
rect 191892 265888 191898 265900
rect 283466 265888 283472 265900
rect 283524 265888 283530 265940
rect 133874 265820 133880 265872
rect 133932 265860 133938 265872
rect 273346 265860 273352 265872
rect 133932 265832 273352 265860
rect 133932 265820 133938 265832
rect 273346 265820 273352 265832
rect 273404 265820 273410 265872
rect 115934 265752 115940 265804
rect 115992 265792 115998 265804
rect 270770 265792 270776 265804
rect 115992 265764 270776 265792
rect 115992 265752 115998 265764
rect 270770 265752 270776 265764
rect 270828 265752 270834 265804
rect 331306 265752 331312 265804
rect 331364 265792 331370 265804
rect 491294 265792 491300 265804
rect 331364 265764 491300 265792
rect 331364 265752 331370 265764
rect 491294 265752 491300 265764
rect 491352 265752 491358 265804
rect 114554 265684 114560 265736
rect 114612 265724 114618 265736
rect 270862 265724 270868 265736
rect 114612 265696 270868 265724
rect 114612 265684 114618 265696
rect 270862 265684 270868 265696
rect 270920 265684 270926 265736
rect 338206 265684 338212 265736
rect 338264 265724 338270 265736
rect 535454 265724 535460 265736
rect 338264 265696 535460 265724
rect 338264 265684 338270 265696
rect 535454 265684 535460 265696
rect 535512 265684 535518 265736
rect 31754 265616 31760 265668
rect 31812 265656 31818 265668
rect 250530 265656 250536 265668
rect 31812 265628 250536 265656
rect 31812 265616 31818 265628
rect 250530 265616 250536 265628
rect 250588 265616 250594 265668
rect 342346 265616 342352 265668
rect 342404 265656 342410 265668
rect 560938 265656 560944 265668
rect 342404 265628 560944 265656
rect 342404 265616 342410 265628
rect 560938 265616 560944 265628
rect 560996 265616 561002 265668
rect 143626 264392 143632 264444
rect 143684 264432 143690 264444
rect 275278 264432 275284 264444
rect 143684 264404 275284 264432
rect 143684 264392 143690 264404
rect 275278 264392 275284 264404
rect 275336 264392 275342 264444
rect 113174 264324 113180 264376
rect 113232 264364 113238 264376
rect 270678 264364 270684 264376
rect 113232 264336 270684 264364
rect 113232 264324 113238 264336
rect 270678 264324 270684 264336
rect 270736 264324 270742 264376
rect 313274 264324 313280 264376
rect 313332 264364 313338 264376
rect 382366 264364 382372 264376
rect 313332 264336 382372 264364
rect 313332 264324 313338 264336
rect 382366 264324 382372 264336
rect 382424 264324 382430 264376
rect 96614 264256 96620 264308
rect 96672 264296 96678 264308
rect 267918 264296 267924 264308
rect 96672 264268 267924 264296
rect 96672 264256 96678 264268
rect 267918 264256 267924 264268
rect 267976 264256 267982 264308
rect 320358 264256 320364 264308
rect 320416 264296 320422 264308
rect 420914 264296 420920 264308
rect 320416 264268 420920 264296
rect 320416 264256 320422 264268
rect 420914 264256 420920 264268
rect 420972 264256 420978 264308
rect 84194 264188 84200 264240
rect 84252 264228 84258 264240
rect 265158 264228 265164 264240
rect 84252 264200 265164 264228
rect 84252 264188 84258 264200
rect 265158 264188 265164 264200
rect 265216 264188 265222 264240
rect 340874 264188 340880 264240
rect 340932 264228 340938 264240
rect 549254 264228 549260 264240
rect 340932 264200 549260 264228
rect 340932 264188 340938 264200
rect 549254 264188 549260 264200
rect 549312 264188 549318 264240
rect 314654 262964 314660 263016
rect 314712 263004 314718 263016
rect 389174 263004 389180 263016
rect 314712 262976 389180 263004
rect 314712 262964 314718 262976
rect 389174 262964 389180 262976
rect 389232 262964 389238 263016
rect 154574 262896 154580 262948
rect 154632 262936 154638 262948
rect 277670 262936 277676 262948
rect 154632 262908 277676 262936
rect 154632 262896 154638 262908
rect 277670 262896 277676 262908
rect 277728 262896 277734 262948
rect 323026 262896 323032 262948
rect 323084 262936 323090 262948
rect 434714 262936 434720 262948
rect 323084 262908 434720 262936
rect 323084 262896 323090 262908
rect 434714 262896 434720 262908
rect 434772 262896 434778 262948
rect 151906 262828 151912 262880
rect 151964 262868 151970 262880
rect 276106 262868 276112 262880
rect 151964 262840 276112 262868
rect 151964 262828 151970 262840
rect 276106 262828 276112 262840
rect 276164 262828 276170 262880
rect 345198 262828 345204 262880
rect 345256 262868 345262 262880
rect 574094 262868 574100 262880
rect 345256 262840 574100 262868
rect 345256 262828 345262 262840
rect 574094 262828 574100 262840
rect 574152 262828 574158 262880
rect 212534 261808 212540 261860
rect 212592 261848 212598 261860
rect 287330 261848 287336 261860
rect 212592 261820 287336 261848
rect 212592 261808 212598 261820
rect 287330 261808 287336 261820
rect 287388 261808 287394 261860
rect 158714 261740 158720 261792
rect 158772 261780 158778 261792
rect 277578 261780 277584 261792
rect 158772 261752 277584 261780
rect 158772 261740 158778 261752
rect 277578 261740 277584 261752
rect 277636 261740 277642 261792
rect 316586 261740 316592 261792
rect 316644 261780 316650 261792
rect 393314 261780 393320 261792
rect 316644 261752 393320 261780
rect 316644 261740 316650 261752
rect 393314 261740 393320 261752
rect 393372 261740 393378 261792
rect 149054 261672 149060 261724
rect 149112 261712 149118 261724
rect 276566 261712 276572 261724
rect 149112 261684 276572 261712
rect 149112 261672 149118 261684
rect 276566 261672 276572 261684
rect 276624 261672 276630 261724
rect 316494 261672 316500 261724
rect 316552 261712 316558 261724
rect 397454 261712 397460 261724
rect 316552 261684 397460 261712
rect 316552 261672 316558 261684
rect 397454 261672 397460 261684
rect 397512 261672 397518 261724
rect 217778 261604 217784 261656
rect 217836 261644 217842 261656
rect 345106 261644 345112 261656
rect 217836 261616 345112 261644
rect 217836 261604 217842 261616
rect 345106 261604 345112 261616
rect 345164 261604 345170 261656
rect 69014 261536 69020 261588
rect 69072 261576 69078 261588
rect 263778 261576 263784 261588
rect 69072 261548 263784 261576
rect 69072 261536 69078 261548
rect 263778 261536 263784 261548
rect 263836 261536 263842 261588
rect 329834 261536 329840 261588
rect 329892 261576 329898 261588
rect 485774 261576 485780 261588
rect 329892 261548 485780 261576
rect 329892 261536 329898 261548
rect 485774 261536 485780 261548
rect 485832 261536 485838 261588
rect 13814 261468 13820 261520
rect 13872 261508 13878 261520
rect 254394 261508 254400 261520
rect 13872 261480 254400 261508
rect 13872 261468 13878 261480
rect 254394 261468 254400 261480
rect 254452 261468 254458 261520
rect 343910 261468 343916 261520
rect 343968 261508 343974 261520
rect 569954 261508 569960 261520
rect 343968 261480 569960 261508
rect 343968 261468 343974 261480
rect 569954 261468 569960 261480
rect 570012 261468 570018 261520
rect 124214 260312 124220 260364
rect 124272 260352 124278 260364
rect 251910 260352 251916 260364
rect 124272 260324 251916 260352
rect 124272 260312 124278 260324
rect 251910 260312 251916 260324
rect 251968 260312 251974 260364
rect 39390 260244 39396 260296
rect 39448 260284 39454 260296
rect 256878 260284 256884 260296
rect 39448 260256 256884 260284
rect 39448 260244 39454 260256
rect 256878 260244 256884 260256
rect 256936 260244 256942 260296
rect 30374 260176 30380 260228
rect 30432 260216 30438 260228
rect 256970 260216 256976 260228
rect 30432 260188 256976 260216
rect 30432 260176 30438 260188
rect 256970 260176 256976 260188
rect 257028 260176 257034 260228
rect 339494 260176 339500 260228
rect 339552 260216 339558 260228
rect 542354 260216 542360 260228
rect 339552 260188 542360 260216
rect 339552 260176 339558 260188
rect 542354 260176 542360 260188
rect 542412 260176 542418 260228
rect 4154 260108 4160 260160
rect 4212 260148 4218 260160
rect 246298 260148 246304 260160
rect 4212 260120 246304 260148
rect 4212 260108 4218 260120
rect 246298 260108 246304 260120
rect 246356 260108 246362 260160
rect 342254 260108 342260 260160
rect 342312 260148 342318 260160
rect 558914 260148 558920 260160
rect 342312 260120 558920 260148
rect 342312 260108 342318 260120
rect 558914 260108 558920 260120
rect 558972 260108 558978 260160
rect 374638 259360 374644 259412
rect 374696 259400 374702 259412
rect 580166 259400 580172 259412
rect 374696 259372 580172 259400
rect 374696 259360 374702 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 176654 258816 176660 258868
rect 176712 258856 176718 258868
rect 266998 258856 267004 258868
rect 176712 258828 267004 258856
rect 176712 258816 176718 258828
rect 266998 258816 267004 258828
rect 267056 258816 267062 258868
rect 173894 258748 173900 258800
rect 173952 258788 173958 258800
rect 280614 258788 280620 258800
rect 173952 258760 280620 258788
rect 173952 258748 173958 258760
rect 280614 258748 280620 258760
rect 280672 258748 280678 258800
rect 316402 258748 316408 258800
rect 316460 258788 316466 258800
rect 398834 258788 398840 258800
rect 316460 258760 398840 258788
rect 316460 258748 316466 258760
rect 398834 258748 398840 258760
rect 398892 258748 398898 258800
rect 217502 258680 217508 258732
rect 217560 258720 217566 258732
rect 346486 258720 346492 258732
rect 217560 258692 346492 258720
rect 217560 258680 217566 258692
rect 346486 258680 346492 258692
rect 346544 258680 346550 258732
rect 117314 257524 117320 257576
rect 117372 257564 117378 257576
rect 260098 257564 260104 257576
rect 117372 257536 260104 257564
rect 117372 257524 117378 257536
rect 260098 257524 260104 257536
rect 260156 257524 260162 257576
rect 106274 257456 106280 257508
rect 106332 257496 106338 257508
rect 261478 257496 261484 257508
rect 106332 257468 261484 257496
rect 106332 257456 106338 257468
rect 261478 257456 261484 257468
rect 261536 257456 261542 257508
rect 23474 257388 23480 257440
rect 23532 257428 23538 257440
rect 251818 257428 251824 257440
rect 23532 257400 251824 257428
rect 23532 257388 23538 257400
rect 251818 257388 251824 257400
rect 251876 257388 251882 257440
rect 316310 257388 316316 257440
rect 316368 257428 316374 257440
rect 391934 257428 391940 257440
rect 316368 257400 391940 257428
rect 316368 257388 316374 257400
rect 391934 257388 391940 257400
rect 391992 257388 391998 257440
rect 25590 257320 25596 257372
rect 25648 257360 25654 257372
rect 255406 257360 255412 257372
rect 25648 257332 255412 257360
rect 25648 257320 25654 257332
rect 255406 257320 255412 257332
rect 255464 257320 255470 257372
rect 316218 257320 316224 257372
rect 316276 257360 316282 257372
rect 396074 257360 396080 257372
rect 316276 257332 396080 257360
rect 316276 257320 316282 257332
rect 396074 257320 396080 257332
rect 396132 257320 396138 257372
rect 218422 256300 218428 256352
rect 218480 256340 218486 256352
rect 287238 256340 287244 256352
rect 218480 256312 287244 256340
rect 218480 256300 218486 256312
rect 287238 256300 287244 256312
rect 287296 256300 287302 256352
rect 217226 256232 217232 256284
rect 217284 256272 217290 256284
rect 350534 256272 350540 256284
rect 217284 256244 350540 256272
rect 217284 256232 217290 256244
rect 350534 256232 350540 256244
rect 350592 256232 350598 256284
rect 122834 256164 122840 256216
rect 122892 256204 122898 256216
rect 271966 256204 271972 256216
rect 122892 256176 271972 256204
rect 122892 256164 122898 256176
rect 271966 256164 271972 256176
rect 272024 256164 272030 256216
rect 318978 256164 318984 256216
rect 319036 256204 319042 256216
rect 413278 256204 413284 256216
rect 319036 256176 413284 256204
rect 319036 256164 319042 256176
rect 413278 256164 413284 256176
rect 413336 256164 413342 256216
rect 118694 256096 118700 256148
rect 118752 256136 118758 256148
rect 272058 256136 272064 256148
rect 118752 256108 272064 256136
rect 118752 256096 118758 256108
rect 272058 256096 272064 256108
rect 272116 256096 272122 256148
rect 320266 256096 320272 256148
rect 320324 256136 320330 256148
rect 425054 256136 425060 256148
rect 320324 256108 425060 256136
rect 320324 256096 320330 256108
rect 425054 256096 425060 256108
rect 425112 256096 425118 256148
rect 77386 256028 77392 256080
rect 77444 256068 77450 256080
rect 265066 256068 265072 256080
rect 77444 256040 265072 256068
rect 77444 256028 77450 256040
rect 265066 256028 265072 256040
rect 265124 256028 265130 256080
rect 321738 256028 321744 256080
rect 321796 256068 321802 256080
rect 431954 256068 431960 256080
rect 321796 256040 431960 256068
rect 321796 256028 321802 256040
rect 431954 256028 431960 256040
rect 432012 256028 432018 256080
rect 17954 255960 17960 256012
rect 18012 256000 18018 256012
rect 255774 256000 255780 256012
rect 18012 255972 255780 256000
rect 18012 255960 18018 255972
rect 255774 255960 255780 255972
rect 255832 255960 255838 256012
rect 324406 255960 324412 256012
rect 324464 256000 324470 256012
rect 445110 256000 445116 256012
rect 324464 255972 445116 256000
rect 324464 255960 324470 255972
rect 445110 255960 445116 255972
rect 445168 255960 445174 256012
rect 169754 254804 169760 254856
rect 169812 254844 169818 254856
rect 280522 254844 280528 254856
rect 169812 254816 280528 254844
rect 169812 254804 169818 254816
rect 280522 254804 280528 254816
rect 280580 254804 280586 254856
rect 311986 254804 311992 254856
rect 312044 254844 312050 254856
rect 372614 254844 372620 254856
rect 312044 254816 372620 254844
rect 312044 254804 312050 254816
rect 372614 254804 372620 254816
rect 372672 254804 372678 254856
rect 3326 254736 3332 254788
rect 3384 254776 3390 254788
rect 8938 254776 8944 254788
rect 3384 254748 8944 254776
rect 3384 254736 3390 254748
rect 8938 254736 8944 254748
rect 8996 254736 9002 254788
rect 110414 254736 110420 254788
rect 110472 254776 110478 254788
rect 269298 254776 269304 254788
rect 110472 254748 269304 254776
rect 110472 254736 110478 254748
rect 269298 254736 269304 254748
rect 269356 254736 269362 254788
rect 317414 254736 317420 254788
rect 317472 254776 317478 254788
rect 404354 254776 404360 254788
rect 317472 254748 404360 254776
rect 317472 254736 317478 254748
rect 404354 254736 404360 254748
rect 404412 254736 404418 254788
rect 88334 254668 88340 254720
rect 88392 254708 88398 254720
rect 253290 254708 253296 254720
rect 88392 254680 253296 254708
rect 88392 254668 88398 254680
rect 253290 254668 253296 254680
rect 253348 254668 253354 254720
rect 328546 254668 328552 254720
rect 328604 254708 328610 254720
rect 474734 254708 474740 254720
rect 328604 254680 474740 254708
rect 328604 254668 328610 254680
rect 474734 254668 474740 254680
rect 474792 254668 474798 254720
rect 91094 254600 91100 254652
rect 91152 254640 91158 254652
rect 266722 254640 266728 254652
rect 91152 254612 266728 254640
rect 91152 254600 91158 254612
rect 266722 254600 266728 254612
rect 266780 254600 266786 254652
rect 343726 254600 343732 254652
rect 343784 254640 343790 254652
rect 564526 254640 564532 254652
rect 343784 254612 564532 254640
rect 343784 254600 343790 254612
rect 564526 254600 564532 254612
rect 564584 254600 564590 254652
rect 86954 254532 86960 254584
rect 87012 254572 87018 254584
rect 266630 254572 266636 254584
rect 87012 254544 266636 254572
rect 87012 254532 87018 254544
rect 266630 254532 266636 254544
rect 266688 254532 266694 254584
rect 343818 254532 343824 254584
rect 343876 254572 343882 254584
rect 567194 254572 567200 254584
rect 343876 254544 567200 254572
rect 343876 254532 343882 254544
rect 567194 254532 567200 254544
rect 567252 254532 567258 254584
rect 303982 253852 303988 253904
rect 304040 253892 304046 253904
rect 364334 253892 364340 253904
rect 304040 253864 364340 253892
rect 304040 253852 304046 253864
rect 364334 253852 364340 253864
rect 364392 253852 364398 253904
rect 303890 253784 303896 253836
rect 303948 253824 303954 253836
rect 365806 253824 365812 253836
rect 303948 253796 365812 253824
rect 303948 253784 303954 253796
rect 365806 253784 365812 253796
rect 365864 253784 365870 253836
rect 301038 253716 301044 253768
rect 301096 253756 301102 253768
rect 367186 253756 367192 253768
rect 301096 253728 367192 253756
rect 301096 253716 301102 253728
rect 367186 253716 367192 253728
rect 367244 253716 367250 253768
rect 300946 253648 300952 253700
rect 301004 253688 301010 253700
rect 368474 253688 368480 253700
rect 301004 253660 368480 253688
rect 301004 253648 301010 253660
rect 368474 253648 368480 253660
rect 368532 253648 368538 253700
rect 316034 253580 316040 253632
rect 316092 253620 316098 253632
rect 394694 253620 394700 253632
rect 316092 253592 394700 253620
rect 316092 253580 316098 253592
rect 394694 253580 394700 253592
rect 394752 253580 394758 253632
rect 176746 253512 176752 253564
rect 176804 253552 176810 253564
rect 280430 253552 280436 253564
rect 176804 253524 280436 253552
rect 176804 253512 176810 253524
rect 280430 253512 280436 253524
rect 280488 253512 280494 253564
rect 316126 253512 316132 253564
rect 316184 253552 316190 253564
rect 398926 253552 398932 253564
rect 316184 253524 398932 253552
rect 316184 253512 316190 253524
rect 398926 253512 398932 253524
rect 398984 253512 398990 253564
rect 217134 253444 217140 253496
rect 217192 253484 217198 253496
rect 348418 253484 348424 253496
rect 217192 253456 348424 253484
rect 217192 253444 217198 253456
rect 348418 253444 348424 253456
rect 348476 253444 348482 253496
rect 118786 253376 118792 253428
rect 118844 253416 118850 253428
rect 271046 253416 271052 253428
rect 118844 253388 271052 253416
rect 118844 253376 118850 253388
rect 271046 253376 271052 253388
rect 271104 253376 271110 253428
rect 332686 253376 332692 253428
rect 332744 253416 332750 253428
rect 496078 253416 496084 253428
rect 332744 253388 496084 253416
rect 332744 253376 332750 253388
rect 496078 253376 496084 253388
rect 496136 253376 496142 253428
rect 110506 253308 110512 253360
rect 110564 253348 110570 253360
rect 270586 253348 270592 253360
rect 110564 253320 270592 253348
rect 110564 253308 110570 253320
rect 270586 253308 270592 253320
rect 270644 253308 270650 253360
rect 332778 253308 332784 253360
rect 332836 253348 332842 253360
rect 499574 253348 499580 253360
rect 332836 253320 499580 253348
rect 332836 253308 332842 253320
rect 499574 253308 499580 253320
rect 499632 253308 499638 253360
rect 95234 253240 95240 253292
rect 95292 253280 95298 253292
rect 267826 253280 267832 253292
rect 95292 253252 267832 253280
rect 95292 253240 95298 253252
rect 267826 253240 267832 253252
rect 267884 253240 267890 253292
rect 334618 253240 334624 253292
rect 334676 253280 334682 253292
rect 506474 253280 506480 253292
rect 334676 253252 506480 253280
rect 334676 253240 334682 253252
rect 506474 253240 506480 253252
rect 506532 253240 506538 253292
rect 73154 253172 73160 253224
rect 73212 253212 73218 253224
rect 263686 253212 263692 253224
rect 73212 253184 263692 253212
rect 73212 253172 73218 253184
rect 263686 253172 263692 253184
rect 263744 253172 263750 253224
rect 336826 253172 336832 253224
rect 336884 253212 336890 253224
rect 528554 253212 528560 253224
rect 336884 253184 528560 253212
rect 336884 253172 336890 253184
rect 528554 253172 528560 253184
rect 528612 253172 528618 253224
rect 302510 253104 302516 253156
rect 302568 253144 302574 253156
rect 360194 253144 360200 253156
rect 302568 253116 360200 253144
rect 302568 253104 302574 253116
rect 360194 253104 360200 253116
rect 360252 253104 360258 253156
rect 302602 253036 302608 253088
rect 302660 253076 302666 253088
rect 358814 253076 358820 253088
rect 302660 253048 358820 253076
rect 302660 253036 302666 253048
rect 358814 253036 358820 253048
rect 358872 253036 358878 253088
rect 172514 252220 172520 252272
rect 172572 252260 172578 252272
rect 280338 252260 280344 252272
rect 172572 252232 280344 252260
rect 172572 252220 172578 252232
rect 280338 252220 280344 252232
rect 280396 252220 280402 252272
rect 160186 252152 160192 252204
rect 160244 252192 160250 252204
rect 277394 252192 277400 252204
rect 160244 252164 277400 252192
rect 160244 252152 160250 252164
rect 277394 252152 277400 252164
rect 277452 252152 277458 252204
rect 321646 252152 321652 252204
rect 321704 252192 321710 252204
rect 427814 252192 427820 252204
rect 321704 252164 427820 252192
rect 321704 252152 321710 252164
rect 427814 252152 427820 252164
rect 427872 252152 427878 252204
rect 155954 252084 155960 252136
rect 156012 252124 156018 252136
rect 277486 252124 277492 252136
rect 156012 252096 277492 252124
rect 156012 252084 156018 252096
rect 277486 252084 277492 252096
rect 277544 252084 277550 252136
rect 321554 252084 321560 252136
rect 321612 252124 321618 252136
rect 432046 252124 432052 252136
rect 321612 252096 432052 252124
rect 321612 252084 321618 252096
rect 432046 252084 432052 252096
rect 432104 252084 432110 252136
rect 218514 252016 218520 252068
rect 218572 252056 218578 252068
rect 347774 252056 347780 252068
rect 218572 252028 347780 252056
rect 218572 252016 218578 252028
rect 347774 252016 347780 252028
rect 347832 252016 347838 252068
rect 60734 251948 60740 252000
rect 60792 251988 60798 252000
rect 253198 251988 253204 252000
rect 60792 251960 253204 251988
rect 60792 251948 60798 251960
rect 253198 251948 253204 251960
rect 253256 251948 253262 252000
rect 325786 251948 325792 252000
rect 325844 251988 325850 252000
rect 454034 251988 454040 252000
rect 325844 251960 454040 251988
rect 325844 251948 325850 251960
rect 454034 251948 454040 251960
rect 454092 251948 454098 252000
rect 49694 251880 49700 251932
rect 49752 251920 49758 251932
rect 259546 251920 259552 251932
rect 49752 251892 259552 251920
rect 49752 251880 49758 251892
rect 259546 251880 259552 251892
rect 259604 251880 259610 251932
rect 327166 251880 327172 251932
rect 327224 251920 327230 251932
rect 466454 251920 466460 251932
rect 327224 251892 466460 251920
rect 327224 251880 327230 251892
rect 466454 251880 466460 251892
rect 466512 251880 466518 251932
rect 46198 251812 46204 251864
rect 46256 251852 46262 251864
rect 260006 251852 260012 251864
rect 46256 251824 260012 251852
rect 46256 251812 46262 251824
rect 260006 251812 260012 251824
rect 260064 251812 260070 251864
rect 334526 251812 334532 251864
rect 334584 251852 334590 251864
rect 509234 251852 509240 251864
rect 334584 251824 509240 251852
rect 334584 251812 334590 251824
rect 509234 251812 509240 251824
rect 509292 251812 509298 251864
rect 309594 251132 309600 251184
rect 309652 251172 309658 251184
rect 365714 251172 365720 251184
rect 309652 251144 365720 251172
rect 309652 251132 309658 251144
rect 365714 251132 365720 251144
rect 365772 251132 365778 251184
rect 306742 251064 306748 251116
rect 306800 251104 306806 251116
rect 363138 251104 363144 251116
rect 306800 251076 363144 251104
rect 306800 251064 306806 251076
rect 363138 251064 363144 251076
rect 363196 251064 363202 251116
rect 306834 250996 306840 251048
rect 306892 251036 306898 251048
rect 363230 251036 363236 251048
rect 306892 251008 363236 251036
rect 306892 250996 306898 251008
rect 363230 250996 363236 251008
rect 363288 250996 363294 251048
rect 308214 250928 308220 250980
rect 308272 250968 308278 250980
rect 365990 250968 365996 250980
rect 308272 250940 365996 250968
rect 308272 250928 308278 250940
rect 365990 250928 365996 250940
rect 366048 250928 366054 250980
rect 305454 250860 305460 250912
rect 305512 250900 305518 250912
rect 363322 250900 363328 250912
rect 305512 250872 363328 250900
rect 305512 250860 305518 250872
rect 363322 250860 363328 250872
rect 363380 250860 363386 250912
rect 209866 250792 209872 250844
rect 209924 250832 209930 250844
rect 286042 250832 286048 250844
rect 209924 250804 286048 250832
rect 209924 250792 209930 250804
rect 286042 250792 286048 250804
rect 286100 250792 286106 250844
rect 302418 250792 302424 250844
rect 302476 250832 302482 250844
rect 360286 250832 360292 250844
rect 302476 250804 360292 250832
rect 302476 250792 302482 250804
rect 360286 250792 360292 250804
rect 360344 250792 360350 250844
rect 135346 250724 135352 250776
rect 135404 250764 135410 250776
rect 273714 250764 273720 250776
rect 135404 250736 273720 250764
rect 135404 250724 135410 250736
rect 273714 250724 273720 250736
rect 273772 250724 273778 250776
rect 306926 250724 306932 250776
rect 306984 250764 306990 250776
rect 365898 250764 365904 250776
rect 306984 250736 365904 250764
rect 306984 250724 306990 250736
rect 365898 250724 365904 250736
rect 365956 250724 365962 250776
rect 70394 250656 70400 250708
rect 70452 250696 70458 250708
rect 264238 250696 264244 250708
rect 70452 250668 264244 250696
rect 70452 250656 70458 250668
rect 264238 250656 264244 250668
rect 264296 250656 264302 250708
rect 311894 250656 311900 250708
rect 311952 250696 311958 250708
rect 374086 250696 374092 250708
rect 311952 250668 374092 250696
rect 311952 250656 311958 250668
rect 374086 250656 374092 250668
rect 374144 250656 374150 250708
rect 66254 250588 66260 250640
rect 66312 250628 66318 250640
rect 262582 250628 262588 250640
rect 66312 250600 262588 250628
rect 66312 250588 66318 250600
rect 262582 250588 262588 250600
rect 262640 250588 262646 250640
rect 318886 250588 318892 250640
rect 318944 250628 318950 250640
rect 416774 250628 416780 250640
rect 318944 250600 416780 250628
rect 318944 250588 318950 250600
rect 416774 250588 416780 250600
rect 416832 250588 416838 250640
rect 62114 250520 62120 250572
rect 62172 250560 62178 250572
rect 262490 250560 262496 250572
rect 62172 250532 262496 250560
rect 62172 250520 62178 250532
rect 262490 250520 262496 250532
rect 262548 250520 262554 250572
rect 331214 250520 331220 250572
rect 331272 250560 331278 250572
rect 492674 250560 492680 250572
rect 331272 250532 492680 250560
rect 331272 250520 331278 250532
rect 492674 250520 492680 250532
rect 492732 250520 492738 250572
rect 52546 250452 52552 250504
rect 52604 250492 52610 250504
rect 260926 250492 260932 250504
rect 52604 250464 260932 250492
rect 52604 250452 52610 250464
rect 260926 250452 260932 250464
rect 260984 250452 260990 250504
rect 345014 250452 345020 250504
rect 345072 250492 345078 250504
rect 576854 250492 576860 250504
rect 345072 250464 576860 250492
rect 345072 250452 345078 250464
rect 576854 250452 576860 250464
rect 576912 250452 576918 250504
rect 309502 250384 309508 250436
rect 309560 250424 309566 250436
rect 361574 250424 361580 250436
rect 309560 250396 361580 250424
rect 309560 250384 309566 250396
rect 361574 250384 361580 250396
rect 361632 250384 361638 250436
rect 185026 249296 185032 249348
rect 185084 249336 185090 249348
rect 282178 249336 282184 249348
rect 185084 249308 282184 249336
rect 185084 249296 185090 249308
rect 282178 249296 282184 249308
rect 282236 249296 282242 249348
rect 318794 249296 318800 249348
rect 318852 249336 318858 249348
rect 414014 249336 414020 249348
rect 318852 249308 414020 249336
rect 318852 249296 318858 249308
rect 414014 249296 414020 249308
rect 414072 249296 414078 249348
rect 85574 249228 85580 249280
rect 85632 249268 85638 249280
rect 266538 249268 266544 249280
rect 85632 249240 266544 249268
rect 85632 249228 85638 249240
rect 266538 249228 266544 249240
rect 266596 249228 266602 249280
rect 338758 249228 338764 249280
rect 338816 249268 338822 249280
rect 458174 249268 458180 249280
rect 338816 249240 458180 249268
rect 338816 249228 338822 249240
rect 458174 249228 458180 249240
rect 458232 249228 458238 249280
rect 82814 249160 82820 249212
rect 82872 249200 82878 249212
rect 264974 249200 264980 249212
rect 82872 249172 264980 249200
rect 82872 249160 82878 249172
rect 264974 249160 264980 249172
rect 265032 249160 265038 249212
rect 327074 249160 327080 249212
rect 327132 249200 327138 249212
rect 460934 249200 460940 249212
rect 327132 249172 460940 249200
rect 327132 249160 327138 249172
rect 460934 249160 460940 249172
rect 460992 249160 460998 249212
rect 59354 249092 59360 249144
rect 59412 249132 59418 249144
rect 262398 249132 262404 249144
rect 59412 249104 262404 249132
rect 59412 249092 59418 249104
rect 262398 249092 262404 249104
rect 262456 249092 262462 249144
rect 328454 249092 328460 249144
rect 328512 249132 328518 249144
rect 477494 249132 477500 249144
rect 328512 249104 477500 249132
rect 328512 249092 328518 249104
rect 477494 249092 477500 249104
rect 477552 249092 477558 249144
rect 57330 249024 57336 249076
rect 57388 249064 57394 249076
rect 261386 249064 261392 249076
rect 57388 249036 261392 249064
rect 57388 249024 57394 249036
rect 261386 249024 261392 249036
rect 261444 249024 261450 249076
rect 335446 249024 335452 249076
rect 335504 249064 335510 249076
rect 520274 249064 520280 249076
rect 335504 249036 520280 249064
rect 335504 249024 335510 249036
rect 520274 249024 520280 249036
rect 520332 249024 520338 249076
rect 308122 248344 308128 248396
rect 308180 248384 308186 248396
rect 364518 248384 364524 248396
rect 308180 248356 364524 248384
rect 308180 248344 308186 248356
rect 364518 248344 364524 248356
rect 364576 248344 364582 248396
rect 305362 248276 305368 248328
rect 305420 248316 305426 248328
rect 362954 248316 362960 248328
rect 305420 248288 362960 248316
rect 305420 248276 305426 248288
rect 362954 248276 362960 248288
rect 363012 248276 363018 248328
rect 306650 248208 306656 248260
rect 306708 248248 306714 248260
rect 364426 248248 364432 248260
rect 306708 248220 364432 248248
rect 306708 248208 306714 248220
rect 364426 248208 364432 248220
rect 364484 248208 364490 248260
rect 305086 248140 305092 248192
rect 305144 248180 305150 248192
rect 363046 248180 363052 248192
rect 305144 248152 363052 248180
rect 305144 248140 305150 248152
rect 363046 248140 363052 248152
rect 363104 248140 363110 248192
rect 198734 248072 198740 248124
rect 198792 248112 198798 248124
rect 284754 248112 284760 248124
rect 198792 248084 284760 248112
rect 198792 248072 198798 248084
rect 284754 248072 284760 248084
rect 284812 248072 284818 248124
rect 302326 248072 302332 248124
rect 302384 248112 302390 248124
rect 362034 248112 362040 248124
rect 302384 248084 362040 248112
rect 302384 248072 302390 248084
rect 362034 248072 362040 248084
rect 362092 248072 362098 248124
rect 175274 248004 175280 248056
rect 175332 248044 175338 248056
rect 280246 248044 280252 248056
rect 175332 248016 280252 248044
rect 175332 248004 175338 248016
rect 280246 248004 280252 248016
rect 280304 248004 280310 248056
rect 302234 248004 302240 248056
rect 302292 248044 302298 248056
rect 371326 248044 371332 248056
rect 302292 248016 371332 248044
rect 302292 248004 302298 248016
rect 371326 248004 371332 248016
rect 371384 248004 371390 248056
rect 140774 247936 140780 247988
rect 140832 247976 140838 247988
rect 275186 247976 275192 247988
rect 140832 247948 275192 247976
rect 140832 247936 140838 247948
rect 275186 247936 275192 247948
rect 275244 247936 275250 247988
rect 320174 247936 320180 247988
rect 320232 247976 320238 247988
rect 423766 247976 423772 247988
rect 320232 247948 423772 247976
rect 320232 247936 320238 247948
rect 423766 247936 423772 247948
rect 423824 247936 423830 247988
rect 89714 247868 89720 247920
rect 89772 247908 89778 247920
rect 266446 247908 266452 247920
rect 89772 247880 266452 247908
rect 89772 247868 89778 247880
rect 266446 247868 266452 247880
rect 266504 247868 266510 247920
rect 325694 247868 325700 247920
rect 325752 247908 325758 247920
rect 455414 247908 455420 247920
rect 325752 247880 455420 247908
rect 325752 247868 325758 247880
rect 455414 247868 455420 247880
rect 455472 247868 455478 247920
rect 41414 247800 41420 247852
rect 41472 247840 41478 247852
rect 258626 247840 258632 247852
rect 41472 247812 258632 247840
rect 41472 247800 41478 247812
rect 258626 247800 258632 247812
rect 258684 247800 258690 247852
rect 332594 247800 332600 247852
rect 332652 247840 332658 247852
rect 502334 247840 502340 247852
rect 332652 247812 502340 247840
rect 332652 247800 332658 247812
rect 502334 247800 502340 247812
rect 502392 247800 502398 247852
rect 35158 247732 35164 247784
rect 35216 247772 35222 247784
rect 256786 247772 256792 247784
rect 35216 247744 256792 247772
rect 35216 247732 35222 247744
rect 256786 247732 256792 247744
rect 256844 247732 256850 247784
rect 334434 247732 334440 247784
rect 334492 247772 334498 247784
rect 511994 247772 512000 247784
rect 334492 247744 512000 247772
rect 334492 247732 334498 247744
rect 511994 247732 512000 247744
rect 512052 247732 512058 247784
rect 8938 247664 8944 247716
rect 8996 247704 9002 247716
rect 252646 247704 252652 247716
rect 8996 247676 252652 247704
rect 8996 247664 9002 247676
rect 252646 247664 252652 247676
rect 252704 247664 252710 247716
rect 336734 247664 336740 247716
rect 336792 247704 336798 247716
rect 524414 247704 524420 247716
rect 336792 247676 524420 247704
rect 336792 247664 336798 247676
rect 524414 247664 524420 247676
rect 524472 247664 524478 247716
rect 309410 247596 309416 247648
rect 309468 247636 309474 247648
rect 364610 247636 364616 247648
rect 309468 247608 364616 247636
rect 309468 247596 309474 247608
rect 364610 247596 364616 247608
rect 364668 247596 364674 247648
rect 355686 247528 355692 247580
rect 355744 247568 355750 247580
rect 369946 247568 369952 247580
rect 355744 247540 369952 247568
rect 355744 247528 355750 247540
rect 369946 247528 369952 247540
rect 370004 247528 370010 247580
rect 217318 246712 217324 246764
rect 217376 246752 217382 246764
rect 346394 246752 346400 246764
rect 217376 246724 346400 246752
rect 217376 246712 217382 246724
rect 346394 246712 346400 246724
rect 346452 246712 346458 246764
rect 121454 246644 121460 246696
rect 121512 246684 121518 246696
rect 272334 246684 272340 246696
rect 121512 246656 272340 246684
rect 121512 246644 121518 246656
rect 272334 246644 272340 246656
rect 272392 246644 272398 246696
rect 300854 246644 300860 246696
rect 300912 246684 300918 246696
rect 366082 246684 366088 246696
rect 300912 246656 366088 246684
rect 300912 246644 300918 246656
rect 366082 246644 366088 246656
rect 366140 246644 366146 246696
rect 109034 246576 109040 246628
rect 109092 246616 109098 246628
rect 269206 246616 269212 246628
rect 109092 246588 269212 246616
rect 109092 246576 109098 246588
rect 269206 246576 269212 246588
rect 269264 246576 269270 246628
rect 322934 246576 322940 246628
rect 322992 246616 322998 246628
rect 438854 246616 438860 246628
rect 322992 246588 438860 246616
rect 322992 246576 322998 246588
rect 438854 246576 438860 246588
rect 438912 246576 438918 246628
rect 85666 246508 85672 246560
rect 85724 246548 85730 246560
rect 266906 246548 266912 246560
rect 85724 246520 266912 246548
rect 85724 246508 85730 246520
rect 266906 246508 266912 246520
rect 266964 246508 266970 246560
rect 334342 246508 334348 246560
rect 334400 246548 334406 246560
rect 505094 246548 505100 246560
rect 334400 246520 505100 246548
rect 334400 246508 334406 246520
rect 505094 246508 505100 246520
rect 505152 246508 505158 246560
rect 64874 246440 64880 246492
rect 64932 246480 64938 246492
rect 262306 246480 262312 246492
rect 64932 246452 262312 246480
rect 64932 246440 64938 246452
rect 262306 246440 262312 246452
rect 262364 246440 262370 246492
rect 334250 246440 334256 246492
rect 334308 246480 334314 246492
rect 507854 246480 507860 246492
rect 334308 246452 507860 246480
rect 334308 246440 334314 246452
rect 507854 246440 507860 246452
rect 507912 246440 507918 246492
rect 38654 246372 38660 246424
rect 38712 246412 38718 246424
rect 250438 246412 250444 246424
rect 38712 246384 250444 246412
rect 38712 246372 38718 246384
rect 250438 246372 250444 246384
rect 250496 246372 250502 246424
rect 334158 246372 334164 246424
rect 334216 246412 334222 246424
rect 510614 246412 510620 246424
rect 334216 246384 510620 246412
rect 334216 246372 334222 246384
rect 510614 246372 510620 246384
rect 510672 246372 510678 246424
rect 6914 246304 6920 246356
rect 6972 246344 6978 246356
rect 252922 246344 252928 246356
rect 6972 246316 252928 246344
rect 6972 246304 6978 246316
rect 252922 246304 252928 246316
rect 252980 246304 252986 246356
rect 335354 246304 335360 246356
rect 335412 246344 335418 246356
rect 516134 246344 516140 246356
rect 335412 246316 516140 246344
rect 335412 246304 335418 246316
rect 516134 246304 516140 246316
rect 516192 246304 516198 246356
rect 355594 245556 355600 245608
rect 355652 245596 355658 245608
rect 369854 245596 369860 245608
rect 355652 245568 369860 245596
rect 355652 245556 355658 245568
rect 369854 245556 369860 245568
rect 369912 245556 369918 245608
rect 355502 245488 355508 245540
rect 355560 245528 355566 245540
rect 372706 245528 372712 245540
rect 355560 245500 372712 245528
rect 355560 245488 355566 245500
rect 372706 245488 372712 245500
rect 372764 245488 372770 245540
rect 307846 245420 307852 245472
rect 307904 245460 307910 245472
rect 361758 245460 361764 245472
rect 307904 245432 361764 245460
rect 307904 245420 307910 245432
rect 361758 245420 361764 245432
rect 361816 245420 361822 245472
rect 307938 245352 307944 245404
rect 307996 245392 308002 245404
rect 361850 245392 361856 245404
rect 307996 245364 361856 245392
rect 307996 245352 308002 245364
rect 361850 245352 361856 245364
rect 361908 245352 361914 245404
rect 203610 245284 203616 245336
rect 203668 245324 203674 245336
rect 283374 245324 283380 245336
rect 203668 245296 283380 245324
rect 203668 245284 203674 245296
rect 283374 245284 283380 245296
rect 283432 245284 283438 245336
rect 307754 245284 307760 245336
rect 307812 245324 307818 245336
rect 361666 245324 361672 245336
rect 307812 245296 361672 245324
rect 307812 245284 307818 245296
rect 361666 245284 361672 245296
rect 361724 245284 361730 245336
rect 171226 245216 171232 245268
rect 171284 245256 171290 245268
rect 280706 245256 280712 245268
rect 171284 245228 280712 245256
rect 171284 245216 171290 245228
rect 280706 245216 280712 245228
rect 280764 245216 280770 245268
rect 306374 245216 306380 245268
rect 306432 245256 306438 245268
rect 361942 245256 361948 245268
rect 306432 245228 361948 245256
rect 306432 245216 306438 245228
rect 361942 245216 361948 245228
rect 362000 245216 362006 245268
rect 168466 245148 168472 245200
rect 168524 245188 168530 245200
rect 279234 245188 279240 245200
rect 168524 245160 279240 245188
rect 168524 245148 168530 245160
rect 279234 245148 279240 245160
rect 279292 245148 279298 245200
rect 324314 245148 324320 245200
rect 324372 245188 324378 245200
rect 445754 245188 445760 245200
rect 324372 245160 445760 245188
rect 324372 245148 324378 245160
rect 445754 245148 445760 245160
rect 445812 245148 445818 245200
rect 104894 245080 104900 245132
rect 104952 245120 104958 245132
rect 269666 245120 269672 245132
rect 104952 245092 269672 245120
rect 104952 245080 104958 245092
rect 269666 245080 269672 245092
rect 269724 245080 269730 245132
rect 334066 245080 334072 245132
rect 334124 245120 334130 245132
rect 503714 245120 503720 245132
rect 334124 245092 503720 245120
rect 334124 245080 334130 245092
rect 503714 245080 503720 245092
rect 503772 245080 503778 245132
rect 100754 245012 100760 245064
rect 100812 245052 100818 245064
rect 268286 245052 268292 245064
rect 100812 245024 268292 245052
rect 100812 245012 100818 245024
rect 268286 245012 268292 245024
rect 268344 245012 268350 245064
rect 333974 245012 333980 245064
rect 334032 245052 334038 245064
rect 506566 245052 506572 245064
rect 334032 245024 506572 245052
rect 334032 245012 334038 245024
rect 506566 245012 506572 245024
rect 506624 245012 506630 245064
rect 60826 244944 60832 244996
rect 60884 244984 60890 244996
rect 262674 244984 262680 244996
rect 60884 244956 262680 244984
rect 60884 244944 60890 244956
rect 262674 244944 262680 244956
rect 262732 244944 262738 244996
rect 338114 244944 338120 244996
rect 338172 244984 338178 244996
rect 534074 244984 534080 244996
rect 338172 244956 534080 244984
rect 338172 244944 338178 244956
rect 534074 244944 534080 244956
rect 534132 244944 534138 244996
rect 27706 244876 27712 244928
rect 27764 244916 27770 244928
rect 257246 244916 257252 244928
rect 27764 244888 257252 244916
rect 27764 244876 27770 244888
rect 257246 244876 257252 244888
rect 257304 244876 257310 244928
rect 343634 244876 343640 244928
rect 343692 244916 343698 244928
rect 571334 244916 571340 244928
rect 343692 244888 571340 244916
rect 343692 244876 343698 244888
rect 571334 244876 571340 244888
rect 571392 244876 571398 244928
rect 355318 244468 355324 244520
rect 355376 244508 355382 244520
rect 363414 244508 363420 244520
rect 355376 244480 363420 244508
rect 355376 244468 355382 244480
rect 363414 244468 363420 244480
rect 363472 244468 363478 244520
rect 355410 244264 355416 244316
rect 355468 244304 355474 244316
rect 363782 244304 363788 244316
rect 355468 244276 363788 244304
rect 355468 244264 355474 244276
rect 363782 244264 363788 244276
rect 363840 244264 363846 244316
rect 303614 243856 303620 243908
rect 303672 243896 303678 243908
rect 364702 243896 364708 243908
rect 303672 243868 364708 243896
rect 303672 243856 303678 243868
rect 364702 243856 364708 243868
rect 364760 243856 364766 243908
rect 299658 243788 299664 243840
rect 299716 243828 299722 243840
rect 362218 243828 362224 243840
rect 299716 243800 362224 243828
rect 299716 243788 299722 243800
rect 362218 243788 362224 243800
rect 362276 243788 362282 243840
rect 299750 243720 299756 243772
rect 299808 243760 299814 243772
rect 362402 243760 362408 243772
rect 299808 243732 362408 243760
rect 299808 243720 299814 243732
rect 362402 243720 362408 243732
rect 362460 243720 362466 243772
rect 298186 243652 298192 243704
rect 298244 243692 298250 243704
rect 361022 243692 361028 243704
rect 298244 243664 361028 243692
rect 298244 243652 298250 243664
rect 361022 243652 361028 243664
rect 361080 243652 361086 243704
rect 219342 243584 219348 243636
rect 219400 243624 219406 243636
rect 297174 243624 297180 243636
rect 219400 243596 297180 243624
rect 219400 243584 219406 243596
rect 297174 243584 297180 243596
rect 297232 243584 297238 243636
rect 299474 243584 299480 243636
rect 299532 243624 299538 243636
rect 366542 243624 366548 243636
rect 299532 243596 366548 243624
rect 299532 243584 299538 243596
rect 366542 243584 366548 243596
rect 366600 243584 366606 243636
rect 217410 243516 217416 243568
rect 217468 243556 217474 243568
rect 297266 243556 297272 243568
rect 217468 243528 297272 243556
rect 217468 243516 217474 243528
rect 297266 243516 297272 243528
rect 297324 243516 297330 243568
rect 299566 243516 299572 243568
rect 299624 243556 299630 243568
rect 369302 243556 369308 243568
rect 299624 243528 369308 243556
rect 299624 243516 299630 243528
rect 369302 243516 369308 243528
rect 369360 243516 369366 243568
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 215938 215268 215944 215280
rect 3384 215240 215944 215268
rect 3384 215228 3390 215240
rect 215938 215228 215944 215240
rect 215996 215228 216002 215280
rect 214374 213868 214380 213920
rect 214432 213908 214438 213920
rect 215938 213908 215944 213920
rect 214432 213880 215944 213908
rect 214432 213868 214438 213880
rect 215938 213868 215944 213880
rect 215996 213868 216002 213920
rect 373350 206932 373356 206984
rect 373408 206972 373414 206984
rect 579614 206972 579620 206984
rect 373408 206944 579620 206972
rect 373408 206932 373414 206944
rect 579614 206932 579620 206944
rect 579672 206932 579678 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 196710 202824 196716 202836
rect 3108 202796 196716 202824
rect 3108 202784 3114 202796
rect 196710 202784 196716 202796
rect 196768 202784 196774 202836
rect 215754 195372 215760 195424
rect 215812 195412 215818 195424
rect 217686 195412 217692 195424
rect 215812 195384 217692 195412
rect 215812 195372 215818 195384
rect 217686 195372 217692 195384
rect 217744 195372 217750 195424
rect 577590 193128 577596 193180
rect 577648 193168 577654 193180
rect 580810 193168 580816 193180
rect 577648 193140 580816 193168
rect 577648 193128 577654 193140
rect 580810 193128 580816 193140
rect 580868 193128 580874 193180
rect 371970 166948 371976 167000
rect 372028 166988 372034 167000
rect 580166 166988 580172 167000
rect 372028 166960 580172 166988
rect 372028 166948 372034 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 358354 160080 358360 160132
rect 358412 160120 358418 160132
rect 363782 160120 363788 160132
rect 358412 160092 363788 160120
rect 358412 160080 358418 160092
rect 363782 160080 363788 160092
rect 363840 160080 363846 160132
rect 322934 159604 322940 159656
rect 322992 159644 322998 159656
rect 358170 159644 358176 159656
rect 322992 159616 358176 159644
rect 322992 159604 322998 159616
rect 358170 159604 358176 159616
rect 358228 159604 358234 159656
rect 318702 159536 318708 159588
rect 318760 159576 318766 159588
rect 358078 159576 358084 159588
rect 318760 159548 358084 159576
rect 318760 159536 318766 159548
rect 358078 159536 358084 159548
rect 358136 159536 358142 159588
rect 213638 159468 213644 159520
rect 213696 159508 213702 159520
rect 256694 159508 256700 159520
rect 213696 159480 256700 159508
rect 213696 159468 213702 159480
rect 256694 159468 256700 159480
rect 256752 159468 256758 159520
rect 314654 159468 314660 159520
rect 314712 159508 314718 159520
rect 357802 159508 357808 159520
rect 314712 159480 357808 159508
rect 314712 159468 314718 159480
rect 357802 159468 357808 159480
rect 357860 159468 357866 159520
rect 211706 159400 211712 159452
rect 211764 159440 211770 159452
rect 259454 159440 259460 159452
rect 211764 159412 259460 159440
rect 211764 159400 211770 159412
rect 259454 159400 259460 159412
rect 259512 159400 259518 159452
rect 310422 159400 310428 159452
rect 310480 159440 310486 159452
rect 357986 159440 357992 159452
rect 310480 159412 357992 159440
rect 310480 159400 310486 159412
rect 357986 159400 357992 159412
rect 358044 159400 358050 159452
rect 215846 159332 215852 159384
rect 215904 159372 215910 159384
rect 263686 159372 263692 159384
rect 215904 159344 263692 159372
rect 215904 159332 215910 159344
rect 263686 159332 263692 159344
rect 263744 159332 263750 159384
rect 304994 159332 305000 159384
rect 305052 159372 305058 159384
rect 356698 159372 356704 159384
rect 305052 159344 356704 159372
rect 305052 159332 305058 159344
rect 356698 159332 356704 159344
rect 356756 159332 356762 159384
rect 300946 159196 300952 159248
rect 301004 159236 301010 159248
rect 357894 159236 357900 159248
rect 301004 159208 357900 159236
rect 301004 159196 301010 159208
rect 357894 159196 357900 159208
rect 357952 159196 357958 159248
rect 295886 159128 295892 159180
rect 295944 159168 295950 159180
rect 370682 159168 370688 159180
rect 295944 159140 370688 159168
rect 295944 159128 295950 159140
rect 370682 159128 370688 159140
rect 370740 159128 370746 159180
rect 288342 159060 288348 159112
rect 288400 159100 288406 159112
rect 365070 159100 365076 159112
rect 288400 159072 365076 159100
rect 288400 159060 288406 159072
rect 365070 159060 365076 159072
rect 365128 159060 365134 159112
rect 279234 158992 279240 159044
rect 279292 159032 279298 159044
rect 360838 159032 360844 159044
rect 279292 159004 360844 159032
rect 279292 158992 279298 159004
rect 360838 158992 360844 159004
rect 360896 158992 360902 159044
rect 278130 158924 278136 158976
rect 278188 158964 278194 158976
rect 360746 158964 360752 158976
rect 278188 158936 360752 158964
rect 278188 158924 278194 158936
rect 360746 158924 360752 158936
rect 360804 158924 360810 158976
rect 277026 158856 277032 158908
rect 277084 158896 277090 158908
rect 360654 158896 360660 158908
rect 277084 158868 360660 158896
rect 277084 158856 277090 158868
rect 360654 158856 360660 158868
rect 360712 158856 360718 158908
rect 275830 158788 275836 158840
rect 275888 158828 275894 158840
rect 359366 158828 359372 158840
rect 275888 158800 359372 158828
rect 275888 158788 275894 158800
rect 359366 158788 359372 158800
rect 359424 158788 359430 158840
rect 211890 158720 211896 158772
rect 211948 158760 211954 158772
rect 239582 158760 239588 158772
rect 211948 158732 239588 158760
rect 211948 158720 211954 158732
rect 239582 158720 239588 158732
rect 239640 158720 239646 158772
rect 274450 158720 274456 158772
rect 274508 158760 274514 158772
rect 359458 158760 359464 158772
rect 274508 158732 359464 158760
rect 274508 158720 274514 158732
rect 359458 158720 359464 158732
rect 359516 158720 359522 158772
rect 213270 158652 213276 158704
rect 213328 158692 213334 158704
rect 238110 158692 238116 158704
rect 213328 158664 238116 158692
rect 213328 158652 213334 158664
rect 238110 158652 238116 158664
rect 238168 158652 238174 158704
rect 298554 158652 298560 158704
rect 298612 158692 298618 158704
rect 304994 158692 305000 158704
rect 298612 158664 305000 158692
rect 298612 158652 298618 158664
rect 304994 158652 305000 158664
rect 305052 158652 305058 158704
rect 306098 158652 306104 158704
rect 306156 158692 306162 158704
rect 314654 158692 314660 158704
rect 306156 158664 314660 158692
rect 306156 158652 306162 158664
rect 314654 158652 314660 158664
rect 314712 158652 314718 158704
rect 212074 158584 212080 158636
rect 212132 158624 212138 158636
rect 230474 158624 230480 158636
rect 212132 158596 230480 158624
rect 212132 158584 212138 158596
rect 230474 158584 230480 158596
rect 230532 158584 230538 158636
rect 308766 158584 308772 158636
rect 308824 158624 308830 158636
rect 318702 158624 318708 158636
rect 308824 158596 318708 158624
rect 308824 158584 308830 158596
rect 318702 158584 318708 158596
rect 318760 158584 318766 158636
rect 214834 158516 214840 158568
rect 214892 158556 214898 158568
rect 235994 158556 236000 158568
rect 214892 158528 236000 158556
rect 214892 158516 214898 158528
rect 235994 158516 236000 158528
rect 236052 158516 236058 158568
rect 262858 158516 262864 158568
rect 262916 158556 262922 158568
rect 367738 158556 367744 158568
rect 262916 158528 367744 158556
rect 262916 158516 262922 158528
rect 367738 158516 367744 158528
rect 367796 158516 367802 158568
rect 213362 158448 213368 158500
rect 213420 158488 213426 158500
rect 234706 158488 234712 158500
rect 213420 158460 234712 158488
rect 213420 158448 213426 158460
rect 234706 158448 234712 158460
rect 234764 158448 234770 158500
rect 259546 158448 259552 158500
rect 259604 158488 259610 158500
rect 364794 158488 364800 158500
rect 259604 158460 364800 158488
rect 259604 158448 259610 158460
rect 364794 158448 364800 158460
rect 364852 158448 364858 158500
rect 219066 158380 219072 158432
rect 219124 158420 219130 158432
rect 242986 158420 242992 158432
rect 219124 158392 242992 158420
rect 219124 158380 219130 158392
rect 242986 158380 242992 158392
rect 243044 158380 243050 158432
rect 263594 158380 263600 158432
rect 263652 158420 263658 158432
rect 362310 158420 362316 158432
rect 263652 158392 362316 158420
rect 263652 158380 263658 158392
rect 362310 158380 362316 158392
rect 362368 158380 362374 158432
rect 214558 158312 214564 158364
rect 214616 158352 214622 158364
rect 242894 158352 242900 158364
rect 214616 158324 242900 158352
rect 214616 158312 214622 158324
rect 242894 158312 242900 158324
rect 242952 158312 242958 158364
rect 268746 158312 268752 158364
rect 268804 158352 268810 158364
rect 357710 158352 357716 158364
rect 268804 158324 357716 158352
rect 268804 158312 268810 158324
rect 357710 158312 357716 158324
rect 357768 158312 357774 158364
rect 214926 158244 214932 158296
rect 214984 158284 214990 158296
rect 245654 158284 245660 158296
rect 214984 158256 245660 158284
rect 214984 158244 214990 158256
rect 245654 158244 245660 158256
rect 245712 158244 245718 158296
rect 269850 158244 269856 158296
rect 269908 158284 269914 158296
rect 357526 158284 357532 158296
rect 269908 158256 357532 158284
rect 269908 158244 269914 158256
rect 357526 158244 357532 158256
rect 357584 158244 357590 158296
rect 216214 158176 216220 158228
rect 216272 158216 216278 158228
rect 247034 158216 247040 158228
rect 216272 158188 247040 158216
rect 216272 158176 216278 158188
rect 247034 158176 247040 158188
rect 247092 158176 247098 158228
rect 271138 158176 271144 158228
rect 271196 158216 271202 158228
rect 357618 158216 357624 158228
rect 271196 158188 357624 158216
rect 271196 158176 271202 158188
rect 357618 158176 357624 158188
rect 357676 158176 357682 158228
rect 217962 158108 217968 158160
rect 218020 158148 218026 158160
rect 251174 158148 251180 158160
rect 218020 158120 251180 158148
rect 218020 158108 218026 158120
rect 251174 158108 251180 158120
rect 251232 158108 251238 158160
rect 303522 158108 303528 158160
rect 303580 158148 303586 158160
rect 310422 158148 310428 158160
rect 303580 158120 310428 158148
rect 303580 158108 303586 158120
rect 310422 158108 310428 158120
rect 310480 158108 310486 158160
rect 321002 158108 321008 158160
rect 321060 158148 321066 158160
rect 360562 158148 360568 158160
rect 321060 158120 360568 158148
rect 321060 158108 321066 158120
rect 360562 158108 360568 158120
rect 360620 158108 360626 158160
rect 219158 158040 219164 158092
rect 219216 158080 219222 158092
rect 252554 158080 252560 158092
rect 219216 158052 252560 158080
rect 219216 158040 219222 158052
rect 252554 158040 252560 158052
rect 252612 158040 252618 158092
rect 313458 158040 313464 158092
rect 313516 158080 313522 158092
rect 359090 158080 359096 158092
rect 313516 158052 359096 158080
rect 313516 158040 313522 158052
rect 359090 158040 359096 158052
rect 359148 158040 359154 158092
rect 216306 157972 216312 158024
rect 216364 158012 216370 158024
rect 249794 158012 249800 158024
rect 216364 157984 249800 158012
rect 216364 157972 216370 157984
rect 249794 157972 249800 157984
rect 249852 157972 249858 158024
rect 315850 157972 315856 158024
rect 315908 158012 315914 158024
rect 359274 158012 359280 158024
rect 315908 157984 359280 158012
rect 315908 157972 315914 157984
rect 359274 157972 359280 157984
rect 359332 157972 359338 158024
rect 216122 157904 216128 157956
rect 216180 157944 216186 157956
rect 233234 157944 233240 157956
rect 216180 157916 233240 157944
rect 216180 157904 216186 157916
rect 233234 157904 233240 157916
rect 233292 157904 233298 157956
rect 318610 157904 318616 157956
rect 318668 157944 318674 157956
rect 359182 157944 359188 157956
rect 318668 157916 359188 157944
rect 318668 157904 318674 157916
rect 359182 157904 359188 157916
rect 359240 157904 359246 157956
rect 218974 157836 218980 157888
rect 219032 157876 219038 157888
rect 234614 157876 234620 157888
rect 219032 157848 234620 157876
rect 219032 157836 219038 157848
rect 234614 157836 234620 157848
rect 234672 157836 234678 157888
rect 272242 157836 272248 157888
rect 272300 157876 272306 157888
rect 322934 157876 322940 157888
rect 272300 157848 322940 157876
rect 272300 157836 272306 157848
rect 322934 157836 322940 157848
rect 322992 157836 322998 157888
rect 323394 157836 323400 157888
rect 323452 157876 323458 157888
rect 360378 157876 360384 157888
rect 323452 157848 360384 157876
rect 323452 157836 323458 157848
rect 360378 157836 360384 157848
rect 360436 157836 360442 157888
rect 214650 157768 214656 157820
rect 214708 157808 214714 157820
rect 229094 157808 229100 157820
rect 214708 157780 229100 157808
rect 214708 157768 214714 157780
rect 229094 157768 229100 157780
rect 229152 157768 229158 157820
rect 325970 157768 325976 157820
rect 326028 157808 326034 157820
rect 360470 157808 360476 157820
rect 326028 157780 360476 157808
rect 326028 157768 326034 157780
rect 360470 157768 360476 157780
rect 360528 157768 360534 157820
rect 240686 157700 240692 157752
rect 240744 157740 240750 157752
rect 372982 157740 372988 157752
rect 240744 157712 372988 157740
rect 240744 157700 240750 157712
rect 372982 157700 372988 157712
rect 373040 157700 373046 157752
rect 261478 157632 261484 157684
rect 261536 157672 261542 157684
rect 366450 157672 366456 157684
rect 261536 157644 366456 157672
rect 261536 157632 261542 157644
rect 366450 157632 366456 157644
rect 366508 157632 366514 157684
rect 248322 157292 248328 157344
rect 248380 157332 248386 157344
rect 370406 157332 370412 157344
rect 248380 157304 370412 157332
rect 248380 157292 248386 157304
rect 370406 157292 370412 157304
rect 370464 157292 370470 157344
rect 252370 157224 252376 157276
rect 252428 157264 252434 157276
rect 369118 157264 369124 157276
rect 252428 157236 369124 157264
rect 252428 157224 252434 157236
rect 369118 157224 369124 157236
rect 369176 157224 369182 157276
rect 250438 157156 250444 157208
rect 250496 157196 250502 157208
rect 366358 157196 366364 157208
rect 250496 157168 366364 157196
rect 250496 157156 250502 157168
rect 366358 157156 366364 157168
rect 366416 157156 366422 157208
rect 254946 157088 254952 157140
rect 255004 157128 255010 157140
rect 363506 157128 363512 157140
rect 255004 157100 363512 157128
rect 255004 157088 255010 157100
rect 363506 157088 363512 157100
rect 363564 157088 363570 157140
rect 257246 157020 257252 157072
rect 257304 157060 257310 157072
rect 366174 157060 366180 157072
rect 257304 157032 366180 157060
rect 257304 157020 257310 157032
rect 366174 157020 366180 157032
rect 366232 157020 366238 157072
rect 259086 156952 259092 157004
rect 259144 156992 259150 157004
rect 366266 156992 366272 157004
rect 259144 156964 366272 156992
rect 259144 156952 259150 156964
rect 366266 156952 366272 156964
rect 366324 156952 366330 157004
rect 255866 156884 255872 156936
rect 255924 156924 255930 156936
rect 360930 156924 360936 156936
rect 255924 156896 360936 156924
rect 255924 156884 255930 156896
rect 360930 156884 360936 156896
rect 360988 156884 360994 156936
rect 271046 156816 271052 156868
rect 271104 156856 271110 156868
rect 374178 156856 374184 156868
rect 271104 156828 374184 156856
rect 271104 156816 271110 156828
rect 374178 156816 374184 156828
rect 374236 156816 374242 156868
rect 276106 156748 276112 156800
rect 276164 156788 276170 156800
rect 369026 156788 369032 156800
rect 276164 156760 369032 156788
rect 276164 156748 276170 156760
rect 369026 156748 369032 156760
rect 369084 156748 369090 156800
rect 281350 156680 281356 156732
rect 281408 156720 281414 156732
rect 371694 156720 371700 156732
rect 281408 156692 371700 156720
rect 281408 156680 281414 156692
rect 371694 156680 371700 156692
rect 371752 156680 371758 156732
rect 286318 156612 286324 156664
rect 286376 156652 286382 156664
rect 371786 156652 371792 156664
rect 286376 156624 371792 156652
rect 286376 156612 286382 156624
rect 371786 156612 371792 156624
rect 371844 156612 371850 156664
rect 274450 156544 274456 156596
rect 274508 156584 274514 156596
rect 358906 156584 358912 156596
rect 274508 156556 358912 156584
rect 274508 156544 274514 156556
rect 358906 156544 358912 156556
rect 358964 156544 358970 156596
rect 293678 156476 293684 156528
rect 293736 156516 293742 156528
rect 371602 156516 371608 156528
rect 293736 156488 371608 156516
rect 293736 156476 293742 156488
rect 371602 156476 371608 156488
rect 371660 156476 371666 156528
rect 311066 156408 311072 156460
rect 311124 156448 311130 156460
rect 358998 156448 359004 156460
rect 311124 156420 359004 156448
rect 311124 156408 311130 156420
rect 358998 156408 359004 156420
rect 359056 156408 359062 156460
rect 248690 155864 248696 155916
rect 248748 155904 248754 155916
rect 368842 155904 368848 155916
rect 248748 155876 368848 155904
rect 248748 155864 248754 155876
rect 368842 155864 368848 155876
rect 368900 155864 368906 155916
rect 211982 155796 211988 155848
rect 212040 155836 212046 155848
rect 237374 155836 237380 155848
rect 212040 155808 237380 155836
rect 212040 155796 212046 155808
rect 237374 155796 237380 155808
rect 237432 155796 237438 155848
rect 252278 155796 252284 155848
rect 252336 155836 252342 155848
rect 370222 155836 370228 155848
rect 252336 155808 370228 155836
rect 252336 155796 252342 155808
rect 370222 155796 370228 155808
rect 370280 155796 370286 155848
rect 213546 155728 213552 155780
rect 213604 155768 213610 155780
rect 241514 155768 241520 155780
rect 213604 155740 241520 155768
rect 213604 155728 213610 155740
rect 241514 155728 241520 155740
rect 241572 155728 241578 155780
rect 253566 155728 253572 155780
rect 253624 155768 253630 155780
rect 363598 155768 363604 155780
rect 253624 155740 363604 155768
rect 253624 155728 253630 155740
rect 363598 155728 363604 155740
rect 363656 155728 363662 155780
rect 216030 155660 216036 155712
rect 216088 155700 216094 155712
rect 248414 155700 248420 155712
rect 216088 155672 248420 155700
rect 216088 155660 216094 155672
rect 248414 155660 248420 155672
rect 248472 155660 248478 155712
rect 260650 155660 260656 155712
rect 260708 155700 260714 155712
rect 367278 155700 367284 155712
rect 260708 155672 367284 155700
rect 260708 155660 260714 155672
rect 367278 155660 367284 155672
rect 367336 155660 367342 155712
rect 213454 155592 213460 155644
rect 213512 155632 213518 155644
rect 253934 155632 253940 155644
rect 213512 155604 253940 155632
rect 213512 155592 213518 155604
rect 253934 155592 253940 155604
rect 253992 155592 253998 155644
rect 261754 155592 261760 155644
rect 261812 155632 261818 155644
rect 367462 155632 367468 155644
rect 261812 155604 367468 155632
rect 261812 155592 261818 155604
rect 367462 155592 367468 155604
rect 367520 155592 367526 155644
rect 210694 155524 210700 155576
rect 210752 155564 210758 155576
rect 267826 155564 267832 155576
rect 210752 155536 267832 155564
rect 210752 155524 210758 155536
rect 267826 155524 267832 155536
rect 267884 155524 267890 155576
rect 268930 155524 268936 155576
rect 268988 155564 268994 155576
rect 372798 155564 372804 155576
rect 268988 155536 372804 155564
rect 268988 155524 268994 155536
rect 372798 155524 372804 155536
rect 372856 155524 372862 155576
rect 210878 155456 210884 155508
rect 210936 155496 210942 155508
rect 255314 155496 255320 155508
rect 210936 155468 255320 155496
rect 210936 155456 210942 155468
rect 255314 155456 255320 155468
rect 255372 155456 255378 155508
rect 264514 155456 264520 155508
rect 264572 155496 264578 155508
rect 367554 155496 367560 155508
rect 264572 155468 367560 155496
rect 264572 155456 264578 155468
rect 367554 155456 367560 155468
rect 367612 155456 367618 155508
rect 219250 155388 219256 155440
rect 219308 155428 219314 155440
rect 264974 155428 264980 155440
rect 219308 155400 264980 155428
rect 219308 155388 219314 155400
rect 264974 155388 264980 155400
rect 265032 155388 265038 155440
rect 266906 155388 266912 155440
rect 266964 155428 266970 155440
rect 370038 155428 370044 155440
rect 266964 155400 370044 155428
rect 266964 155388 266970 155400
rect 370038 155388 370044 155400
rect 370096 155388 370102 155440
rect 214466 155320 214472 155372
rect 214524 155360 214530 155372
rect 260834 155360 260840 155372
rect 214524 155332 260840 155360
rect 214524 155320 214530 155332
rect 260834 155320 260840 155332
rect 260892 155320 260898 155372
rect 265986 155320 265992 155372
rect 266044 155360 266050 155372
rect 367370 155360 367376 155372
rect 266044 155332 367376 155360
rect 266044 155320 266050 155332
rect 367370 155320 367376 155332
rect 367428 155320 367434 155372
rect 218790 155252 218796 155304
rect 218848 155292 218854 155304
rect 266354 155292 266360 155304
rect 218848 155264 266360 155292
rect 218848 155252 218854 155264
rect 266354 155252 266360 155264
rect 266412 155252 266418 155304
rect 267642 155252 267648 155304
rect 267700 155292 267706 155304
rect 368566 155292 368572 155304
rect 267700 155264 368572 155292
rect 267700 155252 267706 155264
rect 368566 155252 368572 155264
rect 368624 155252 368630 155304
rect 212166 155184 212172 155236
rect 212224 155224 212230 155236
rect 273254 155224 273260 155236
rect 212224 155196 273260 155224
rect 212224 155184 212230 155196
rect 273254 155184 273260 155196
rect 273312 155184 273318 155236
rect 274542 155184 274548 155236
rect 274600 155224 274606 155236
rect 368750 155224 368756 155236
rect 274600 155196 368756 155224
rect 274600 155184 274606 155196
rect 368750 155184 368756 155196
rect 368808 155184 368814 155236
rect 217686 155116 217692 155168
rect 217744 155156 217750 155168
rect 277394 155156 277400 155168
rect 217744 155128 277400 155156
rect 217744 155116 217750 155128
rect 277394 155116 277400 155128
rect 277452 155116 277458 155168
rect 278682 155116 278688 155168
rect 278740 155156 278746 155168
rect 368934 155156 368940 155168
rect 278740 155128 368940 155156
rect 278740 155116 278746 155128
rect 368934 155116 368940 155128
rect 368992 155116 368998 155168
rect 217410 155048 217416 155100
rect 217468 155088 217474 155100
rect 278774 155088 278780 155100
rect 217468 155060 278780 155088
rect 217468 155048 217474 155060
rect 278774 155048 278780 155060
rect 278832 155048 278838 155100
rect 283926 155048 283932 155100
rect 283984 155088 283990 155100
rect 371510 155088 371516 155100
rect 283984 155060 371516 155088
rect 283984 155048 283990 155060
rect 371510 155048 371516 155060
rect 371568 155048 371574 155100
rect 217870 154980 217876 155032
rect 217928 155020 217934 155032
rect 274634 155020 274640 155032
rect 217928 154992 274640 155020
rect 217928 154980 217934 154992
rect 274634 154980 274640 154992
rect 274692 154980 274698 155032
rect 291010 154980 291016 155032
rect 291068 155020 291074 155032
rect 372062 155020 372068 155032
rect 291068 154992 372068 155020
rect 291068 154980 291074 154992
rect 372062 154980 372068 154992
rect 372120 154980 372126 155032
rect 253658 154504 253664 154556
rect 253716 154544 253722 154556
rect 371418 154544 371424 154556
rect 253716 154516 371424 154544
rect 253716 154504 253722 154516
rect 371418 154504 371424 154516
rect 371476 154504 371482 154556
rect 256234 154436 256240 154488
rect 256292 154476 256298 154488
rect 359550 154476 359556 154488
rect 256292 154448 359556 154476
rect 256292 154436 256298 154448
rect 359550 154436 359556 154448
rect 359608 154436 359614 154488
rect 345750 154232 345756 154284
rect 345808 154272 345814 154284
rect 366542 154272 366548 154284
rect 345808 154244 366548 154272
rect 345808 154232 345814 154244
rect 366542 154232 366548 154244
rect 366600 154232 366606 154284
rect 295334 154164 295340 154216
rect 295392 154204 295398 154216
rect 362218 154204 362224 154216
rect 295392 154176 362224 154204
rect 295392 154164 295398 154176
rect 362218 154164 362224 154176
rect 362276 154164 362282 154216
rect 299566 154096 299572 154148
rect 299624 154136 299630 154148
rect 370498 154136 370504 154148
rect 299624 154108 370504 154136
rect 299624 154096 299630 154108
rect 370498 154096 370504 154108
rect 370556 154096 370562 154148
rect 288434 154028 288440 154080
rect 288492 154068 288498 154080
rect 361022 154068 361028 154080
rect 288492 154040 361028 154068
rect 288492 154028 288498 154040
rect 361022 154028 361028 154040
rect 361080 154028 361086 154080
rect 298094 153960 298100 154012
rect 298152 154000 298158 154012
rect 372890 154000 372896 154012
rect 298152 153972 372896 154000
rect 298152 153960 298158 153972
rect 372890 153960 372896 153972
rect 372948 153960 372954 154012
rect 293954 153892 293960 153944
rect 294012 153932 294018 153944
rect 369302 153932 369308 153944
rect 294012 153904 369308 153932
rect 294012 153892 294018 153904
rect 369302 153892 369308 153904
rect 369360 153892 369366 153944
rect 285674 153824 285680 153876
rect 285732 153864 285738 153876
rect 367830 153864 367836 153876
rect 285732 153836 367836 153864
rect 285732 153824 285738 153836
rect 367830 153824 367836 153836
rect 367888 153824 367894 153876
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 199378 150396 199384 150408
rect 3568 150368 199384 150396
rect 3568 150356 3574 150368
rect 199378 150356 199384 150368
rect 199436 150356 199442 150408
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 203518 137952 203524 137964
rect 3568 137924 203524 137952
rect 3568 137912 3574 137924
rect 203518 137912 203524 137924
rect 203576 137912 203582 137964
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 197998 97968 198004 97980
rect 3476 97940 198004 97968
rect 3476 97928 3482 97940
rect 197998 97928 198004 97940
rect 198056 97928 198062 97980
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 206278 85524 206284 85536
rect 3200 85496 206284 85524
rect 3200 85484 3206 85496
rect 206278 85484 206284 85496
rect 206336 85484 206342 85536
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 207658 71720 207664 71732
rect 3476 71692 207664 71720
rect 3476 71680 3482 71692
rect 207658 71680 207664 71692
rect 207716 71680 207722 71732
rect 378778 60664 378784 60716
rect 378836 60704 378842 60716
rect 580166 60704 580172 60716
rect 378836 60676 580172 60704
rect 378836 60664 378842 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 25498 59344 25504 59356
rect 3108 59316 25504 59344
rect 3108 59304 3114 59316
rect 25498 59304 25504 59316
rect 25556 59304 25562 59356
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 82078 45540 82084 45552
rect 3476 45512 82084 45540
rect 3476 45500 3482 45512
rect 82078 45500 82084 45512
rect 82136 45500 82142 45552
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 88978 33096 88984 33108
rect 3568 33068 88984 33096
rect 3568 33056 3574 33068
rect 88978 33056 88984 33068
rect 89036 33056 89042 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 192570 20652 192576 20664
rect 3476 20624 192576 20652
rect 3476 20612 3482 20624
rect 192570 20612 192576 20624
rect 192628 20612 192634 20664
rect 160094 11704 160100 11756
rect 160152 11744 160158 11756
rect 161290 11744 161296 11756
rect 160152 11716 161296 11744
rect 160152 11704 160158 11716
rect 161290 11704 161296 11716
rect 161348 11704 161354 11756
rect 176654 11704 176660 11756
rect 176712 11744 176718 11756
rect 177850 11744 177856 11756
rect 176712 11716 177856 11744
rect 176712 11704 176718 11716
rect 177850 11704 177856 11716
rect 177908 11704 177914 11756
rect 184934 11704 184940 11756
rect 184992 11744 184998 11756
rect 186130 11744 186136 11756
rect 184992 11716 186136 11744
rect 184992 11704 184998 11716
rect 186130 11704 186136 11716
rect 186188 11704 186194 11756
rect 201494 11704 201500 11756
rect 201552 11744 201558 11756
rect 202690 11744 202696 11756
rect 201552 11716 202696 11744
rect 201552 11704 201558 11716
rect 202690 11704 202696 11716
rect 202748 11704 202754 11756
rect 234614 11704 234620 11756
rect 234672 11744 234678 11756
rect 235810 11744 235816 11756
rect 234672 11716 235816 11744
rect 234672 11704 234678 11716
rect 235810 11704 235816 11716
rect 235868 11704 235874 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 319714 9392 319720 9444
rect 319772 9432 319778 9444
rect 365806 9432 365812 9444
rect 319772 9404 365812 9432
rect 319772 9392 319778 9404
rect 365806 9392 365812 9404
rect 365864 9392 365870 9444
rect 316218 9324 316224 9376
rect 316276 9364 316282 9376
rect 364702 9364 364708 9376
rect 316276 9336 364708 9364
rect 316276 9324 316282 9336
rect 364702 9324 364708 9336
rect 364760 9324 364766 9376
rect 322106 9256 322112 9308
rect 322164 9296 322170 9308
rect 372706 9296 372712 9308
rect 322164 9268 372712 9296
rect 322164 9256 322170 9268
rect 372706 9256 372712 9268
rect 372764 9256 372770 9308
rect 303154 9188 303160 9240
rect 303212 9228 303218 9240
rect 358262 9228 358268 9240
rect 303212 9200 358268 9228
rect 303212 9188 303218 9200
rect 358262 9188 358268 9200
rect 358320 9188 358326 9240
rect 306742 9120 306748 9172
rect 306800 9160 306806 9172
rect 368474 9160 368480 9172
rect 306800 9132 368480 9160
rect 306800 9120 306806 9132
rect 368474 9120 368480 9132
rect 368532 9120 368538 9172
rect 309042 9052 309048 9104
rect 309100 9092 309106 9104
rect 369946 9092 369952 9104
rect 309100 9064 369952 9092
rect 309100 9052 309106 9064
rect 369946 9052 369952 9064
rect 370004 9052 370010 9104
rect 305546 8984 305552 9036
rect 305604 9024 305610 9036
rect 367186 9024 367192 9036
rect 305604 8996 367192 9024
rect 305604 8984 305610 8996
rect 367186 8984 367192 8996
rect 367244 8984 367250 9036
rect 304350 8916 304356 8968
rect 304408 8956 304414 8968
rect 366082 8956 366088 8968
rect 304408 8928 366088 8956
rect 304408 8916 304414 8928
rect 366082 8916 366088 8928
rect 366140 8916 366146 8968
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 200758 6848 200764 6860
rect 3476 6820 200764 6848
rect 3476 6808 3482 6820
rect 200758 6808 200764 6820
rect 200816 6808 200822 6860
rect 337470 6808 337476 6860
rect 337528 6848 337534 6860
rect 363138 6848 363144 6860
rect 337528 6820 363144 6848
rect 337528 6808 337534 6820
rect 363138 6808 363144 6820
rect 363196 6808 363202 6860
rect 333882 6740 333888 6792
rect 333940 6780 333946 6792
rect 363230 6780 363236 6792
rect 333940 6752 363236 6780
rect 333940 6740 333946 6752
rect 363230 6740 363236 6752
rect 363288 6740 363294 6792
rect 577498 6740 577504 6792
rect 577556 6780 577562 6792
rect 580258 6780 580264 6792
rect 577556 6752 580264 6780
rect 577556 6740 577562 6752
rect 580258 6740 580264 6752
rect 580316 6740 580322 6792
rect 330386 6672 330392 6724
rect 330444 6712 330450 6724
rect 363322 6712 363328 6724
rect 330444 6684 363328 6712
rect 330444 6672 330450 6684
rect 363322 6672 363328 6684
rect 363380 6672 363386 6724
rect 318518 6604 318524 6656
rect 318576 6644 318582 6656
rect 364334 6644 364340 6656
rect 318576 6616 364340 6644
rect 318576 6604 318582 6616
rect 364334 6604 364340 6616
rect 364392 6604 364398 6656
rect 313826 6536 313832 6588
rect 313884 6576 313890 6588
rect 360286 6576 360292 6588
rect 313884 6548 360292 6576
rect 313884 6536 313890 6548
rect 360286 6536 360292 6548
rect 360344 6536 360350 6588
rect 317322 6468 317328 6520
rect 317380 6508 317386 6520
rect 363414 6508 363420 6520
rect 317380 6480 363420 6508
rect 317380 6468 317386 6480
rect 363414 6468 363420 6480
rect 363472 6468 363478 6520
rect 315022 6400 315028 6452
rect 315080 6440 315086 6452
rect 362034 6440 362040 6452
rect 315080 6412 362040 6440
rect 315080 6400 315086 6412
rect 362034 6400 362040 6412
rect 362092 6400 362098 6452
rect 312630 6332 312636 6384
rect 312688 6372 312694 6384
rect 360194 6372 360200 6384
rect 312688 6344 360200 6372
rect 312688 6332 312694 6344
rect 360194 6332 360200 6344
rect 360252 6332 360258 6384
rect 311434 6264 311440 6316
rect 311492 6304 311498 6316
rect 358814 6304 358820 6316
rect 311492 6276 358820 6304
rect 311492 6264 311498 6276
rect 358814 6264 358820 6276
rect 358872 6264 358878 6316
rect 307938 6196 307944 6248
rect 307996 6236 308002 6248
rect 369854 6236 369860 6248
rect 307996 6208 369860 6236
rect 307996 6196 308002 6208
rect 369854 6196 369860 6208
rect 369912 6196 369918 6248
rect 310238 6128 310244 6180
rect 310296 6168 310302 6180
rect 371326 6168 371332 6180
rect 310296 6140 371332 6168
rect 310296 6128 310302 6140
rect 371326 6128 371332 6140
rect 371384 6128 371390 6180
rect 340966 6060 340972 6112
rect 341024 6100 341030 6112
rect 365898 6100 365904 6112
rect 341024 6072 365904 6100
rect 341024 6060 341030 6072
rect 365898 6060 365904 6072
rect 365956 6060 365962 6112
rect 344554 5992 344560 6044
rect 344612 6032 344618 6044
rect 365990 6032 365996 6044
rect 344612 6004 365996 6032
rect 344612 5992 344618 6004
rect 365990 5992 365996 6004
rect 366048 5992 366054 6044
rect 350442 5924 350448 5976
rect 350500 5964 350506 5976
rect 364610 5964 364616 5976
rect 350500 5936 364616 5964
rect 350500 5924 350506 5936
rect 364610 5924 364616 5936
rect 364668 5924 364674 5976
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 8938 4128 8944 4140
rect 6512 4100 8944 4128
rect 6512 4088 6518 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 44266 4088 44272 4140
rect 44324 4128 44330 4140
rect 46198 4128 46204 4140
rect 44324 4100 46204 4128
rect 44324 4088 44330 4100
rect 46198 4088 46204 4100
rect 46256 4088 46262 4140
rect 180242 4088 180248 4140
rect 180300 4128 180306 4140
rect 181438 4128 181444 4140
rect 180300 4100 181444 4128
rect 180300 4088 180306 4100
rect 181438 4088 181444 4100
rect 181496 4088 181502 4140
rect 216398 4088 216404 4140
rect 216456 4128 216462 4140
rect 240502 4128 240508 4140
rect 216456 4100 240508 4128
rect 216456 4088 216462 4100
rect 240502 4088 240508 4100
rect 240560 4088 240566 4140
rect 336274 4088 336280 4140
rect 336332 4128 336338 4140
rect 364426 4128 364432 4140
rect 336332 4100 364432 4128
rect 336332 4088 336338 4100
rect 364426 4088 364432 4100
rect 364484 4088 364490 4140
rect 428550 4088 428556 4140
rect 428608 4128 428614 4140
rect 434438 4128 434444 4140
rect 428608 4100 434444 4128
rect 428608 4088 428614 4100
rect 434438 4088 434444 4100
rect 434496 4088 434502 4140
rect 460198 4088 460204 4140
rect 460256 4128 460262 4140
rect 462774 4128 462780 4140
rect 460256 4100 462780 4128
rect 460256 4088 460262 4100
rect 462774 4088 462780 4100
rect 462832 4088 462838 4140
rect 468478 4088 468484 4140
rect 468536 4128 468542 4140
rect 471054 4128 471060 4140
rect 468536 4100 471060 4128
rect 468536 4088 468542 4100
rect 471054 4088 471060 4100
rect 471112 4088 471118 4140
rect 478230 4088 478236 4140
rect 478288 4128 478294 4140
rect 482830 4128 482836 4140
rect 478288 4100 482836 4128
rect 478288 4088 478294 4100
rect 482830 4088 482836 4100
rect 482888 4088 482894 4140
rect 536190 4088 536196 4140
rect 536248 4128 536254 4140
rect 538398 4128 538404 4140
rect 536248 4100 538404 4128
rect 536248 4088 536254 4100
rect 538398 4088 538404 4100
rect 538456 4088 538462 4140
rect 51350 4020 51356 4072
rect 51408 4060 51414 4072
rect 57238 4060 57244 4072
rect 51408 4032 57244 4060
rect 51408 4020 51414 4032
rect 57238 4020 57244 4032
rect 57296 4020 57302 4072
rect 212350 4020 212356 4072
rect 212408 4060 212414 4072
rect 245194 4060 245200 4072
rect 212408 4032 245200 4060
rect 212408 4020 212414 4032
rect 245194 4020 245200 4032
rect 245252 4020 245258 4072
rect 332686 4020 332692 4072
rect 332744 4060 332750 4072
rect 363046 4060 363052 4072
rect 332744 4032 363052 4060
rect 332744 4020 332750 4032
rect 363046 4020 363052 4032
rect 363104 4020 363110 4072
rect 213730 3952 213736 4004
rect 213788 3992 213794 4004
rect 258258 3992 258264 4004
rect 213788 3964 258264 3992
rect 213788 3952 213794 3964
rect 258258 3952 258264 3964
rect 258316 3952 258322 4004
rect 329190 3952 329196 4004
rect 329248 3992 329254 4004
rect 362954 3992 362960 4004
rect 329248 3964 362960 3992
rect 329248 3952 329254 3964
rect 362954 3952 362960 3964
rect 363012 3952 363018 4004
rect 213822 3884 213828 3936
rect 213880 3924 213886 3936
rect 260650 3924 260656 3936
rect 213880 3896 260656 3924
rect 213880 3884 213886 3896
rect 260650 3884 260656 3896
rect 260708 3884 260714 3936
rect 301958 3884 301964 3936
rect 302016 3924 302022 3936
rect 352558 3924 352564 3936
rect 302016 3896 352564 3924
rect 302016 3884 302022 3896
rect 352558 3884 352564 3896
rect 352616 3884 352622 3936
rect 4062 3816 4068 3868
rect 4120 3856 4126 3868
rect 7558 3856 7564 3868
rect 4120 3828 7564 3856
rect 4120 3816 4126 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 215018 3816 215024 3868
rect 215076 3856 215082 3868
rect 262950 3856 262956 3868
rect 215076 3828 262956 3856
rect 215076 3816 215082 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 291378 3816 291384 3868
rect 291436 3856 291442 3868
rect 345750 3856 345756 3868
rect 291436 3828 345756 3856
rect 291436 3816 291442 3828
rect 345750 3816 345756 3828
rect 345808 3816 345814 3868
rect 354030 3816 354036 3868
rect 354088 3856 354094 3868
rect 363782 3856 363788 3868
rect 354088 3828 363788 3856
rect 354088 3816 354094 3828
rect 363782 3816 363788 3828
rect 363840 3816 363846 3868
rect 440878 3816 440884 3868
rect 440936 3856 440942 3868
rect 443822 3856 443828 3868
rect 440936 3828 443828 3856
rect 440936 3816 440942 3828
rect 443822 3816 443828 3828
rect 443880 3816 443886 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 519538 3856 519544 3868
rect 516836 3828 519544 3856
rect 516836 3816 516842 3828
rect 519538 3816 519544 3828
rect 519596 3816 519602 3868
rect 566458 3816 566464 3868
rect 566516 3856 566522 3868
rect 569126 3856 569132 3868
rect 566516 3828 569132 3856
rect 566516 3816 566522 3828
rect 569126 3816 569132 3828
rect 569184 3816 569190 3868
rect 211062 3748 211068 3800
rect 211120 3788 211126 3800
rect 268838 3788 268844 3800
rect 211120 3760 268844 3788
rect 211120 3748 211126 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 292574 3748 292580 3800
rect 292632 3788 292638 3800
rect 348418 3788 348424 3800
rect 292632 3760 348424 3788
rect 292632 3748 292638 3760
rect 348418 3748 348424 3760
rect 348476 3748 348482 3800
rect 349246 3748 349252 3800
rect 349304 3788 349310 3800
rect 361850 3788 361856 3800
rect 349304 3760 361856 3788
rect 349304 3748 349310 3760
rect 361850 3748 361856 3760
rect 361908 3748 361914 3800
rect 30098 3680 30104 3732
rect 30156 3720 30162 3732
rect 39390 3720 39396 3732
rect 30156 3692 39396 3720
rect 30156 3680 30162 3692
rect 39390 3680 39396 3692
rect 39448 3680 39454 3732
rect 69106 3680 69112 3732
rect 69164 3720 69170 3732
rect 71038 3720 71044 3732
rect 69164 3692 71044 3720
rect 69164 3680 69170 3692
rect 71038 3680 71044 3692
rect 71096 3680 71102 3732
rect 135254 3680 135260 3732
rect 135312 3720 135318 3732
rect 136450 3720 136456 3732
rect 135312 3692 136456 3720
rect 135312 3680 135318 3692
rect 136450 3680 136456 3692
rect 136508 3680 136514 3732
rect 212258 3680 212264 3732
rect 212316 3720 212322 3732
rect 272426 3720 272432 3732
rect 212316 3692 272432 3720
rect 212316 3680 212322 3692
rect 272426 3680 272432 3692
rect 272484 3680 272490 3732
rect 299566 3680 299572 3732
rect 299624 3720 299630 3732
rect 300762 3720 300768 3732
rect 299624 3692 300768 3720
rect 299624 3680 299630 3692
rect 300762 3680 300768 3692
rect 300820 3680 300826 3732
rect 301774 3680 301780 3732
rect 301832 3720 301838 3732
rect 353938 3720 353944 3732
rect 301832 3692 353944 3720
rect 301832 3680 301838 3692
rect 353938 3680 353944 3692
rect 353996 3680 354002 3732
rect 445018 3680 445024 3732
rect 445076 3720 445082 3732
rect 458082 3720 458088 3732
rect 445076 3692 458088 3720
rect 445076 3680 445082 3692
rect 458082 3680 458088 3692
rect 458140 3680 458146 3732
rect 489178 3680 489184 3732
rect 489236 3720 489242 3732
rect 491110 3720 491116 3732
rect 489236 3692 491116 3720
rect 489236 3680 489242 3692
rect 491110 3680 491116 3692
rect 491168 3680 491174 3732
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 32398 3652 32404 3664
rect 1728 3624 32404 3652
rect 1728 3612 1734 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 37182 3612 37188 3664
rect 37240 3652 37246 3664
rect 43438 3652 43444 3664
rect 37240 3624 43444 3652
rect 37240 3612 37246 3624
rect 43438 3612 43444 3624
rect 43496 3612 43502 3664
rect 46658 3612 46664 3664
rect 46716 3652 46722 3664
rect 170490 3652 170496 3664
rect 46716 3624 170496 3652
rect 46716 3612 46722 3624
rect 170490 3612 170496 3624
rect 170548 3612 170554 3664
rect 187326 3612 187332 3664
rect 187384 3652 187390 3664
rect 196618 3652 196624 3664
rect 187384 3624 196624 3652
rect 187384 3612 187390 3624
rect 196618 3612 196624 3624
rect 196676 3612 196682 3664
rect 215938 3612 215944 3664
rect 215996 3652 216002 3664
rect 276014 3652 276020 3664
rect 215996 3624 276020 3652
rect 215996 3612 216002 3624
rect 276014 3612 276020 3624
rect 276072 3612 276078 3664
rect 285398 3612 285404 3664
rect 285456 3652 285462 3664
rect 345658 3652 345664 3664
rect 285456 3624 345664 3652
rect 285456 3612 285462 3624
rect 345658 3612 345664 3624
rect 345716 3612 345722 3664
rect 346946 3612 346952 3664
rect 347004 3652 347010 3664
rect 363874 3652 363880 3664
rect 347004 3624 363880 3652
rect 347004 3612 347010 3624
rect 363874 3612 363880 3624
rect 363932 3612 363938 3664
rect 427078 3612 427084 3664
rect 427136 3652 427142 3664
rect 440326 3652 440332 3664
rect 427136 3624 440332 3652
rect 427136 3612 427142 3624
rect 440326 3612 440332 3624
rect 440384 3612 440390 3664
rect 476758 3612 476764 3664
rect 476816 3652 476822 3664
rect 476816 3624 480254 3652
rect 476816 3612 476822 3624
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 21358 3584 21364 3596
rect 20680 3556 21364 3584
rect 20680 3544 20686 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 171778 3584 171784 3596
rect 25372 3556 171784 3584
rect 25372 3544 25378 3556
rect 171778 3544 171784 3556
rect 171836 3544 171842 3596
rect 183738 3544 183744 3596
rect 183796 3584 183802 3596
rect 188338 3584 188344 3596
rect 183796 3556 188344 3584
rect 183796 3544 183802 3556
rect 188338 3544 188344 3556
rect 188396 3544 188402 3596
rect 195606 3544 195612 3596
rect 195664 3584 195670 3596
rect 203610 3584 203616 3596
rect 195664 3556 203616 3584
rect 195664 3544 195670 3556
rect 203610 3544 203616 3556
rect 203668 3544 203674 3596
rect 216582 3544 216588 3596
rect 216640 3584 216646 3596
rect 284294 3584 284300 3596
rect 216640 3556 284300 3584
rect 216640 3544 216646 3556
rect 284294 3544 284300 3556
rect 284352 3544 284358 3596
rect 287790 3544 287796 3596
rect 287848 3584 287854 3596
rect 354122 3584 354128 3596
rect 287848 3556 354128 3584
rect 287848 3544 287854 3556
rect 354122 3544 354128 3556
rect 354180 3544 354186 3596
rect 355226 3544 355232 3596
rect 355284 3584 355290 3596
rect 365714 3584 365720 3596
rect 355284 3556 365720 3584
rect 355284 3544 355290 3556
rect 365714 3544 365720 3556
rect 365772 3544 365778 3596
rect 377398 3544 377404 3596
rect 377456 3584 377462 3596
rect 411898 3584 411904 3596
rect 377456 3556 411904 3584
rect 377456 3544 377462 3556
rect 411898 3544 411904 3556
rect 411956 3544 411962 3596
rect 421558 3544 421564 3596
rect 421616 3584 421622 3596
rect 427262 3584 427268 3596
rect 421616 3556 427268 3584
rect 421616 3544 421622 3556
rect 427262 3544 427268 3556
rect 427320 3544 427326 3596
rect 442258 3544 442264 3596
rect 442316 3584 442322 3596
rect 445018 3584 445024 3596
rect 442316 3556 445024 3584
rect 442316 3544 442322 3556
rect 445018 3544 445024 3556
rect 445076 3544 445082 3596
rect 458818 3544 458824 3596
rect 458876 3584 458882 3596
rect 465166 3584 465172 3596
rect 458876 3556 465172 3584
rect 458876 3544 458882 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 469858 3584 469864 3596
rect 467156 3556 469864 3584
rect 467156 3544 467162 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 470566 3556 475240 3584
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 13078 3516 13084 3528
rect 12400 3488 13084 3516
rect 12400 3476 12406 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 170398 3516 170404 3528
rect 15988 3488 170404 3516
rect 15988 3476 15994 3488
rect 170398 3476 170404 3488
rect 170456 3476 170462 3528
rect 219342 3476 219348 3528
rect 219400 3516 219406 3528
rect 280706 3516 280712 3528
rect 219400 3488 280712 3516
rect 219400 3476 219406 3488
rect 280706 3476 280712 3488
rect 280764 3476 280770 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 357434 3516 357440 3528
rect 281960 3488 357440 3516
rect 281960 3476 281966 3488
rect 357434 3476 357440 3488
rect 357492 3476 357498 3528
rect 374086 3476 374092 3528
rect 374144 3516 374150 3528
rect 375282 3516 375288 3528
rect 374144 3488 375288 3516
rect 374144 3476 374150 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 381538 3476 381544 3528
rect 381596 3516 381602 3528
rect 381596 3488 423628 3516
rect 381596 3476 381602 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 171134 3448 171140 3460
rect 624 3420 171140 3448
rect 624 3408 630 3420
rect 171134 3408 171140 3420
rect 171192 3408 171198 3460
rect 190822 3408 190828 3460
rect 190880 3448 190886 3460
rect 199470 3448 199476 3460
rect 190880 3420 199476 3448
rect 190880 3408 190886 3420
rect 199470 3408 199476 3420
rect 199528 3408 199534 3460
rect 215110 3408 215116 3460
rect 215168 3448 215174 3460
rect 277118 3448 277124 3460
rect 215168 3420 277124 3448
rect 215168 3408 215174 3420
rect 277118 3408 277124 3420
rect 277176 3408 277182 3460
rect 283098 3408 283104 3460
rect 283156 3448 283162 3460
rect 367094 3448 367100 3460
rect 283156 3420 367100 3448
rect 283156 3408 283162 3420
rect 367094 3408 367100 3420
rect 367152 3408 367158 3460
rect 373258 3408 373264 3460
rect 373316 3448 373322 3460
rect 384758 3448 384764 3460
rect 373316 3420 384764 3448
rect 373316 3408 373322 3420
rect 384758 3408 384764 3420
rect 384816 3408 384822 3460
rect 387058 3408 387064 3460
rect 387116 3448 387122 3460
rect 388254 3448 388260 3460
rect 387116 3420 388260 3448
rect 387116 3408 387122 3420
rect 388254 3408 388260 3420
rect 388312 3408 388318 3460
rect 390554 3408 390560 3460
rect 390612 3448 390618 3460
rect 391842 3448 391848 3460
rect 390612 3420 391848 3448
rect 390612 3408 390618 3420
rect 391842 3408 391848 3420
rect 391900 3408 391906 3460
rect 393286 3420 412634 3448
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 35158 3380 35164 3392
rect 33652 3352 35164 3380
rect 33652 3340 33658 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 57330 3380 57336 3392
rect 56100 3352 57336 3380
rect 56100 3340 56106 3352
rect 57330 3340 57336 3352
rect 57388 3340 57394 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 212442 3340 212448 3392
rect 212500 3380 212506 3392
rect 227530 3380 227536 3392
rect 212500 3352 227536 3380
rect 212500 3340 212506 3352
rect 227530 3340 227536 3352
rect 227588 3340 227594 3392
rect 297266 3340 297272 3392
rect 297324 3380 297330 3392
rect 301774 3380 301780 3392
rect 297324 3352 301780 3380
rect 297324 3340 297330 3352
rect 301774 3340 301780 3352
rect 301832 3340 301838 3392
rect 338666 3340 338672 3392
rect 338724 3380 338730 3392
rect 361942 3380 361948 3392
rect 338724 3352 361948 3380
rect 338724 3340 338730 3352
rect 361942 3340 361948 3352
rect 362000 3340 362006 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 388438 3340 388444 3392
rect 388496 3380 388502 3392
rect 393286 3380 393314 3420
rect 388496 3352 393314 3380
rect 388496 3340 388502 3352
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 57238 3272 57244 3324
rect 57296 3312 57302 3324
rect 58618 3312 58624 3324
rect 57296 3284 58624 3312
rect 57296 3272 57302 3284
rect 58618 3272 58624 3284
rect 58676 3272 58682 3324
rect 208578 3272 208584 3324
rect 208636 3312 208642 3324
rect 211798 3312 211804 3324
rect 208636 3284 211804 3312
rect 208636 3272 208642 3284
rect 211798 3272 211804 3284
rect 211856 3272 211862 3324
rect 215202 3272 215208 3324
rect 215260 3312 215266 3324
rect 222746 3312 222752 3324
rect 215260 3284 222752 3312
rect 215260 3272 215266 3284
rect 222746 3272 222752 3284
rect 222804 3272 222810 3324
rect 343358 3272 343364 3324
rect 343416 3312 343422 3324
rect 364518 3312 364524 3324
rect 343416 3284 364524 3312
rect 343416 3272 343422 3284
rect 364518 3272 364524 3284
rect 364576 3272 364582 3324
rect 412606 3312 412634 3420
rect 414658 3408 414664 3460
rect 414716 3448 414722 3460
rect 416682 3448 416688 3460
rect 414716 3420 416688 3448
rect 414716 3408 414722 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 423600 3380 423628 3488
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 431954 3476 431960 3528
rect 432012 3516 432018 3528
rect 433242 3516 433248 3528
rect 432012 3488 433248 3516
rect 432012 3476 432018 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 439498 3476 439504 3528
rect 439556 3516 439562 3528
rect 441522 3516 441528 3528
rect 439556 3488 441528 3516
rect 439556 3476 439562 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 448514 3476 448520 3528
rect 448572 3516 448578 3528
rect 449802 3516 449808 3528
rect 448572 3488 449808 3516
rect 448572 3476 448578 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 454678 3476 454684 3528
rect 454736 3516 454742 3528
rect 456886 3516 456892 3528
rect 454736 3488 456892 3516
rect 454736 3476 454742 3488
rect 456886 3476 456892 3488
rect 456944 3476 456950 3528
rect 462958 3476 462964 3528
rect 463016 3516 463022 3528
rect 470566 3516 470594 3556
rect 463016 3488 470594 3516
rect 463016 3476 463022 3488
rect 471238 3476 471244 3528
rect 471296 3516 471302 3528
rect 473446 3516 473452 3528
rect 471296 3488 473452 3516
rect 471296 3476 471302 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 475212 3516 475240 3556
rect 475378 3544 475384 3596
rect 475436 3584 475442 3596
rect 476942 3584 476948 3596
rect 475436 3556 476948 3584
rect 475436 3544 475442 3556
rect 476942 3544 476948 3556
rect 477000 3544 477006 3596
rect 480226 3584 480254 3624
rect 484026 3584 484032 3596
rect 480226 3556 484032 3584
rect 484026 3544 484032 3556
rect 484084 3544 484090 3596
rect 500218 3544 500224 3596
rect 500276 3584 500282 3596
rect 501782 3584 501788 3596
rect 500276 3556 501788 3584
rect 500276 3544 500282 3556
rect 501782 3544 501788 3556
rect 501840 3544 501846 3596
rect 511258 3544 511264 3596
rect 511316 3584 511322 3596
rect 513558 3584 513564 3596
rect 511316 3556 513564 3584
rect 511316 3544 511322 3556
rect 513558 3544 513564 3556
rect 513616 3544 513622 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 527726 3584 527732 3596
rect 525116 3556 527732 3584
rect 525116 3544 525122 3556
rect 527726 3544 527732 3556
rect 527784 3544 527790 3596
rect 533706 3584 533712 3596
rect 528526 3556 533712 3584
rect 479334 3516 479340 3528
rect 475212 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 496078 3476 496084 3528
rect 496136 3516 496142 3528
rect 497090 3516 497096 3528
rect 496136 3488 497096 3516
rect 496136 3476 496142 3488
rect 497090 3476 497096 3488
rect 497148 3476 497154 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 520918 3476 520924 3528
rect 520976 3516 520982 3528
rect 523034 3516 523040 3528
rect 520976 3488 523040 3516
rect 520976 3476 520982 3488
rect 523034 3476 523040 3488
rect 523092 3476 523098 3528
rect 527818 3476 527824 3528
rect 527876 3516 527882 3528
rect 528526 3516 528554 3556
rect 533706 3544 533712 3556
rect 533764 3544 533770 3596
rect 549898 3544 549904 3596
rect 549956 3584 549962 3596
rect 551462 3584 551468 3596
rect 549956 3556 551468 3584
rect 549956 3544 549962 3556
rect 551462 3544 551468 3556
rect 551520 3544 551526 3596
rect 527876 3488 528554 3516
rect 527876 3476 527882 3488
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 545758 3476 545764 3528
rect 545816 3516 545822 3528
rect 546678 3516 546684 3528
rect 545816 3488 546684 3516
rect 545816 3476 545822 3488
rect 546678 3476 546684 3488
rect 546736 3476 546742 3528
rect 570598 3476 570604 3528
rect 570656 3516 570662 3528
rect 572714 3516 572720 3528
rect 570656 3488 572720 3516
rect 570656 3476 570662 3488
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 580994 3448 581000 3460
rect 431926 3420 581000 3448
rect 429654 3380 429660 3392
rect 423600 3352 429660 3380
rect 429654 3340 429660 3352
rect 429712 3340 429718 3392
rect 431926 3312 431954 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 493318 3340 493324 3392
rect 493376 3380 493382 3392
rect 499390 3380 499396 3392
rect 493376 3352 499396 3380
rect 493376 3340 493382 3352
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 542998 3340 543004 3392
rect 543056 3380 543062 3392
rect 549070 3380 549076 3392
rect 543056 3352 549076 3380
rect 543056 3340 543062 3352
rect 549070 3340 549076 3352
rect 549128 3340 549134 3392
rect 412606 3284 431954 3312
rect 446398 3272 446404 3324
rect 446456 3312 446462 3324
rect 452102 3312 452108 3324
rect 446456 3284 452108 3312
rect 446456 3272 446462 3284
rect 452102 3272 452108 3284
rect 452160 3272 452166 3324
rect 509878 3272 509884 3324
rect 509936 3312 509942 3324
rect 514754 3312 514760 3324
rect 509936 3284 514760 3312
rect 509936 3272 509942 3284
rect 514754 3272 514760 3284
rect 514812 3272 514818 3324
rect 216490 3204 216496 3256
rect 216548 3244 216554 3256
rect 226334 3244 226340 3256
rect 216548 3216 226340 3244
rect 216548 3204 216554 3216
rect 226334 3204 226340 3216
rect 226392 3204 226398 3256
rect 342162 3204 342168 3256
rect 342220 3244 342226 3256
rect 361666 3244 361672 3256
rect 342220 3216 361672 3244
rect 342220 3204 342226 3216
rect 361666 3204 361672 3216
rect 361724 3204 361730 3256
rect 404998 3204 405004 3256
rect 405056 3244 405062 3256
rect 408402 3244 408408 3256
rect 405056 3216 408408 3244
rect 405056 3204 405062 3216
rect 408402 3204 408408 3216
rect 408460 3204 408466 3256
rect 554038 3204 554044 3256
rect 554096 3244 554102 3256
rect 557350 3244 557356 3256
rect 554096 3216 557356 3244
rect 554096 3204 554102 3216
rect 557350 3204 557356 3216
rect 557408 3204 557414 3256
rect 345750 3136 345756 3188
rect 345808 3176 345814 3188
rect 361758 3176 361764 3188
rect 345808 3148 361764 3176
rect 345808 3136 345814 3148
rect 361758 3136 361764 3148
rect 361816 3136 361822 3188
rect 371878 3136 371884 3188
rect 371936 3176 371942 3188
rect 376478 3176 376484 3188
rect 371936 3148 376484 3176
rect 371936 3136 371942 3148
rect 376478 3136 376484 3148
rect 376536 3136 376542 3188
rect 435358 3136 435364 3188
rect 435416 3176 435422 3188
rect 437934 3176 437940 3188
rect 435416 3148 437940 3176
rect 435416 3136 435422 3148
rect 437934 3136 437940 3148
rect 437992 3136 437998 3188
rect 485038 3136 485044 3188
rect 485096 3176 485102 3188
rect 487614 3176 487620 3188
rect 485096 3148 487620 3176
rect 485096 3136 485102 3148
rect 487614 3136 487620 3148
rect 487672 3136 487678 3188
rect 534718 3136 534724 3188
rect 534776 3176 534782 3188
rect 537202 3176 537208 3188
rect 534776 3148 537208 3176
rect 534776 3136 534782 3148
rect 537202 3136 537208 3148
rect 537260 3136 537266 3188
rect 560938 3136 560944 3188
rect 560996 3176 561002 3188
rect 563238 3176 563244 3188
rect 560996 3148 563244 3176
rect 560996 3136 561002 3148
rect 563238 3136 563244 3148
rect 563296 3136 563302 3188
rect 352834 3068 352840 3120
rect 352892 3108 352898 3120
rect 362494 3108 362500 3120
rect 352892 3080 362500 3108
rect 352892 3068 352898 3080
rect 362494 3068 362500 3080
rect 362552 3068 362558 3120
rect 445110 3068 445116 3120
rect 445168 3108 445174 3120
rect 447410 3108 447416 3120
rect 445168 3080 447416 3108
rect 445168 3068 445174 3080
rect 447410 3068 447416 3080
rect 447468 3068 447474 3120
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 25590 3040 25596 3052
rect 19484 3012 25596 3040
rect 19484 3000 19490 3012
rect 25590 3000 25596 3012
rect 25648 3000 25654 3052
rect 413278 3000 413284 3052
rect 413336 3040 413342 3052
rect 415486 3040 415492 3052
rect 413336 3012 415492 3040
rect 413336 3000 413342 3012
rect 415486 3000 415492 3012
rect 415544 3000 415550 3052
rect 417510 3000 417516 3052
rect 417568 3040 417574 3052
rect 420178 3040 420184 3052
rect 417568 3012 420184 3040
rect 417568 3000 417574 3012
rect 420178 3000 420184 3012
rect 420236 3000 420242 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 486510 3000 486516 3052
rect 486568 3040 486574 3052
rect 488810 3040 488816 3052
rect 486568 3012 488816 3040
rect 486568 3000 486574 3012
rect 488810 3000 488816 3012
rect 488868 3000 488874 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 522298 3000 522304 3052
rect 522356 3040 522362 3052
rect 524230 3040 524236 3052
rect 522356 3012 524236 3040
rect 522356 3000 522362 3012
rect 524230 3000 524236 3012
rect 524288 3000 524294 3052
rect 538858 3000 538864 3052
rect 538916 3040 538922 3052
rect 540790 3040 540796 3052
rect 538916 3012 540796 3040
rect 538916 3000 538922 3012
rect 540790 3000 540796 3012
rect 540848 3000 540854 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565630 3040 565636 3052
rect 563756 3012 565636 3040
rect 563756 3000 563762 3012
rect 565630 3000 565636 3012
rect 565688 3000 565694 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 396718 2932 396724 2984
rect 396776 2972 396782 2984
rect 402514 2972 402520 2984
rect 396776 2944 402520 2972
rect 396776 2932 396782 2944
rect 402514 2932 402520 2944
rect 402572 2932 402578 2984
rect 540238 2932 540244 2984
rect 540296 2972 540302 2984
rect 541986 2972 541992 2984
rect 540296 2944 541992 2972
rect 540296 2932 540302 2944
rect 541986 2932 541992 2944
rect 542044 2932 542050 2984
rect 552750 2932 552756 2984
rect 552808 2972 552814 2984
rect 554958 2972 554964 2984
rect 552808 2944 554964 2972
rect 552808 2932 552814 2944
rect 554958 2932 554964 2944
rect 555016 2932 555022 2984
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 219348 700408 219400 700460
rect 267648 700408 267700 700460
rect 217968 700340 218020 700392
rect 283840 700340 283892 700392
rect 348792 700340 348844 700392
rect 358820 700340 358872 700392
rect 8116 700272 8168 700324
rect 98644 700272 98696 700324
rect 217876 700272 217928 700324
rect 300124 700272 300176 700324
rect 332508 700272 332560 700324
rect 357440 700272 357492 700324
rect 359464 700272 359516 700324
rect 429844 700272 429896 700324
rect 442264 700272 442316 700324
rect 559656 700272 559708 700324
rect 105452 699728 105504 699780
rect 108304 699728 108356 699780
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 137836 699660 137888 699712
rect 140044 699660 140096 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 391204 696940 391256 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 21364 683136 21416 683188
rect 381544 683136 381596 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 215944 670692 215996 670744
rect 377404 670692 377456 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 28264 656888 28316 656940
rect 373264 643084 373316 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 3148 618264 3200 618316
rect 214564 618264 214616 618316
rect 363604 616836 363656 616888
rect 580172 616836 580224 616888
rect 3424 606024 3476 606076
rect 7564 606024 7616 606076
rect 374644 590656 374696 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 57244 579640 57296 579692
rect 378784 576852 378836 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 211804 565836 211856 565888
rect 217784 565088 217836 565140
rect 234620 565088 234672 565140
rect 367744 563048 367796 563100
rect 580172 563048 580224 563100
rect 3424 553664 3476 553716
rect 8944 553664 8996 553716
rect 369124 536800 369176 536852
rect 579896 536800 579948 536852
rect 3424 527144 3476 527196
rect 35164 527144 35216 527196
rect 371884 524424 371936 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 210424 514768 210476 514820
rect 358084 510620 358136 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 13084 500964 13136 501016
rect 360844 484372 360896 484424
rect 580172 484372 580224 484424
rect 217876 478592 217928 478644
rect 269948 478592 270000 478644
rect 217968 478524 218020 478576
rect 271236 478524 271288 478576
rect 268660 478456 268712 478508
rect 357440 478456 357492 478508
rect 269304 478388 269356 478440
rect 358820 478388 358872 478440
rect 217416 478320 217468 478372
rect 308588 478320 308640 478372
rect 218980 478252 219032 478304
rect 314476 478252 314528 478304
rect 256884 478184 256936 478236
rect 374644 478184 374696 478236
rect 7564 478116 7616 478168
rect 282368 478116 282420 478168
rect 241428 476824 241480 476876
rect 238484 476756 238536 476808
rect 237288 476688 237340 476740
rect 239404 476688 239456 476740
rect 316408 476756 316460 476808
rect 311256 476688 311308 476740
rect 242808 476620 242860 476672
rect 319076 476620 319128 476672
rect 271788 476552 271840 476604
rect 330208 476552 330260 476604
rect 266268 476484 266320 476536
rect 326896 476484 326948 476536
rect 256608 476416 256660 476468
rect 318432 476416 318484 476468
rect 318708 476416 318760 476468
rect 336004 476416 336056 476468
rect 262128 476348 262180 476400
rect 323032 476348 323084 476400
rect 326988 476348 327040 476400
rect 338764 476348 338816 476400
rect 309048 476280 309100 476332
rect 329104 476280 329156 476332
rect 311808 476212 311860 476264
rect 331864 476212 331916 476264
rect 315948 476144 316000 476196
rect 334624 476144 334676 476196
rect 240048 476076 240100 476128
rect 313832 476076 313884 476128
rect 314568 476076 314620 476128
rect 333244 476076 333296 476128
rect 321468 475532 321520 475584
rect 355324 475532 355376 475584
rect 274548 475464 274600 475516
rect 331496 475464 331548 475516
rect 219164 475396 219216 475448
rect 321652 475396 321704 475448
rect 255596 475328 255648 475380
rect 371884 475328 371936 475380
rect 3424 474716 3476 474768
rect 287612 474716 287664 474768
rect 264796 474240 264848 474292
rect 297364 474240 297416 474292
rect 274456 474172 274508 474224
rect 353116 474172 353168 474224
rect 219072 474104 219124 474156
rect 317144 474104 317196 474156
rect 252928 474036 252980 474088
rect 360844 474036 360896 474088
rect 153200 473968 153252 474020
rect 275192 473968 275244 474020
rect 253756 472812 253808 472864
rect 329564 472812 329616 472864
rect 217508 472744 217560 472796
rect 323676 472744 323728 472796
rect 254860 472676 254912 472728
rect 369124 472676 369176 472728
rect 8944 472608 8996 472660
rect 284392 472608 284444 472660
rect 302148 472608 302200 472660
rect 345940 472608 345992 472660
rect 259276 471384 259328 471436
rect 294604 471384 294656 471436
rect 217600 471316 217652 471368
rect 327540 471316 327592 471368
rect 13084 471248 13136 471300
rect 286324 471248 286376 471300
rect 286508 471248 286560 471300
rect 338028 471248 338080 471300
rect 253572 470568 253624 470620
rect 580172 470568 580224 470620
rect 248236 470024 248288 470076
rect 310520 470024 310572 470076
rect 257988 469956 258040 470008
rect 333428 469956 333480 470008
rect 257528 469888 257580 469940
rect 378784 469888 378836 469940
rect 35164 469820 35216 469872
rect 285680 469820 285732 469872
rect 293868 469820 293920 469872
rect 341984 469820 342036 469872
rect 253848 468732 253900 468784
rect 301504 468732 301556 468784
rect 280068 468664 280120 468716
rect 356704 468664 356756 468716
rect 219256 468596 219308 468648
rect 319720 468596 319772 468648
rect 264704 468528 264756 468580
rect 462320 468528 462372 468580
rect 57244 468460 57296 468512
rect 283748 468460 283800 468512
rect 248328 467304 248380 467356
rect 320364 467304 320416 467356
rect 217692 467236 217744 467288
rect 325608 467236 325660 467288
rect 262772 467168 262824 467220
rect 527180 467168 527232 467220
rect 4804 467100 4856 467152
rect 281724 467100 281776 467152
rect 299388 467100 299440 467152
rect 344560 467100 344612 467152
rect 275928 465876 275980 465928
rect 354404 465876 354456 465928
rect 218888 465808 218940 465860
rect 307300 465808 307352 465860
rect 258816 465740 258868 465792
rect 373264 465740 373316 465792
rect 21364 465672 21416 465724
rect 279792 465672 279844 465724
rect 291108 465672 291160 465724
rect 340696 465672 340748 465724
rect 246948 464448 247000 464500
rect 317788 464448 317840 464500
rect 218060 464380 218112 464432
rect 273260 464380 273312 464432
rect 274364 464380 274416 464432
rect 351828 464380 351880 464432
rect 266728 464312 266780 464364
rect 396724 464312 396776 464364
rect 324228 463156 324280 463208
rect 357716 463156 357768 463208
rect 252376 463088 252428 463140
rect 326252 463088 326304 463140
rect 255228 463020 255280 463072
rect 330852 463020 330904 463072
rect 260840 462952 260892 463004
rect 391204 462952 391256 463004
rect 3240 462340 3292 462392
rect 288992 462340 289044 462392
rect 211804 461796 211856 461848
rect 285036 461796 285088 461848
rect 262036 461728 262088 461780
rect 338672 461728 338724 461780
rect 268016 461660 268068 461712
rect 364340 461660 364392 461712
rect 71780 461592 71832 461644
rect 276480 461592 276532 461644
rect 288348 461592 288400 461644
rect 339408 461592 339460 461644
rect 250996 460436 251048 460488
rect 313188 460436 313240 460488
rect 239404 460368 239456 460420
rect 309232 460368 309284 460420
rect 277216 460300 277268 460352
rect 355692 460300 355744 460352
rect 265992 460232 266044 460284
rect 359464 460232 359516 460284
rect 98644 460164 98696 460216
rect 278504 460164 278556 460216
rect 215944 459008 215996 459060
rect 281080 459008 281132 459060
rect 260656 458940 260708 458992
rect 337384 458940 337436 458992
rect 140044 458872 140096 458924
rect 274548 458872 274600 458924
rect 281448 458872 281500 458924
rect 335452 458872 335504 458924
rect 264060 458804 264112 458856
rect 494060 458804 494112 458856
rect 249708 457580 249760 457632
rect 322296 457580 322348 457632
rect 256516 457512 256568 457564
rect 332140 457512 332192 457564
rect 28264 457444 28316 457496
rect 280436 457444 280488 457496
rect 306288 457444 306340 457496
rect 348516 457444 348568 457496
rect 252284 456764 252336 456816
rect 580172 456764 580224 456816
rect 201500 456220 201552 456272
rect 272616 456220 272668 456272
rect 259368 456152 259420 456204
rect 334808 456152 334860 456204
rect 262128 456084 262180 456136
rect 442264 456084 442316 456136
rect 88340 456016 88392 456068
rect 277124 456016 277176 456068
rect 277308 456016 277360 456068
rect 332784 456016 332836 456068
rect 268936 454860 268988 454912
rect 293224 454860 293276 454912
rect 296628 454860 296680 454912
rect 343272 454860 343324 454912
rect 244188 454792 244240 454844
rect 309876 454792 309928 454844
rect 260104 454724 260156 454776
rect 377404 454724 377456 454776
rect 40040 454656 40092 454708
rect 277860 454656 277912 454708
rect 278596 454656 278648 454708
rect 357072 454656 357124 454708
rect 214564 453568 214616 453620
rect 283012 453568 283064 453620
rect 251088 453500 251140 453552
rect 324320 453500 324372 453552
rect 271696 453432 271748 453484
rect 349160 453432 349212 453484
rect 169760 453364 169812 453416
rect 273904 453364 273956 453416
rect 258172 453296 258224 453348
rect 363604 453296 363656 453348
rect 252468 452140 252520 452192
rect 328276 452140 328328 452192
rect 210424 452072 210476 452124
rect 286968 452072 287020 452124
rect 273168 452004 273220 452056
rect 350540 452004 350592 452056
rect 255964 451936 256016 451988
rect 367744 451936 367796 451988
rect 108304 451868 108356 451920
rect 275836 451868 275888 451920
rect 278688 450712 278740 450764
rect 334164 450712 334216 450764
rect 254216 450644 254268 450696
rect 358084 450644 358136 450696
rect 261484 450576 261536 450628
rect 381544 450576 381596 450628
rect 25504 450508 25556 450560
rect 279148 450508 279200 450560
rect 245476 449692 245528 449744
rect 312544 449692 312596 449744
rect 245568 449624 245620 449676
rect 315120 449624 315172 449676
rect 267648 449556 267700 449608
rect 343916 449556 343968 449608
rect 266176 449488 266228 449540
rect 342628 449488 342680 449540
rect 263508 449420 263560 449472
rect 340052 449420 340104 449472
rect 264888 449352 264940 449404
rect 341340 449352 341392 449404
rect 269028 449284 269080 449336
rect 346584 449284 346636 449336
rect 270408 449216 270460 449268
rect 347872 449216 347924 449268
rect 267556 449148 267608 449200
rect 345296 449148 345348 449200
rect 303528 448060 303580 448112
rect 347228 448060 347280 448112
rect 284208 447992 284260 448044
rect 336740 447992 336792 448044
rect 237196 447924 237248 447976
rect 311900 447924 311952 447976
rect 260748 447856 260800 447908
rect 336096 447856 336148 447908
rect 217324 447788 217376 447840
rect 307944 447788 307996 447840
rect 267372 446632 267424 446684
rect 412640 446632 412692 446684
rect 265348 446564 265400 446616
rect 477500 446564 477552 446616
rect 263416 446496 263468 446548
rect 542360 446496 542412 446548
rect 4160 446428 4212 446480
rect 288256 446428 288308 446480
rect 259460 446360 259512 446412
rect 580264 446360 580316 446412
rect 203524 446156 203576 446208
rect 300124 446156 300176 446208
rect 199384 446088 199436 446140
rect 300768 446088 300820 446140
rect 200764 446020 200816 446072
rect 306012 446020 306064 446072
rect 250996 445952 251048 446004
rect 362592 445952 362644 446004
rect 249708 445884 249760 445936
rect 363604 445884 363656 445936
rect 235908 445816 235960 445868
rect 378784 445816 378836 445868
rect 82084 445748 82136 445800
rect 303988 445748 304040 445800
rect 231124 444932 231176 444984
rect 290280 444932 290332 444984
rect 225604 444864 225656 444916
rect 295524 444864 295576 444916
rect 215944 444796 215996 444848
rect 297456 444796 297508 444848
rect 245752 444728 245804 444780
rect 374644 444728 374696 444780
rect 240508 444660 240560 444712
rect 371976 444660 372028 444712
rect 100024 444592 100076 444644
rect 291568 444592 291620 444644
rect 95884 444524 95936 444576
rect 293500 444524 293552 444576
rect 7564 444456 7616 444508
rect 289636 444456 289688 444508
rect 244464 444388 244516 444440
rect 578884 444388 578936 444440
rect 355324 444320 355376 444372
rect 356428 444320 356480 444372
rect 356704 444320 356756 444372
rect 358360 444320 358412 444372
rect 248328 444116 248380 444168
rect 362408 444116 362460 444168
rect 245108 444048 245160 444100
rect 362224 444048 362276 444100
rect 334624 443980 334676 444032
rect 353760 443980 353812 444032
rect 243084 443912 243136 443964
rect 251180 443912 251232 443964
rect 333244 443912 333296 443964
rect 352472 443912 352524 443964
rect 94504 443844 94556 443896
rect 294880 443844 294932 443896
rect 301504 443844 301556 443896
rect 315764 443844 315816 443896
rect 331864 443844 331916 443896
rect 351184 443844 351236 443896
rect 230480 443776 230532 443828
rect 259460 443776 259512 443828
rect 294604 443776 294656 443828
rect 321008 443776 321060 443828
rect 336004 443776 336056 443828
rect 355048 443776 355100 443828
rect 219348 443708 219400 443760
rect 270592 443708 270644 443760
rect 297364 443708 297416 443760
rect 324964 443708 325016 443760
rect 329104 443708 329156 443760
rect 349804 443708 349856 443760
rect 217784 443640 217836 443692
rect 271972 443640 272024 443692
rect 293224 443640 293276 443692
rect 328920 443640 328972 443692
rect 338764 443640 338816 443692
rect 359004 443640 359056 443692
rect 243728 443572 243780 443624
rect 276112 443572 276164 443624
rect 251272 443504 251324 443556
rect 301412 443504 301464 443556
rect 229744 443436 229796 443488
rect 292856 443436 292908 443488
rect 228364 443368 228416 443420
rect 294144 443368 294196 443420
rect 239220 443300 239272 443352
rect 329748 443300 329800 443352
rect 196716 443232 196768 443284
rect 298744 443232 298796 443284
rect 250352 443164 250404 443216
rect 362500 443164 362552 443216
rect 237196 443096 237248 443148
rect 245568 443096 245620 443148
rect 359648 443096 359700 443148
rect 388444 443096 388496 443148
rect 276020 443028 276072 443080
rect 292212 443028 292264 443080
rect 360292 443028 360344 443080
rect 581092 443028 581144 443080
rect 235264 442960 235316 443012
rect 242900 442960 242952 443012
rect 246396 442960 246448 443012
rect 277400 442960 277452 443012
rect 280068 442960 280120 443012
rect 296168 442960 296220 443012
rect 360936 442960 360988 443012
rect 582380 442960 582432 443012
rect 329748 442620 329800 442672
rect 580724 442620 580776 442672
rect 3516 442552 3568 442604
rect 280068 442552 280120 442604
rect 300860 442552 300912 442604
rect 580632 442552 580684 442604
rect 3608 442484 3660 442536
rect 276020 442484 276072 442536
rect 279976 442484 280028 442536
rect 580264 442484 580316 442536
rect 276112 442416 276164 442468
rect 580816 442416 580868 442468
rect 251180 442348 251232 442400
rect 580908 442348 580960 442400
rect 245568 442280 245620 442332
rect 580540 442280 580592 442332
rect 242900 442212 242952 442264
rect 580448 442212 580500 442264
rect 231216 442144 231268 442196
rect 290924 442144 290976 442196
rect 206284 442076 206336 442128
rect 302056 442076 302108 442128
rect 198004 442008 198056 442060
rect 302700 442008 302752 442060
rect 192576 441940 192628 441992
rect 306656 441940 306708 441992
rect 248972 441872 249024 441924
rect 363696 441872 363748 441924
rect 140780 441804 140832 441856
rect 255964 441804 256016 441856
rect 247040 441736 247092 441788
rect 362316 441736 362368 441788
rect 8944 441668 8996 441720
rect 296812 441668 296864 441720
rect 241152 441600 241204 441652
rect 577596 441600 577648 441652
rect 283840 441192 283892 441244
rect 242348 441124 242400 441176
rect 248052 441124 248104 441176
rect 3424 440852 3476 440904
rect 251272 441056 251324 441108
rect 207664 440648 207716 440700
rect 242348 440988 242400 441040
rect 242716 440988 242768 441040
rect 247868 440988 247920 441040
rect 248052 440988 248104 441040
rect 252008 440988 252060 441040
rect 277400 440988 277452 441040
rect 283104 440988 283156 441040
rect 283564 440988 283616 441040
rect 283840 441056 283892 441108
rect 289268 441396 289320 441448
rect 284576 441328 284628 441380
rect 304908 441328 304960 441380
rect 284852 441260 284904 441312
rect 288900 441260 288952 441312
rect 284024 441192 284076 441244
rect 303068 441260 303120 441312
rect 298652 441192 298704 441244
rect 288900 441124 288952 441176
rect 284024 441056 284076 441108
rect 284576 440988 284628 441040
rect 284852 440988 284904 441040
rect 289268 440988 289320 441040
rect 88984 440376 89036 440428
rect 25504 440308 25556 440360
rect 304356 440988 304408 441040
rect 305000 440988 305052 441040
rect 580172 440852 580224 440904
rect 364984 440580 365036 440632
rect 377404 440512 377456 440564
rect 373356 440444 373408 440496
rect 97632 438132 97684 438184
rect 230480 438132 230532 438184
rect 362592 431876 362644 431928
rect 579804 431876 579856 431928
rect 3332 423580 3384 423632
rect 7564 423580 7616 423632
rect 364984 419432 365036 419484
rect 579988 419432 580040 419484
rect 3332 411204 3384 411256
rect 231216 411204 231268 411256
rect 362500 405628 362552 405680
rect 579804 405628 579856 405680
rect 3332 398760 3384 398812
rect 231124 398760 231176 398812
rect 363696 379448 363748 379500
rect 580080 379448 580132 379500
rect 3700 375980 3752 376032
rect 229744 375980 229796 376032
rect 154764 374892 154816 374944
rect 170404 374892 170456 374944
rect 116124 374824 116176 374876
rect 170956 374824 171008 374876
rect 103244 374756 103296 374808
rect 225696 374756 225748 374808
rect 100668 374688 100720 374740
rect 229836 374688 229888 374740
rect 147036 374620 147088 374672
rect 174728 374620 174780 374672
rect 139308 374552 139360 374604
rect 171784 374552 171836 374604
rect 121276 374484 121328 374536
rect 170772 374484 170824 374536
rect 165528 374416 165580 374468
rect 226984 374416 227036 374468
rect 167644 374348 167696 374400
rect 229744 374348 229796 374400
rect 108396 374280 108448 374332
rect 175924 374280 175976 374332
rect 131580 374212 131632 374264
rect 228456 374212 228508 374264
rect 126428 374144 126480 374196
rect 231124 374144 231176 374196
rect 162492 374008 162544 374060
rect 170496 374008 170548 374060
rect 32404 373056 32456 373108
rect 165068 373056 165120 373108
rect 165528 373056 165580 373108
rect 123852 372988 123904 373040
rect 170588 372988 170640 373040
rect 118700 372920 118752 372972
rect 174544 372920 174596 372972
rect 105820 372852 105872 372904
rect 174636 372852 174688 372904
rect 149612 372784 149664 372836
rect 228548 372784 228600 372836
rect 136732 372716 136784 372768
rect 224224 372716 224276 372768
rect 110972 372648 111024 372700
rect 228640 372648 228692 372700
rect 157340 372580 157392 372632
rect 173164 372580 173216 372632
rect 3332 372512 3384 372564
rect 100024 372512 100076 372564
rect 97816 371696 97868 371748
rect 97724 371628 97776 371680
rect 113456 371696 113508 371748
rect 115756 371696 115808 371748
rect 134064 371764 134116 371816
rect 133834 371696 133886 371748
rect 143172 371696 143224 371748
rect 144368 371696 144420 371748
rect 99840 371560 99892 371612
rect 97908 371492 97960 371544
rect 113456 371560 113508 371612
rect 113824 371560 113876 371612
rect 115756 371560 115808 371612
rect 129188 371560 129240 371612
rect 135168 371628 135220 371680
rect 145012 371628 145064 371680
rect 133834 371560 133886 371612
rect 143172 371560 143224 371612
rect 143264 371560 143316 371612
rect 144368 371560 144420 371612
rect 144736 371560 144788 371612
rect 144920 371560 144972 371612
rect 153016 371628 153068 371680
rect 152556 371560 152608 371612
rect 173256 371696 173308 371748
rect 229928 371628 229980 371680
rect 231216 371560 231268 371612
rect 231400 371492 231452 371544
rect 231308 371424 231360 371476
rect 230020 371356 230072 371408
rect 230112 371288 230164 371340
rect 231492 371220 231544 371272
rect 172336 368500 172388 368552
rect 227076 368500 227128 368552
rect 169944 367888 169996 367940
rect 170680 367888 170732 367940
rect 172428 365712 172480 365764
rect 231584 365712 231636 365764
rect 363604 365644 363656 365696
rect 580080 365644 580132 365696
rect 171692 357416 171744 357468
rect 228732 357416 228784 357468
rect 172428 354696 172480 354748
rect 230204 354696 230256 354748
rect 362408 353200 362460 353252
rect 579988 353200 580040 353252
rect 172428 351908 172480 351960
rect 227168 351908 227220 351960
rect 171692 350480 171744 350532
rect 171876 350480 171928 350532
rect 171140 349120 171192 349172
rect 171876 349120 171928 349172
rect 192484 349120 192536 349172
rect 172428 346400 172480 346452
rect 220084 346400 220136 346452
rect 172428 342252 172480 342304
rect 231676 342252 231728 342304
rect 172428 336744 172480 336796
rect 230296 336744 230348 336796
rect 172428 333956 172480 334008
rect 228824 333956 228876 334008
rect 172428 331236 172480 331288
rect 230388 331236 230440 331288
rect 172428 328448 172480 328500
rect 225788 328448 225840 328500
rect 171416 325660 171468 325712
rect 232228 325660 232280 325712
rect 362316 325592 362368 325644
rect 580080 325592 580132 325644
rect 172428 320152 172480 320204
rect 231768 320152 231820 320204
rect 3332 320084 3384 320136
rect 95884 320084 95936 320136
rect 172428 317432 172480 317484
rect 231860 317432 231912 317484
rect 172428 314644 172480 314696
rect 231952 314644 232004 314696
rect 377404 313216 377456 313268
rect 579988 313216 580040 313268
rect 230940 312944 230992 312996
rect 231308 312944 231360 312996
rect 231400 312672 231452 312724
rect 231676 312672 231728 312724
rect 172428 311856 172480 311908
rect 231860 311856 231912 311908
rect 231768 311788 231820 311840
rect 232044 311788 232096 311840
rect 172152 311312 172204 311364
rect 231032 311312 231084 311364
rect 171784 311244 171836 311296
rect 232136 311244 232188 311296
rect 171968 311176 172020 311228
rect 231768 311176 231820 311228
rect 192484 311108 192536 311160
rect 232228 311108 232280 311160
rect 171876 310564 171928 310616
rect 228824 310632 228876 310684
rect 226984 310496 227036 310548
rect 233148 310564 233200 310616
rect 232136 310496 232188 310548
rect 232780 310496 232832 310548
rect 233700 310496 233752 310548
rect 255412 310496 255464 310548
rect 255596 310496 255648 310548
rect 273536 310496 273588 310548
rect 273720 310496 273772 310548
rect 232596 310360 232648 310412
rect 231952 310292 232004 310344
rect 235540 310292 235592 310344
rect 231860 310224 231912 310276
rect 236276 310224 236328 310276
rect 230296 310156 230348 310208
rect 238944 310156 238996 310208
rect 172428 310020 172480 310072
rect 235908 310088 235960 310140
rect 231032 310020 231084 310072
rect 231952 310020 232004 310072
rect 172244 309952 172296 310004
rect 239496 309952 239548 310004
rect 232964 309884 233016 309936
rect 244464 309884 244516 309936
rect 230204 309816 230256 309868
rect 238760 309816 238812 309868
rect 230388 309612 230440 309664
rect 241796 309612 241848 309664
rect 228732 309476 228784 309528
rect 242992 309476 243044 309528
rect 231584 309408 231636 309460
rect 247500 309408 247552 309460
rect 315948 309408 316000 309460
rect 316408 309408 316460 309460
rect 232044 309340 232096 309392
rect 249616 309340 249668 309392
rect 231676 309272 231728 309324
rect 236552 309272 236604 309324
rect 231400 309204 231452 309256
rect 252836 309204 252888 309256
rect 170680 309136 170732 309188
rect 234160 309136 234212 309188
rect 236552 309136 236604 309188
rect 249800 309136 249852 309188
rect 354220 309136 354272 309188
rect 229928 309068 229980 309120
rect 233608 309068 233660 309120
rect 235816 309068 235868 309120
rect 238576 309068 238628 309120
rect 347688 309068 347740 309120
rect 231492 309000 231544 309052
rect 235356 309000 235408 309052
rect 348700 309000 348752 309052
rect 231216 308932 231268 308984
rect 235724 308932 235776 308984
rect 230020 308864 230072 308916
rect 238208 308864 238260 308916
rect 231860 308796 231912 308848
rect 241612 308864 241664 308916
rect 231952 308728 232004 308780
rect 245844 308796 245896 308848
rect 173164 308660 173216 308712
rect 248144 308728 248196 308780
rect 247960 308660 248012 308712
rect 254400 308660 254452 308712
rect 230940 308592 230992 308644
rect 240324 308592 240376 308644
rect 253204 308592 253256 308644
rect 262404 308932 262456 308984
rect 314844 308932 314896 308984
rect 315028 308932 315080 308984
rect 326712 308932 326764 308984
rect 338856 308932 338908 308984
rect 348516 308932 348568 308984
rect 352104 308932 352156 308984
rect 355692 309068 355744 309120
rect 367744 309068 367796 309120
rect 366272 309000 366324 309052
rect 170588 308524 170640 308576
rect 242348 308524 242400 308576
rect 250444 308524 250496 308576
rect 259000 308524 259052 308576
rect 253296 308456 253348 308508
rect 267004 308864 267056 308916
rect 310336 308864 310388 308916
rect 260380 308796 260432 308848
rect 268752 308796 268804 308848
rect 314660 308796 314712 308848
rect 315396 308796 315448 308848
rect 317420 308864 317472 308916
rect 317972 308864 318024 308916
rect 319076 308864 319128 308916
rect 319352 308864 319404 308916
rect 367652 308932 367704 308984
rect 303804 308728 303856 308780
rect 355232 308728 355284 308780
rect 371424 308864 371476 308916
rect 356520 308796 356572 308848
rect 357164 308728 357216 308780
rect 304540 308660 304592 308712
rect 355508 308660 355560 308712
rect 367376 308660 367428 308712
rect 260104 308592 260156 308644
rect 271604 308592 271656 308644
rect 302516 308592 302568 308644
rect 355692 308592 355744 308644
rect 356060 308592 356112 308644
rect 367560 308592 367612 308644
rect 271236 308524 271288 308576
rect 273444 308524 273496 308576
rect 302332 308524 302384 308576
rect 355600 308524 355652 308576
rect 357256 308524 357308 308576
rect 368572 308524 368624 308576
rect 267004 308456 267056 308508
rect 281264 308456 281316 308508
rect 301504 308456 301556 308508
rect 355416 308456 355468 308508
rect 360200 308456 360252 308508
rect 360844 308456 360896 308508
rect 224224 308388 224276 308440
rect 237012 308388 237064 308440
rect 174544 308320 174596 308372
rect 250352 308320 250404 308372
rect 228548 308252 228600 308304
rect 230112 308184 230164 308236
rect 242164 308184 242216 308236
rect 246764 308184 246816 308236
rect 246304 308116 246356 308168
rect 253480 308116 253532 308168
rect 252192 308048 252244 308100
rect 272708 308388 272760 308440
rect 301320 308388 301372 308440
rect 356520 308388 356572 308440
rect 356888 308388 356940 308440
rect 370044 308456 370096 308508
rect 312268 308320 312320 308372
rect 313004 308320 313056 308372
rect 313924 308320 313976 308372
rect 314936 308320 314988 308372
rect 315856 308320 315908 308372
rect 316132 308320 316184 308372
rect 316960 308320 317012 308372
rect 317604 308320 317656 308372
rect 318340 308320 318392 308372
rect 319168 308320 319220 308372
rect 319812 308320 319864 308372
rect 320180 308320 320232 308372
rect 321192 308320 321244 308372
rect 355324 308320 355376 308372
rect 367468 308320 367520 308372
rect 312176 308252 312228 308304
rect 312452 308252 312504 308304
rect 313372 308252 313424 308304
rect 314752 308252 314804 308304
rect 315672 308252 315724 308304
rect 316592 308252 316644 308304
rect 317696 308252 317748 308304
rect 317880 308252 317932 308304
rect 318984 308252 319036 308304
rect 319628 308252 319680 308304
rect 320364 308252 320416 308304
rect 320640 308252 320692 308304
rect 353852 308252 353904 308304
rect 366180 308252 366232 308304
rect 311900 308184 311952 308236
rect 313188 308184 313240 308236
rect 313280 308184 313332 308236
rect 314292 308184 314344 308236
rect 314660 308184 314712 308236
rect 315488 308184 315540 308236
rect 311992 308116 312044 308168
rect 312452 308116 312504 308168
rect 315028 308116 315080 308168
rect 315304 308116 315356 308168
rect 316224 308116 316276 308168
rect 317328 308184 317380 308236
rect 318064 308184 318116 308236
rect 318800 308184 318852 308236
rect 319444 308184 319496 308236
rect 354956 308184 355008 308236
rect 367284 308184 367336 308236
rect 317696 308116 317748 308168
rect 318708 308116 318760 308168
rect 318892 308116 318944 308168
rect 319996 308116 320048 308168
rect 320272 308116 320324 308168
rect 320640 308116 320692 308168
rect 354588 308116 354640 308168
rect 364800 308116 364852 308168
rect 259736 308048 259788 308100
rect 260012 308048 260064 308100
rect 317512 308048 317564 308100
rect 318524 308048 318576 308100
rect 245752 307980 245804 308032
rect 251916 307980 251968 308032
rect 269488 307980 269540 308032
rect 269764 307980 269816 308032
rect 285680 307980 285732 308032
rect 285956 307980 286008 308032
rect 311992 307980 312044 308032
rect 312820 307980 312872 308032
rect 316500 307980 316552 308032
rect 316776 307980 316828 308032
rect 320272 307980 320324 308032
rect 321376 307980 321428 308032
rect 360292 307980 360344 308032
rect 360660 307980 360712 308032
rect 251824 307912 251876 307964
rect 256516 307912 256568 307964
rect 317788 307912 317840 307964
rect 318156 307912 318208 307964
rect 320456 307912 320508 307964
rect 321008 307912 321060 307964
rect 360476 307912 360528 307964
rect 361212 307912 361264 307964
rect 244004 307844 244056 307896
rect 249248 307844 249300 307896
rect 250536 307844 250588 307896
rect 242808 307776 242860 307828
rect 243544 307776 243596 307828
rect 247776 307776 247828 307828
rect 248512 307776 248564 307828
rect 250904 307776 250956 307828
rect 251364 307776 251416 307828
rect 253388 307844 253440 307896
rect 259552 307844 259604 307896
rect 261760 307844 261812 307896
rect 269856 307844 269908 307896
rect 337016 307844 337068 307896
rect 337292 307844 337344 307896
rect 353392 307844 353444 307896
rect 360936 307844 360988 307896
rect 257804 307776 257856 307828
rect 348424 307776 348476 307828
rect 350356 307776 350408 307828
rect 353024 307776 353076 307828
rect 363512 307776 363564 307828
rect 227168 307708 227220 307760
rect 243728 307708 243780 307760
rect 225788 307640 225840 307692
rect 241980 307640 242032 307692
rect 229836 307572 229888 307624
rect 252284 307572 252336 307624
rect 175924 307504 175976 307556
rect 244832 307504 244884 307556
rect 220084 307436 220136 307488
rect 242532 307436 242584 307488
rect 229744 307368 229796 307420
rect 251732 307368 251784 307420
rect 228456 307300 228508 307352
rect 247132 307300 247184 307352
rect 315396 307300 315448 307352
rect 373264 307300 373316 307352
rect 172428 307232 172480 307284
rect 246948 307232 247000 307284
rect 313556 307232 313608 307284
rect 313832 307232 313884 307284
rect 317972 307232 318024 307284
rect 402980 307232 403032 307284
rect 170496 307164 170548 307216
rect 249984 307164 250036 307216
rect 295616 307164 295668 307216
rect 295892 307164 295944 307216
rect 323676 307164 323728 307216
rect 427084 307164 427136 307216
rect 170588 307096 170640 307148
rect 238392 307096 238444 307148
rect 313556 307096 313608 307148
rect 314476 307096 314528 307148
rect 330116 307096 330168 307148
rect 480260 307096 480312 307148
rect 200120 307028 200172 307080
rect 284944 307028 284996 307080
rect 316408 307028 316460 307080
rect 317144 307028 317196 307080
rect 340420 307028 340472 307080
rect 543740 307028 543792 307080
rect 170404 306960 170456 307012
rect 239680 306960 239732 307012
rect 262588 306960 262640 307012
rect 267924 306960 267976 307012
rect 276388 306960 276440 307012
rect 292764 306960 292816 307012
rect 293408 306960 293460 307012
rect 321836 306960 321888 307012
rect 322112 306960 322164 307012
rect 262680 306756 262732 306808
rect 268016 306756 268068 306808
rect 287060 306824 287112 306876
rect 287336 306824 287388 306876
rect 276480 306756 276532 306808
rect 277676 306688 277728 306740
rect 324412 306688 324464 306740
rect 325056 306688 325108 306740
rect 260840 306552 260892 306604
rect 261300 306552 261352 306604
rect 238944 306484 238996 306536
rect 239864 306484 239916 306536
rect 255320 306484 255372 306536
rect 255872 306484 255924 306536
rect 267832 306484 267884 306536
rect 268108 306484 268160 306536
rect 295800 306552 295852 306604
rect 327172 306552 327224 306604
rect 327632 306552 327684 306604
rect 357532 306552 357584 306604
rect 357992 306552 358044 306604
rect 278780 306484 278832 306536
rect 279792 306484 279844 306536
rect 282736 306484 282788 306536
rect 288532 306484 288584 306536
rect 294236 306484 294288 306536
rect 239036 306416 239088 306468
rect 240048 306416 240100 306468
rect 255504 306416 255556 306468
rect 255964 306416 256016 306468
rect 259552 306416 259604 306468
rect 260656 306416 260708 306468
rect 260932 306416 260984 306468
rect 261208 306416 261260 306468
rect 263600 306416 263652 306468
rect 263876 306416 263928 306468
rect 264152 306416 264204 306468
rect 264428 306416 264480 306468
rect 266636 306416 266688 306468
rect 266912 306416 266964 306468
rect 270684 306416 270736 306468
rect 270960 306416 271012 306468
rect 273720 306416 273772 306468
rect 274456 306416 274508 306468
rect 277676 306416 277728 306468
rect 279056 306416 279108 306468
rect 279424 306416 279476 306468
rect 280344 306416 280396 306468
rect 280804 306416 280856 306468
rect 286048 306416 286100 306468
rect 286232 306416 286284 306468
rect 237380 306348 237432 306400
rect 237932 306348 237984 306400
rect 238852 306348 238904 306400
rect 239312 306348 239364 306400
rect 240232 306348 240284 306400
rect 241428 306348 241480 306400
rect 243084 306348 243136 306400
rect 244096 306348 244148 306400
rect 248512 306348 248564 306400
rect 248880 306348 248932 306400
rect 249892 306348 249944 306400
rect 250996 306348 251048 306400
rect 251732 306348 251784 306400
rect 252100 306348 252152 306400
rect 252652 306348 252704 306400
rect 253664 306348 253716 306400
rect 255596 306348 255648 306400
rect 256148 306348 256200 306400
rect 256792 306348 256844 306400
rect 257988 306348 258040 306400
rect 259644 306348 259696 306400
rect 260472 306348 260524 306400
rect 261300 306348 261352 306400
rect 261852 306348 261904 306400
rect 264060 306348 264112 306400
rect 264888 306348 264940 306400
rect 265072 306348 265124 306400
rect 265256 306348 265308 306400
rect 265348 306348 265400 306400
rect 265624 306348 265676 306400
rect 267740 306348 267792 306400
rect 268108 306348 268160 306400
rect 269212 306348 269264 306400
rect 270224 306348 270276 306400
rect 272248 306348 272300 306400
rect 273076 306348 273128 306400
rect 273628 306348 273680 306400
rect 274088 306348 274140 306400
rect 274916 306348 274968 306400
rect 275560 306348 275612 306400
rect 276112 306348 276164 306400
rect 277308 306348 277360 306400
rect 277400 306348 277452 306400
rect 278412 306348 278464 306400
rect 278872 306348 278924 306400
rect 279148 306348 279200 306400
rect 282920 306348 282972 306400
rect 283748 306348 283800 306400
rect 284392 306348 284444 306400
rect 285128 306348 285180 306400
rect 285680 306348 285732 306400
rect 3332 306280 3384 306332
rect 94504 306280 94556 306332
rect 219072 306280 219124 306332
rect 284208 306280 284260 306332
rect 284668 306280 284720 306332
rect 285496 306280 285548 306332
rect 287428 306280 287480 306332
rect 291568 306280 291620 306332
rect 292212 306280 292264 306332
rect 293132 306280 293184 306332
rect 293684 306280 293736 306332
rect 296720 306484 296772 306536
rect 297180 306484 297232 306536
rect 296904 306416 296956 306468
rect 297364 306416 297416 306468
rect 306840 306416 306892 306468
rect 310612 306416 310664 306468
rect 310888 306416 310940 306468
rect 325792 306416 325844 306468
rect 326436 306416 326488 306468
rect 328552 306416 328604 306468
rect 329380 306416 329432 306468
rect 331312 306416 331364 306468
rect 331772 306416 331824 306468
rect 336832 306416 336884 306468
rect 337200 306416 337252 306468
rect 339684 306416 339736 306468
rect 339960 306416 340012 306468
rect 340880 306416 340932 306468
rect 341432 306416 341484 306468
rect 345020 306416 345072 306468
rect 345480 306416 345532 306468
rect 295800 306348 295852 306400
rect 299664 306348 299716 306400
rect 300400 306348 300452 306400
rect 300860 306348 300912 306400
rect 301688 306348 301740 306400
rect 302424 306348 302476 306400
rect 303252 306348 303304 306400
rect 303804 306348 303856 306400
rect 304632 306348 304684 306400
rect 295524 306280 295576 306332
rect 295984 306280 296036 306332
rect 298100 306280 298152 306332
rect 298652 306280 298704 306332
rect 299572 306280 299624 306332
rect 300216 306280 300268 306332
rect 302516 306280 302568 306332
rect 303068 306280 303120 306332
rect 303712 306280 303764 306332
rect 304356 306280 304408 306332
rect 216496 306212 216548 306264
rect 171692 306144 171744 306196
rect 245476 306144 245528 306196
rect 247224 306144 247276 306196
rect 247868 306144 247920 306196
rect 251364 306144 251416 306196
rect 252468 306144 252520 306196
rect 254032 306144 254084 306196
rect 254768 306144 254820 306196
rect 255688 306144 255740 306196
rect 256332 306144 256384 306196
rect 258080 306144 258132 306196
rect 258540 306144 258592 306196
rect 259736 306144 259788 306196
rect 260288 306144 260340 306196
rect 262588 306144 262640 306196
rect 263324 306144 263376 306196
rect 263692 306144 263744 306196
rect 264520 306144 264572 306196
rect 266728 306144 266780 306196
rect 267372 306144 267424 306196
rect 267924 306144 267976 306196
rect 268292 306144 268344 306196
rect 269120 306144 269172 306196
rect 269488 306144 269540 306196
rect 270868 306144 270920 306196
rect 271052 306144 271104 306196
rect 271972 306144 272024 306196
rect 272524 306144 272576 306196
rect 273352 306144 273404 306196
rect 274272 306144 274324 306196
rect 277492 306144 277544 306196
rect 277860 306144 277912 306196
rect 279240 306144 279292 306196
rect 279976 306144 280028 306196
rect 280068 306144 280120 306196
rect 281540 306144 281592 306196
rect 283380 306212 283432 306264
rect 284024 306212 284076 306264
rect 284576 306212 284628 306264
rect 285312 306212 285364 306264
rect 285864 306212 285916 306264
rect 286140 306212 286192 306264
rect 286876 306212 286928 306264
rect 287152 306212 287204 306264
rect 287244 306212 287296 306264
rect 287980 306212 288032 306264
rect 294236 306212 294288 306264
rect 297180 306212 297232 306264
rect 297916 306212 297968 306264
rect 300952 306212 301004 306264
rect 302056 306212 302108 306264
rect 302332 306212 302384 306264
rect 303436 306212 303488 306264
rect 305460 306212 305512 306264
rect 305920 306212 305972 306264
rect 306656 306212 306708 306264
rect 328736 306348 328788 306400
rect 329564 306348 329616 306400
rect 329840 306348 329892 306400
rect 331128 306348 331180 306400
rect 331220 306348 331272 306400
rect 332232 306348 332284 306400
rect 332600 306348 332652 306400
rect 332876 306348 332928 306400
rect 333060 306348 333112 306400
rect 333612 306348 333664 306400
rect 335360 306348 335412 306400
rect 336096 306348 336148 306400
rect 336740 306348 336792 306400
rect 337384 306348 337436 306400
rect 345112 306348 345164 306400
rect 346216 306348 346268 306400
rect 347780 306348 347832 306400
rect 349068 306348 349120 306400
rect 307944 306280 307996 306332
rect 308956 306280 309008 306332
rect 310980 306280 311032 306332
rect 311440 306280 311492 306332
rect 321836 306280 321888 306332
rect 322664 306280 322716 306332
rect 325700 306280 325752 306332
rect 326160 306280 326212 306332
rect 327540 306280 327592 306332
rect 327816 306280 327868 306332
rect 328644 306280 328696 306332
rect 329104 306280 329156 306332
rect 329932 306280 329984 306332
rect 330944 306280 330996 306332
rect 331312 306280 331364 306332
rect 332048 306280 332100 306332
rect 332968 306280 333020 306332
rect 333244 306280 333296 306332
rect 335544 306280 335596 306332
rect 336280 306280 336332 306332
rect 336924 306280 336976 306332
rect 337752 306280 337804 306332
rect 338120 306280 338172 306332
rect 338948 306280 339000 306332
rect 342260 306280 342312 306332
rect 342904 306280 342956 306332
rect 343824 306280 343876 306332
rect 344284 306280 344336 306332
rect 345020 306280 345072 306332
rect 345756 306280 345808 306332
rect 347872 306280 347924 306332
rect 348240 306280 348292 306332
rect 350540 306280 350592 306332
rect 351552 306280 351604 306332
rect 353208 306280 353260 306332
rect 362316 306484 362368 306536
rect 357624 306416 357676 306468
rect 308036 306212 308088 306264
rect 308588 306212 308640 306264
rect 311072 306212 311124 306264
rect 311624 306212 311676 306264
rect 321560 306212 321612 306264
rect 322020 306212 322072 306264
rect 322940 306212 322992 306264
rect 323492 306212 323544 306264
rect 325884 306212 325936 306264
rect 326896 306212 326948 306264
rect 328828 306212 328880 306264
rect 329012 306212 329064 306264
rect 332600 306212 332652 306264
rect 333796 306212 333848 306264
rect 335452 306212 335504 306264
rect 336648 306212 336700 306264
rect 336832 306212 336884 306264
rect 337936 306212 337988 306264
rect 338488 306212 338540 306264
rect 339316 306212 339368 306264
rect 339684 306212 339736 306264
rect 340052 306212 340104 306264
rect 341064 306212 341116 306264
rect 341432 306212 341484 306264
rect 342720 306212 342772 306264
rect 343272 306212 343324 306264
rect 289084 306144 289136 306196
rect 295708 306144 295760 306196
rect 296536 306144 296588 306196
rect 301044 306144 301096 306196
rect 301872 306144 301924 306196
rect 303988 306144 304040 306196
rect 305368 306144 305420 306196
rect 305736 306144 305788 306196
rect 306380 306144 306432 306196
rect 306840 306144 306892 306196
rect 307852 306144 307904 306196
rect 308404 306144 308456 306196
rect 310704 306144 310756 306196
rect 311348 306144 311400 306196
rect 321744 306144 321796 306196
rect 322480 306144 322532 306196
rect 324596 306144 324648 306196
rect 325608 306144 325660 306196
rect 328644 306144 328696 306196
rect 329196 306144 329248 306196
rect 332784 306144 332836 306196
rect 333428 306144 333480 306196
rect 333980 306144 334032 306196
rect 334440 306144 334492 306196
rect 334532 306144 334584 306196
rect 334900 306144 334952 306196
rect 338212 306144 338264 306196
rect 338672 306144 338724 306196
rect 339500 306144 339552 306196
rect 340236 306144 340288 306196
rect 340972 306144 341024 306196
rect 341524 306144 341576 306196
rect 215208 306076 215260 306128
rect 282736 306076 282788 306128
rect 295616 306076 295668 306128
rect 296352 306076 296404 306128
rect 219164 306008 219216 306060
rect 282552 306008 282604 306060
rect 283656 306008 283708 306060
rect 293500 306008 293552 306060
rect 305000 306076 305052 306128
rect 305644 306076 305696 306128
rect 306564 306076 306616 306128
rect 307300 306076 307352 306128
rect 309232 306076 309284 306128
rect 309692 306076 309744 306128
rect 310796 306076 310848 306128
rect 311808 306076 311860 306128
rect 321560 306076 321612 306128
rect 322296 306076 322348 306128
rect 323216 306076 323268 306128
rect 324044 306076 324096 306128
rect 324504 306076 324556 306128
rect 325240 306076 325292 306128
rect 327172 306076 327224 306128
rect 327908 306076 327960 306128
rect 328460 306076 328512 306128
rect 329012 306076 329064 306128
rect 334164 306076 334216 306128
rect 335084 306076 335136 306128
rect 339592 306076 339644 306128
rect 340604 306076 340656 306128
rect 341064 306076 341116 306128
rect 341800 306076 341852 306128
rect 342444 306076 342496 306128
rect 343088 306076 343140 306128
rect 305092 306008 305144 306060
rect 306288 306008 306340 306060
rect 306380 306008 306432 306060
rect 307208 306008 307260 306060
rect 309140 306008 309192 306060
rect 309600 306008 309652 306060
rect 323124 306008 323176 306060
rect 323860 306008 323912 306060
rect 327264 306008 327316 306060
rect 328276 306008 328328 306060
rect 334440 306008 334492 306060
rect 335268 306008 335320 306060
rect 338212 306008 338264 306060
rect 339132 306008 339184 306060
rect 340972 306008 341024 306060
rect 341984 306008 342036 306060
rect 342352 306008 342404 306060
rect 343364 306008 343416 306060
rect 345296 306212 345348 306264
rect 356520 306212 356572 306264
rect 356796 306212 356848 306264
rect 357808 306348 357860 306400
rect 357992 306348 358044 306400
rect 359648 306348 359700 306400
rect 366364 306280 366416 306332
rect 357716 306212 357768 306264
rect 356336 306144 356388 306196
rect 371608 306212 371660 306264
rect 357440 306076 357492 306128
rect 357900 306076 357952 306128
rect 354036 306008 354088 306060
rect 368940 306144 368992 306196
rect 359280 306076 359332 306128
rect 359740 306076 359792 306128
rect 359832 306076 359884 306128
rect 369032 306076 369084 306128
rect 359372 306008 359424 306060
rect 359924 306008 359976 306060
rect 362316 306008 362368 306060
rect 368756 306008 368808 306060
rect 214932 305940 214984 305992
rect 282368 305940 282420 305992
rect 284208 305940 284260 305992
rect 291844 305940 291896 305992
rect 303988 305940 304040 305992
rect 328460 305940 328512 305992
rect 329748 305940 329800 305992
rect 343916 305940 343968 305992
rect 344192 305940 344244 305992
rect 345204 305940 345256 305992
rect 345296 305940 345348 305992
rect 345848 305940 345900 305992
rect 354772 305940 354824 305992
rect 371516 305940 371568 305992
rect 216312 305872 216364 305924
rect 282736 305872 282788 305924
rect 284944 305872 284996 305924
rect 292672 305872 292724 305924
rect 355140 305872 355192 305924
rect 371792 305872 371844 305924
rect 213828 305804 213880 305856
rect 170404 305736 170456 305788
rect 255136 305736 255188 305788
rect 256976 305736 257028 305788
rect 257620 305736 257672 305788
rect 258264 305736 258316 305788
rect 258816 305736 258868 305788
rect 261024 305736 261076 305788
rect 261484 305736 261536 305788
rect 262312 305736 262364 305788
rect 263140 305736 263192 305788
rect 263968 305736 264020 305788
rect 264704 305736 264756 305788
rect 266820 305736 266872 305788
rect 267556 305736 267608 305788
rect 270776 305736 270828 305788
rect 271420 305736 271472 305788
rect 277584 305804 277636 305856
rect 278228 305804 278280 305856
rect 278872 305804 278924 305856
rect 279608 305804 279660 305856
rect 280436 305804 280488 305856
rect 281080 305804 281132 305856
rect 281816 305804 281868 305856
rect 282276 305804 282328 305856
rect 294696 305804 294748 305856
rect 343916 305804 343968 305856
rect 344652 305804 344704 305856
rect 353576 305804 353628 305856
rect 359832 305804 359884 305856
rect 359924 305804 359976 305856
rect 369124 305804 369176 305856
rect 284852 305736 284904 305788
rect 292396 305736 292448 305788
rect 354404 305736 354456 305788
rect 371700 305736 371752 305788
rect 195980 305668 196032 305720
rect 284300 305668 284352 305720
rect 287428 305668 287480 305720
rect 287796 305668 287848 305720
rect 293040 305668 293092 305720
rect 293868 305668 293920 305720
rect 351184 305668 351236 305720
rect 359648 305668 359700 305720
rect 359740 305668 359792 305720
rect 370228 305668 370280 305720
rect 178040 305600 178092 305652
rect 280068 305600 280120 305652
rect 280252 305600 280304 305652
rect 280896 305600 280948 305652
rect 281724 305600 281776 305652
rect 282828 305600 282880 305652
rect 283196 305600 283248 305652
rect 283932 305600 283984 305652
rect 298192 305600 298244 305652
rect 299204 305600 299256 305652
rect 347136 305600 347188 305652
rect 370412 305600 370464 305652
rect 218980 305532 219032 305584
rect 290648 305532 290700 305584
rect 352288 305532 352340 305584
rect 359924 305532 359976 305584
rect 360016 305532 360068 305584
rect 363604 305532 363656 305584
rect 218888 305464 218940 305516
rect 289544 305464 289596 305516
rect 309324 305464 309376 305516
rect 310152 305464 310204 305516
rect 355784 305464 355836 305516
rect 365076 305464 365128 305516
rect 172152 305396 172204 305448
rect 235172 305396 235224 305448
rect 235908 305396 235960 305448
rect 236644 305396 236696 305448
rect 247684 305396 247736 305448
rect 247960 305396 248012 305448
rect 256884 305396 256936 305448
rect 257436 305396 257488 305448
rect 261116 305396 261168 305448
rect 262036 305396 262088 305448
rect 266452 305396 266504 305448
rect 267188 305396 267240 305448
rect 271052 305396 271104 305448
rect 271788 305396 271840 305448
rect 276388 305396 276440 305448
rect 276940 305396 276992 305448
rect 280160 305396 280212 305448
rect 280528 305396 280580 305448
rect 282736 305396 282788 305448
rect 284944 305396 284996 305448
rect 349436 305396 349488 305448
rect 97448 305328 97500 305380
rect 256700 305328 256752 305380
rect 257344 305328 257396 305380
rect 282368 305328 282420 305380
rect 284852 305328 284904 305380
rect 359188 305396 359240 305448
rect 360108 305396 360160 305448
rect 359556 305328 359608 305380
rect 352656 305260 352708 305312
rect 360016 305260 360068 305312
rect 343640 305192 343692 305244
rect 344836 305192 344888 305244
rect 351736 305192 351788 305244
rect 359740 305192 359792 305244
rect 97448 305124 97500 305176
rect 276020 305056 276072 305108
rect 277124 305056 277176 305108
rect 97632 304920 97684 304972
rect 97908 304920 97960 304972
rect 172336 304920 172388 304972
rect 245200 304920 245252 304972
rect 294144 304852 294196 304904
rect 294328 304852 294380 304904
rect 294328 304716 294380 304768
rect 295064 304716 295116 304768
rect 258356 304648 258408 304700
rect 259184 304648 259236 304700
rect 264980 304648 265032 304700
rect 265900 304648 265952 304700
rect 169944 304580 169996 304632
rect 237196 304580 237248 304632
rect 274640 304580 274692 304632
rect 275744 304580 275796 304632
rect 169852 304512 169904 304564
rect 243176 304512 243228 304564
rect 290188 304512 290240 304564
rect 291016 304512 291068 304564
rect 172244 304444 172296 304496
rect 246028 304444 246080 304496
rect 324228 304444 324280 304496
rect 440884 304444 440936 304496
rect 171416 304376 171468 304428
rect 249432 304376 249484 304428
rect 250352 304376 250404 304428
rect 250812 304376 250864 304428
rect 299940 304376 299992 304428
rect 300768 304376 300820 304428
rect 326436 304376 326488 304428
rect 452660 304376 452712 304428
rect 207020 304308 207072 304360
rect 285680 304308 285732 304360
rect 331772 304308 331824 304360
rect 485044 304308 485096 304360
rect 189080 304240 189132 304292
rect 283104 304240 283156 304292
rect 303896 304240 303948 304292
rect 304172 304240 304224 304292
rect 335912 304240 335964 304292
rect 514024 304240 514076 304292
rect 252744 304172 252796 304224
rect 253112 304172 253164 304224
rect 262496 304172 262548 304224
rect 262772 304172 262824 304224
rect 295340 304172 295392 304224
rect 296168 304172 296220 304224
rect 252928 303832 252980 303884
rect 253848 303832 253900 303884
rect 269304 303696 269356 303748
rect 270408 303696 270460 303748
rect 265164 303628 265216 303680
rect 266268 303628 266320 303680
rect 217968 303560 218020 303612
rect 292856 303560 292908 303612
rect 355876 303560 355928 303612
rect 372068 303560 372120 303612
rect 216404 303492 216456 303544
rect 291384 303492 291436 303544
rect 347964 303492 348016 303544
rect 367928 303492 367980 303544
rect 214840 303424 214892 303476
rect 290832 303424 290884 303476
rect 352472 303424 352524 303476
rect 372804 303424 372856 303476
rect 212448 303356 212500 303408
rect 289360 303356 289412 303408
rect 350172 303356 350224 303408
rect 370596 303356 370648 303408
rect 219256 303288 219308 303340
rect 295432 303288 295484 303340
rect 352840 303288 352892 303340
rect 374184 303288 374236 303340
rect 216220 303220 216272 303272
rect 292580 303220 292632 303272
rect 351920 303220 351972 303272
rect 374368 303220 374420 303272
rect 214564 303152 214616 303204
rect 292028 303152 292080 303204
rect 299848 303152 299900 303204
rect 300584 303152 300636 303204
rect 348884 303152 348936 303204
rect 372988 303152 373040 303204
rect 212080 303084 212132 303136
rect 289912 303084 289964 303136
rect 349620 303084 349672 303136
rect 374276 303084 374328 303136
rect 169760 303016 169812 303068
rect 251548 303016 251600 303068
rect 301136 303016 301188 303068
rect 363696 303016 363748 303068
rect 213644 302948 213696 303000
rect 294052 302948 294104 303000
rect 298376 302948 298428 303000
rect 367100 302948 367152 303000
rect 184940 302880 184992 302932
rect 282644 302880 282696 302932
rect 298836 302880 298888 302932
rect 367836 302880 367888 302932
rect 214656 302812 214708 302864
rect 289728 302812 289780 302864
rect 350724 302812 350776 302864
rect 366456 302812 366508 302864
rect 216128 302744 216180 302796
rect 290280 302744 290332 302796
rect 341156 302744 341208 302796
rect 342168 302744 342220 302796
rect 356612 302744 356664 302796
rect 370688 302744 370740 302796
rect 214748 302676 214800 302728
rect 288164 302676 288216 302728
rect 351368 302676 351420 302728
rect 362316 302676 362368 302728
rect 269580 302472 269632 302524
rect 270040 302472 270092 302524
rect 334256 302472 334308 302524
rect 334716 302472 334768 302524
rect 236460 302268 236512 302320
rect 236184 302200 236236 302252
rect 172428 302132 172480 302184
rect 240140 302132 240192 302184
rect 210976 301724 211028 301776
rect 295340 301724 295392 301776
rect 212172 301656 212224 301708
rect 296812 301656 296864 301708
rect 312268 301656 312320 301708
rect 374000 301656 374052 301708
rect 211896 301588 211948 301640
rect 347964 301588 348016 301640
rect 358820 301588 358872 301640
rect 359004 301588 359056 301640
rect 171784 301520 171836 301572
rect 257344 301520 257396 301572
rect 331588 301520 331640 301572
rect 494060 301520 494112 301572
rect 193220 301452 193272 301504
rect 282920 301452 282972 301504
rect 338672 301452 338724 301504
rect 529940 301452 529992 301504
rect 276296 300840 276348 300892
rect 276572 300840 276624 300892
rect 97448 300772 97500 300824
rect 249984 300772 250036 300824
rect 99104 300704 99156 300756
rect 251364 300704 251416 300756
rect 97080 300636 97132 300688
rect 245752 300636 245804 300688
rect 313832 300636 313884 300688
rect 376760 300636 376812 300688
rect 97816 300568 97868 300620
rect 246212 300568 246264 300620
rect 298284 300568 298336 300620
rect 365168 300568 365220 300620
rect 99380 300500 99432 300552
rect 247132 300500 247184 300552
rect 299848 300500 299900 300552
rect 369216 300500 369268 300552
rect 97908 300432 97960 300484
rect 242808 300432 242860 300484
rect 301136 300432 301188 300484
rect 370504 300432 370556 300484
rect 98920 300364 98972 300416
rect 243360 300364 243412 300416
rect 299940 300364 299992 300416
rect 372896 300364 372948 300416
rect 97724 300296 97776 300348
rect 242716 300296 242768 300348
rect 320824 300296 320876 300348
rect 422300 300296 422352 300348
rect 99840 300228 99892 300280
rect 240416 300228 240468 300280
rect 333152 300228 333204 300280
rect 498292 300228 498344 300280
rect 99472 300160 99524 300212
rect 241060 300160 241112 300212
rect 339868 300160 339920 300212
rect 538864 300160 538916 300212
rect 97632 300092 97684 300144
rect 237564 300092 237616 300144
rect 341524 300092 341576 300144
rect 545764 300092 545816 300144
rect 98828 300024 98880 300076
rect 233332 300024 233384 300076
rect 205640 299956 205692 300008
rect 285772 299956 285824 300008
rect 213368 299888 213420 299940
rect 290280 299888 290332 299940
rect 99012 299412 99064 299464
rect 240508 299412 240560 299464
rect 98644 299344 98696 299396
rect 240232 299344 240284 299396
rect 98552 299276 98604 299328
rect 238944 299276 238996 299328
rect 104532 299208 104584 299260
rect 234988 299208 235040 299260
rect 114836 299140 114888 299192
rect 244464 299140 244516 299192
rect 119988 299072 120040 299124
rect 247224 299072 247276 299124
rect 117412 299004 117464 299056
rect 243084 299004 243136 299056
rect 130292 298936 130344 298988
rect 250352 298936 250404 298988
rect 319352 298936 319404 298988
rect 377404 298936 377456 298988
rect 125140 298868 125192 298920
rect 238852 298868 238904 298920
rect 315120 298868 315172 298920
rect 385040 298868 385092 298920
rect 140596 298800 140648 298852
rect 250628 298800 250680 298852
rect 333060 298800 333112 298852
rect 500224 298800 500276 298852
rect 156052 298732 156104 298784
rect 251732 298732 251784 298784
rect 341432 298732 341484 298784
rect 547972 298732 548024 298784
rect 145748 298664 145800 298716
rect 236184 298664 236236 298716
rect 161204 298596 161256 298648
rect 247776 298596 247828 298648
rect 163780 298528 163832 298580
rect 234712 298528 234764 298580
rect 158628 298052 158680 298104
rect 166356 298052 166408 298104
rect 170588 298052 170640 298104
rect 169852 297984 169904 298036
rect 132868 297916 132920 297968
rect 251456 297916 251508 297968
rect 122564 297848 122616 297900
rect 237932 297848 237984 297900
rect 138020 297780 138072 297832
rect 239128 297780 239180 297832
rect 148324 297712 148376 297764
rect 236276 297712 236328 297764
rect 100024 297644 100076 297696
rect 172244 297644 172296 297696
rect 214472 297644 214524 297696
rect 294420 297644 294472 297696
rect 322204 297644 322256 297696
rect 381544 297644 381596 297696
rect 101956 297576 102008 297628
rect 171416 297576 171468 297628
rect 213736 297576 213788 297628
rect 294236 297576 294288 297628
rect 319260 297576 319312 297628
rect 412640 297576 412692 297628
rect 107108 297508 107160 297560
rect 169944 297508 169996 297560
rect 213276 297508 213328 297560
rect 346584 297508 346636 297560
rect 135444 297440 135496 297492
rect 171692 297440 171744 297492
rect 210884 297440 210936 297492
rect 293040 297440 293092 297492
rect 327632 297440 327684 297492
rect 463700 297440 463752 297492
rect 143172 297372 143224 297424
rect 211712 297372 211764 297424
rect 294144 297372 294196 297424
rect 342812 297372 342864 297424
rect 557540 297372 557592 297424
rect 172152 297304 172204 297356
rect 213460 297304 213512 297356
rect 293132 297304 293184 297356
rect 215852 297236 215904 297288
rect 295248 297236 295300 297288
rect 216036 297168 216088 297220
rect 293224 297168 293276 297220
rect 98736 297100 98788 297152
rect 236368 297100 236420 297152
rect 112260 297032 112312 297084
rect 235908 297032 235960 297084
rect 126980 296624 127032 296676
rect 243544 296624 243596 296676
rect 153200 296556 153252 296608
rect 248604 296556 248656 296608
rect 209780 296216 209832 296268
rect 286232 296216 286284 296268
rect 129740 296148 129792 296200
rect 273812 296148 273864 296200
rect 318064 296148 318116 296200
rect 400220 296148 400272 296200
rect 125600 296080 125652 296132
rect 272432 296080 272484 296132
rect 322020 296080 322072 296132
rect 421564 296080 421616 296132
rect 63500 296012 63552 296064
rect 262772 296012 262824 296064
rect 335820 296012 335872 296064
rect 516784 296012 516836 296064
rect 16580 295944 16632 295996
rect 255872 295944 255924 295996
rect 344192 295944 344244 295996
rect 563704 295944 563756 295996
rect 217876 295264 217928 295316
rect 296996 295264 297048 295316
rect 215760 295196 215812 295248
rect 297088 295196 297140 295248
rect 215116 295128 215168 295180
rect 296904 295128 296956 295180
rect 214380 295060 214432 295112
rect 296720 295060 296772 295112
rect 212264 294992 212316 295044
rect 295708 294992 295760 295044
rect 211068 294924 211120 294976
rect 295524 294924 295576 294976
rect 210700 294856 210752 294908
rect 295800 294856 295852 294908
rect 210792 294788 210844 294840
rect 295616 294788 295668 294840
rect 168380 294720 168432 294772
rect 278780 294720 278832 294772
rect 313740 294720 313792 294772
rect 380900 294720 380952 294772
rect 135260 294652 135312 294704
rect 274732 294652 274784 294704
rect 329104 294652 329156 294704
rect 468484 294652 468536 294704
rect 43444 294584 43496 294636
rect 258448 294584 258500 294636
rect 337200 294584 337252 294636
rect 525800 294584 525852 294636
rect 215024 294516 215076 294568
rect 294328 294516 294380 294568
rect 218796 294448 218848 294500
rect 295892 294448 295944 294500
rect 3332 293904 3384 293956
rect 228364 293904 228416 293956
rect 317788 293496 317840 293548
rect 405740 293496 405792 293548
rect 218704 293428 218756 293480
rect 349712 293428 349764 293480
rect 202880 293360 202932 293412
rect 284668 293360 284720 293412
rect 329012 293360 329064 293412
rect 467104 293360 467156 293412
rect 71044 293292 71096 293344
rect 263600 293292 263652 293344
rect 335728 293292 335780 293344
rect 509884 293292 509936 293344
rect 52460 293224 52512 293276
rect 260840 293224 260892 293276
rect 338580 293224 338632 293276
rect 527824 293224 527876 293276
rect 315028 292000 315080 292052
rect 387064 292000 387116 292052
rect 161480 291932 161532 291984
rect 279148 291932 279200 291984
rect 327540 291932 327592 291984
rect 464344 291932 464396 291984
rect 128360 291864 128412 291916
rect 271144 291864 271196 291916
rect 330116 291864 330168 291916
rect 478144 291864 478196 291916
rect 22100 291796 22152 291848
rect 255688 291796 255740 291848
rect 338488 291796 338540 291848
rect 534724 291796 534776 291848
rect 151820 290708 151872 290760
rect 276020 290708 276072 290760
rect 317696 290708 317748 290760
rect 408500 290708 408552 290760
rect 217692 290640 217744 290692
rect 348516 290640 348568 290692
rect 143540 290572 143592 290624
rect 274640 290572 274692 290624
rect 320640 290572 320692 290624
rect 418160 290572 418212 290624
rect 44180 290504 44232 290556
rect 259828 290504 259880 290556
rect 341248 290504 341300 290556
rect 543004 290504 543056 290556
rect 13084 290436 13136 290488
rect 254308 290436 254360 290488
rect 341340 290436 341392 290488
rect 549904 290436 549956 290488
rect 201500 289280 201552 289332
rect 284576 289280 284628 289332
rect 132500 289212 132552 289264
rect 273628 289212 273680 289264
rect 321928 289212 321980 289264
rect 430580 289212 430632 289264
rect 103520 289144 103572 289196
rect 269764 289144 269816 289196
rect 331496 289144 331548 289196
rect 490012 289144 490064 289196
rect 9680 289076 9732 289128
rect 254216 289076 254268 289128
rect 341156 289076 341208 289128
rect 552664 289076 552716 289128
rect 181444 287784 181496 287836
rect 281908 287784 281960 287836
rect 327448 287784 327500 287836
rect 460204 287784 460256 287836
rect 139400 287716 139452 287768
rect 275100 287716 275152 287768
rect 342628 287716 342680 287768
rect 554044 287716 554096 287768
rect 27620 287648 27672 287700
rect 257160 287648 257212 287700
rect 342720 287648 342772 287700
rect 561680 287648 561732 287700
rect 312176 286560 312228 286612
rect 371240 286560 371292 286612
rect 199476 286492 199528 286544
rect 283288 286492 283340 286544
rect 323400 286492 323452 286544
rect 435364 286492 435416 286544
rect 146300 286424 146352 286476
rect 276480 286424 276532 286476
rect 324872 286424 324924 286476
rect 448520 286424 448572 286476
rect 46940 286356 46992 286408
rect 259736 286356 259788 286408
rect 328920 286356 328972 286408
rect 471980 286356 472032 286408
rect 8300 286288 8352 286340
rect 254124 286288 254176 286340
rect 344100 286288 344152 286340
rect 566464 286288 566516 286340
rect 150440 285132 150492 285184
rect 276388 285132 276440 285184
rect 313648 285132 313700 285184
rect 378140 285132 378192 285184
rect 81440 285064 81492 285116
rect 265532 285064 265584 285116
rect 313556 285064 313608 285116
rect 382280 285064 382332 285116
rect 40040 284996 40092 285048
rect 258356 284996 258408 285048
rect 323308 284996 323360 285048
rect 436100 284996 436152 285048
rect 2780 284928 2832 284980
rect 252836 284928 252888 284980
rect 345480 284928 345532 284980
rect 575480 284928 575532 284980
rect 153200 283840 153252 283892
rect 277860 283840 277912 283892
rect 314936 283840 314988 283892
rect 390560 283840 390612 283892
rect 217600 283772 217652 283824
rect 350632 283772 350684 283824
rect 138020 283704 138072 283756
rect 275008 283704 275060 283756
rect 324780 283704 324832 283756
rect 442264 283704 442316 283756
rect 58624 283636 58676 283688
rect 261300 283636 261352 283688
rect 337108 283636 337160 283688
rect 521660 283636 521712 283688
rect 20720 283568 20772 283620
rect 255596 283568 255648 283620
rect 339776 283568 339828 283620
rect 536104 283568 536156 283620
rect 313464 282412 313516 282464
rect 371884 282412 371936 282464
rect 157340 282344 157392 282396
rect 277768 282344 277820 282396
rect 319168 282344 319220 282396
rect 414664 282344 414716 282396
rect 131120 282276 131172 282328
rect 273536 282276 273588 282328
rect 327356 282276 327408 282328
rect 458824 282276 458876 282328
rect 107660 282208 107712 282260
rect 269580 282208 269632 282260
rect 328828 282208 328880 282260
rect 471244 282208 471296 282260
rect 39304 282140 39356 282192
rect 258264 282140 258316 282192
rect 342536 282140 342588 282192
rect 556252 282140 556304 282192
rect 320548 280984 320600 281036
rect 417424 280984 417476 281036
rect 142160 280916 142212 280968
rect 274916 280916 274968 280968
rect 326068 280916 326120 280968
rect 445024 280916 445076 280968
rect 126980 280848 127032 280900
rect 272248 280848 272300 280900
rect 330024 280848 330076 280900
rect 481732 280848 481784 280900
rect 26240 280780 26292 280832
rect 257068 280780 257120 280832
rect 345388 280780 345440 280832
rect 571984 280780 572036 280832
rect 319076 279624 319128 279676
rect 409880 279624 409932 279676
rect 165620 279556 165672 279608
rect 279056 279556 279108 279608
rect 320456 279556 320508 279608
rect 423680 279556 423732 279608
rect 57244 279488 57296 279540
rect 261208 279488 261260 279540
rect 332968 279488 333020 279540
rect 493324 279488 493376 279540
rect 21364 279420 21416 279472
rect 255504 279420 255556 279472
rect 338396 279420 338448 279472
rect 531320 279420 531372 279472
rect 188344 278264 188396 278316
rect 281816 278264 281868 278316
rect 147680 278196 147732 278248
rect 276296 278196 276348 278248
rect 321836 278196 321888 278248
rect 428464 278196 428516 278248
rect 98000 278128 98052 278180
rect 268200 278128 268252 278180
rect 323216 278128 323268 278180
rect 441620 278128 441672 278180
rect 71780 278060 71832 278112
rect 264152 278060 264204 278112
rect 335636 278060 335688 278112
rect 511264 278060 511316 278112
rect 42800 277992 42852 278044
rect 253388 277992 253440 278044
rect 345296 277992 345348 278044
rect 578240 277992 578292 278044
rect 196624 276904 196676 276956
rect 281724 276904 281776 276956
rect 136640 276836 136692 276888
rect 274824 276836 274876 276888
rect 317604 276836 317656 276888
rect 407212 276836 407264 276888
rect 102140 276768 102192 276820
rect 269488 276768 269540 276820
rect 323124 276768 323176 276820
rect 439504 276768 439556 276820
rect 78680 276700 78732 276752
rect 265440 276700 265492 276752
rect 337016 276700 337068 276752
rect 522304 276700 522356 276752
rect 35900 276632 35952 276684
rect 258172 276632 258224 276684
rect 342444 276632 342496 276684
rect 560300 276632 560352 276684
rect 193312 275544 193364 275596
rect 283196 275544 283248 275596
rect 127072 275476 127124 275528
rect 273444 275476 273496 275528
rect 317512 275476 317564 275528
rect 405004 275476 405056 275528
rect 111800 275408 111852 275460
rect 270960 275408 271012 275460
rect 324688 275408 324740 275460
rect 448612 275408 448664 275460
rect 93860 275340 93912 275392
rect 268108 275340 268160 275392
rect 325976 275340 326028 275392
rect 454684 275340 454736 275392
rect 11060 275272 11112 275324
rect 247684 275272 247736 275324
rect 336924 275272 336976 275324
rect 525064 275272 525116 275324
rect 324596 274184 324648 274236
rect 446404 274184 446456 274236
rect 197360 274116 197412 274168
rect 284484 274116 284536 274168
rect 324504 274116 324556 274168
rect 449900 274116 449952 274168
rect 162860 274048 162912 274100
rect 278964 274048 279016 274100
rect 325884 274048 325936 274100
rect 459560 274048 459612 274100
rect 120080 273980 120132 274032
rect 272156 273980 272208 274032
rect 338304 273980 338356 274032
rect 531412 273980 531464 274032
rect 93952 273912 94004 273964
rect 268016 273912 268068 273964
rect 362224 273912 362276 273964
rect 580172 273912 580224 273964
rect 201592 272756 201644 272808
rect 284392 272756 284444 272808
rect 187700 272688 187752 272740
rect 283104 272688 283156 272740
rect 102232 272620 102284 272672
rect 269396 272620 269448 272672
rect 80060 272552 80112 272604
rect 265348 272552 265400 272604
rect 328736 272552 328788 272604
rect 475384 272552 475436 272604
rect 57980 272484 58032 272536
rect 261116 272484 261168 272536
rect 339684 272484 339736 272536
rect 540244 272484 540296 272536
rect 211804 271396 211856 271448
rect 285864 271396 285916 271448
rect 180800 271328 180852 271380
rect 282092 271328 282144 271380
rect 99380 271260 99432 271312
rect 260196 271260 260248 271312
rect 314844 271260 314896 271312
rect 386420 271260 386472 271312
rect 77300 271192 77352 271244
rect 265256 271192 265308 271244
rect 329932 271192 329984 271244
rect 484400 271192 484452 271244
rect 53840 271124 53892 271176
rect 261024 271124 261076 271176
rect 339592 271124 339644 271176
rect 545120 271124 545172 271176
rect 167000 269968 167052 270020
rect 278872 269968 278924 270020
rect 314752 269968 314804 270020
rect 390652 269968 390704 270020
rect 92480 269900 92532 269952
rect 266820 269900 266872 269952
rect 331404 269900 331456 269952
rect 486424 269900 486476 269952
rect 75920 269832 75972 269884
rect 264060 269832 264112 269884
rect 335544 269832 335596 269884
rect 517520 269832 517572 269884
rect 14464 269764 14516 269816
rect 254032 269764 254084 269816
rect 341064 269764 341116 269816
rect 552020 269764 552072 269816
rect 144920 268472 144972 268524
rect 276204 268472 276256 268524
rect 74540 268404 74592 268456
rect 263968 268404 264020 268456
rect 327264 268404 327316 268456
rect 467840 268404 467892 268456
rect 7564 268336 7616 268388
rect 252744 268336 252796 268388
rect 328644 268336 328696 268388
rect 473452 268336 473504 268388
rect 2964 267656 3016 267708
rect 225604 267656 225656 267708
rect 218612 267180 218664 267232
rect 347872 267180 347924 267232
rect 332876 267112 332928 267164
rect 495440 267112 495492 267164
rect 67640 267044 67692 267096
rect 263876 267044 263928 267096
rect 340972 267044 341024 267096
rect 553400 267044 553452 267096
rect 48320 266976 48372 267028
rect 259644 266976 259696 267028
rect 344008 266976 344060 267028
rect 565820 266976 565872 267028
rect 191840 265888 191892 265940
rect 283472 265888 283524 265940
rect 133880 265820 133932 265872
rect 273352 265820 273404 265872
rect 115940 265752 115992 265804
rect 270776 265752 270828 265804
rect 331312 265752 331364 265804
rect 491300 265752 491352 265804
rect 114560 265684 114612 265736
rect 270868 265684 270920 265736
rect 338212 265684 338264 265736
rect 535460 265684 535512 265736
rect 31760 265616 31812 265668
rect 250536 265616 250588 265668
rect 342352 265616 342404 265668
rect 560944 265616 560996 265668
rect 143632 264392 143684 264444
rect 275284 264392 275336 264444
rect 113180 264324 113232 264376
rect 270684 264324 270736 264376
rect 313280 264324 313332 264376
rect 382372 264324 382424 264376
rect 96620 264256 96672 264308
rect 267924 264256 267976 264308
rect 320364 264256 320416 264308
rect 420920 264256 420972 264308
rect 84200 264188 84252 264240
rect 265164 264188 265216 264240
rect 340880 264188 340932 264240
rect 549260 264188 549312 264240
rect 314660 262964 314712 263016
rect 389180 262964 389232 263016
rect 154580 262896 154632 262948
rect 277676 262896 277728 262948
rect 323032 262896 323084 262948
rect 434720 262896 434772 262948
rect 151912 262828 151964 262880
rect 276112 262828 276164 262880
rect 345204 262828 345256 262880
rect 574100 262828 574152 262880
rect 212540 261808 212592 261860
rect 287336 261808 287388 261860
rect 158720 261740 158772 261792
rect 277584 261740 277636 261792
rect 316592 261740 316644 261792
rect 393320 261740 393372 261792
rect 149060 261672 149112 261724
rect 276572 261672 276624 261724
rect 316500 261672 316552 261724
rect 397460 261672 397512 261724
rect 217784 261604 217836 261656
rect 345112 261604 345164 261656
rect 69020 261536 69072 261588
rect 263784 261536 263836 261588
rect 329840 261536 329892 261588
rect 485780 261536 485832 261588
rect 13820 261468 13872 261520
rect 254400 261468 254452 261520
rect 343916 261468 343968 261520
rect 569960 261468 570012 261520
rect 124220 260312 124272 260364
rect 251916 260312 251968 260364
rect 39396 260244 39448 260296
rect 256884 260244 256936 260296
rect 30380 260176 30432 260228
rect 256976 260176 257028 260228
rect 339500 260176 339552 260228
rect 542360 260176 542412 260228
rect 4160 260108 4212 260160
rect 246304 260108 246356 260160
rect 342260 260108 342312 260160
rect 558920 260108 558972 260160
rect 374644 259360 374696 259412
rect 580172 259360 580224 259412
rect 176660 258816 176712 258868
rect 267004 258816 267056 258868
rect 173900 258748 173952 258800
rect 280620 258748 280672 258800
rect 316408 258748 316460 258800
rect 398840 258748 398892 258800
rect 217508 258680 217560 258732
rect 346492 258680 346544 258732
rect 117320 257524 117372 257576
rect 260104 257524 260156 257576
rect 106280 257456 106332 257508
rect 261484 257456 261536 257508
rect 23480 257388 23532 257440
rect 251824 257388 251876 257440
rect 316316 257388 316368 257440
rect 391940 257388 391992 257440
rect 25596 257320 25648 257372
rect 255412 257320 255464 257372
rect 316224 257320 316276 257372
rect 396080 257320 396132 257372
rect 218428 256300 218480 256352
rect 287244 256300 287296 256352
rect 217232 256232 217284 256284
rect 350540 256232 350592 256284
rect 122840 256164 122892 256216
rect 271972 256164 272024 256216
rect 318984 256164 319036 256216
rect 413284 256164 413336 256216
rect 118700 256096 118752 256148
rect 272064 256096 272116 256148
rect 320272 256096 320324 256148
rect 425060 256096 425112 256148
rect 77392 256028 77444 256080
rect 265072 256028 265124 256080
rect 321744 256028 321796 256080
rect 431960 256028 432012 256080
rect 17960 255960 18012 256012
rect 255780 255960 255832 256012
rect 324412 255960 324464 256012
rect 445116 255960 445168 256012
rect 169760 254804 169812 254856
rect 280528 254804 280580 254856
rect 311992 254804 312044 254856
rect 372620 254804 372672 254856
rect 3332 254736 3384 254788
rect 8944 254736 8996 254788
rect 110420 254736 110472 254788
rect 269304 254736 269356 254788
rect 317420 254736 317472 254788
rect 404360 254736 404412 254788
rect 88340 254668 88392 254720
rect 253296 254668 253348 254720
rect 328552 254668 328604 254720
rect 474740 254668 474792 254720
rect 91100 254600 91152 254652
rect 266728 254600 266780 254652
rect 343732 254600 343784 254652
rect 564532 254600 564584 254652
rect 86960 254532 87012 254584
rect 266636 254532 266688 254584
rect 343824 254532 343876 254584
rect 567200 254532 567252 254584
rect 303988 253852 304040 253904
rect 364340 253852 364392 253904
rect 303896 253784 303948 253836
rect 365812 253784 365864 253836
rect 301044 253716 301096 253768
rect 367192 253716 367244 253768
rect 300952 253648 301004 253700
rect 368480 253648 368532 253700
rect 316040 253580 316092 253632
rect 394700 253580 394752 253632
rect 176752 253512 176804 253564
rect 280436 253512 280488 253564
rect 316132 253512 316184 253564
rect 398932 253512 398984 253564
rect 217140 253444 217192 253496
rect 348424 253444 348476 253496
rect 118792 253376 118844 253428
rect 271052 253376 271104 253428
rect 332692 253376 332744 253428
rect 496084 253376 496136 253428
rect 110512 253308 110564 253360
rect 270592 253308 270644 253360
rect 332784 253308 332836 253360
rect 499580 253308 499632 253360
rect 95240 253240 95292 253292
rect 267832 253240 267884 253292
rect 334624 253240 334676 253292
rect 506480 253240 506532 253292
rect 73160 253172 73212 253224
rect 263692 253172 263744 253224
rect 336832 253172 336884 253224
rect 528560 253172 528612 253224
rect 302516 253104 302568 253156
rect 360200 253104 360252 253156
rect 302608 253036 302660 253088
rect 358820 253036 358872 253088
rect 172520 252220 172572 252272
rect 280344 252220 280396 252272
rect 160192 252152 160244 252204
rect 277400 252152 277452 252204
rect 321652 252152 321704 252204
rect 427820 252152 427872 252204
rect 155960 252084 156012 252136
rect 277492 252084 277544 252136
rect 321560 252084 321612 252136
rect 432052 252084 432104 252136
rect 218520 252016 218572 252068
rect 347780 252016 347832 252068
rect 60740 251948 60792 252000
rect 253204 251948 253256 252000
rect 325792 251948 325844 252000
rect 454040 251948 454092 252000
rect 49700 251880 49752 251932
rect 259552 251880 259604 251932
rect 327172 251880 327224 251932
rect 466460 251880 466512 251932
rect 46204 251812 46256 251864
rect 260012 251812 260064 251864
rect 334532 251812 334584 251864
rect 509240 251812 509292 251864
rect 309600 251132 309652 251184
rect 365720 251132 365772 251184
rect 306748 251064 306800 251116
rect 363144 251064 363196 251116
rect 306840 250996 306892 251048
rect 363236 250996 363288 251048
rect 308220 250928 308272 250980
rect 365996 250928 366048 250980
rect 305460 250860 305512 250912
rect 363328 250860 363380 250912
rect 209872 250792 209924 250844
rect 286048 250792 286100 250844
rect 302424 250792 302476 250844
rect 360292 250792 360344 250844
rect 135352 250724 135404 250776
rect 273720 250724 273772 250776
rect 306932 250724 306984 250776
rect 365904 250724 365956 250776
rect 70400 250656 70452 250708
rect 264244 250656 264296 250708
rect 311900 250656 311952 250708
rect 374092 250656 374144 250708
rect 66260 250588 66312 250640
rect 262588 250588 262640 250640
rect 318892 250588 318944 250640
rect 416780 250588 416832 250640
rect 62120 250520 62172 250572
rect 262496 250520 262548 250572
rect 331220 250520 331272 250572
rect 492680 250520 492732 250572
rect 52552 250452 52604 250504
rect 260932 250452 260984 250504
rect 345020 250452 345072 250504
rect 576860 250452 576912 250504
rect 309508 250384 309560 250436
rect 361580 250384 361632 250436
rect 185032 249296 185084 249348
rect 282184 249296 282236 249348
rect 318800 249296 318852 249348
rect 414020 249296 414072 249348
rect 85580 249228 85632 249280
rect 266544 249228 266596 249280
rect 338764 249228 338816 249280
rect 458180 249228 458232 249280
rect 82820 249160 82872 249212
rect 264980 249160 265032 249212
rect 327080 249160 327132 249212
rect 460940 249160 460992 249212
rect 59360 249092 59412 249144
rect 262404 249092 262456 249144
rect 328460 249092 328512 249144
rect 477500 249092 477552 249144
rect 57336 249024 57388 249076
rect 261392 249024 261444 249076
rect 335452 249024 335504 249076
rect 520280 249024 520332 249076
rect 308128 248344 308180 248396
rect 364524 248344 364576 248396
rect 305368 248276 305420 248328
rect 362960 248276 363012 248328
rect 306656 248208 306708 248260
rect 364432 248208 364484 248260
rect 305092 248140 305144 248192
rect 363052 248140 363104 248192
rect 198740 248072 198792 248124
rect 284760 248072 284812 248124
rect 302332 248072 302384 248124
rect 362040 248072 362092 248124
rect 175280 248004 175332 248056
rect 280252 248004 280304 248056
rect 302240 248004 302292 248056
rect 371332 248004 371384 248056
rect 140780 247936 140832 247988
rect 275192 247936 275244 247988
rect 320180 247936 320232 247988
rect 423772 247936 423824 247988
rect 89720 247868 89772 247920
rect 266452 247868 266504 247920
rect 325700 247868 325752 247920
rect 455420 247868 455472 247920
rect 41420 247800 41472 247852
rect 258632 247800 258684 247852
rect 332600 247800 332652 247852
rect 502340 247800 502392 247852
rect 35164 247732 35216 247784
rect 256792 247732 256844 247784
rect 334440 247732 334492 247784
rect 512000 247732 512052 247784
rect 8944 247664 8996 247716
rect 252652 247664 252704 247716
rect 336740 247664 336792 247716
rect 524420 247664 524472 247716
rect 309416 247596 309468 247648
rect 364616 247596 364668 247648
rect 355692 247528 355744 247580
rect 369952 247528 370004 247580
rect 217324 246712 217376 246764
rect 346400 246712 346452 246764
rect 121460 246644 121512 246696
rect 272340 246644 272392 246696
rect 300860 246644 300912 246696
rect 366088 246644 366140 246696
rect 109040 246576 109092 246628
rect 269212 246576 269264 246628
rect 322940 246576 322992 246628
rect 438860 246576 438912 246628
rect 85672 246508 85724 246560
rect 266912 246508 266964 246560
rect 334348 246508 334400 246560
rect 505100 246508 505152 246560
rect 64880 246440 64932 246492
rect 262312 246440 262364 246492
rect 334256 246440 334308 246492
rect 507860 246440 507912 246492
rect 38660 246372 38712 246424
rect 250444 246372 250496 246424
rect 334164 246372 334216 246424
rect 510620 246372 510672 246424
rect 6920 246304 6972 246356
rect 252928 246304 252980 246356
rect 335360 246304 335412 246356
rect 516140 246304 516192 246356
rect 355600 245556 355652 245608
rect 369860 245556 369912 245608
rect 355508 245488 355560 245540
rect 372712 245488 372764 245540
rect 307852 245420 307904 245472
rect 361764 245420 361816 245472
rect 307944 245352 307996 245404
rect 361856 245352 361908 245404
rect 203616 245284 203668 245336
rect 283380 245284 283432 245336
rect 307760 245284 307812 245336
rect 361672 245284 361724 245336
rect 171232 245216 171284 245268
rect 280712 245216 280764 245268
rect 306380 245216 306432 245268
rect 361948 245216 362000 245268
rect 168472 245148 168524 245200
rect 279240 245148 279292 245200
rect 324320 245148 324372 245200
rect 445760 245148 445812 245200
rect 104900 245080 104952 245132
rect 269672 245080 269724 245132
rect 334072 245080 334124 245132
rect 503720 245080 503772 245132
rect 100760 245012 100812 245064
rect 268292 245012 268344 245064
rect 333980 245012 334032 245064
rect 506572 245012 506624 245064
rect 60832 244944 60884 244996
rect 262680 244944 262732 244996
rect 338120 244944 338172 244996
rect 534080 244944 534132 244996
rect 27712 244876 27764 244928
rect 257252 244876 257304 244928
rect 343640 244876 343692 244928
rect 571340 244876 571392 244928
rect 355324 244468 355376 244520
rect 363420 244468 363472 244520
rect 355416 244264 355468 244316
rect 363788 244264 363840 244316
rect 303620 243856 303672 243908
rect 364708 243856 364760 243908
rect 299664 243788 299716 243840
rect 362224 243788 362276 243840
rect 299756 243720 299808 243772
rect 362408 243720 362460 243772
rect 298192 243652 298244 243704
rect 361028 243652 361080 243704
rect 219348 243584 219400 243636
rect 297180 243584 297232 243636
rect 299480 243584 299532 243636
rect 366548 243584 366600 243636
rect 217416 243516 217468 243568
rect 297272 243516 297324 243568
rect 299572 243516 299624 243568
rect 369308 243516 369360 243568
rect 3332 215228 3384 215280
rect 215944 215228 215996 215280
rect 214380 213868 214432 213920
rect 215944 213868 215996 213920
rect 373356 206932 373408 206984
rect 579620 206932 579672 206984
rect 3056 202784 3108 202836
rect 196716 202784 196768 202836
rect 215760 195372 215812 195424
rect 217692 195372 217744 195424
rect 577596 193128 577648 193180
rect 580816 193128 580868 193180
rect 371976 166948 372028 167000
rect 580172 166948 580224 167000
rect 358360 160080 358412 160132
rect 363788 160080 363840 160132
rect 322940 159604 322992 159656
rect 358176 159604 358228 159656
rect 318708 159536 318760 159588
rect 358084 159536 358136 159588
rect 213644 159468 213696 159520
rect 256700 159468 256752 159520
rect 314660 159468 314712 159520
rect 357808 159468 357860 159520
rect 211712 159400 211764 159452
rect 259460 159400 259512 159452
rect 310428 159400 310480 159452
rect 357992 159400 358044 159452
rect 215852 159332 215904 159384
rect 263692 159332 263744 159384
rect 305000 159332 305052 159384
rect 356704 159332 356756 159384
rect 300952 159196 301004 159248
rect 357900 159196 357952 159248
rect 295892 159128 295944 159180
rect 370688 159128 370740 159180
rect 288348 159060 288400 159112
rect 365076 159060 365128 159112
rect 279240 158992 279292 159044
rect 360844 158992 360896 159044
rect 278136 158924 278188 158976
rect 360752 158924 360804 158976
rect 277032 158856 277084 158908
rect 360660 158856 360712 158908
rect 275836 158788 275888 158840
rect 359372 158788 359424 158840
rect 211896 158720 211948 158772
rect 239588 158720 239640 158772
rect 274456 158720 274508 158772
rect 359464 158720 359516 158772
rect 213276 158652 213328 158704
rect 238116 158652 238168 158704
rect 298560 158652 298612 158704
rect 305000 158652 305052 158704
rect 306104 158652 306156 158704
rect 314660 158652 314712 158704
rect 212080 158584 212132 158636
rect 230480 158584 230532 158636
rect 308772 158584 308824 158636
rect 318708 158584 318760 158636
rect 214840 158516 214892 158568
rect 236000 158516 236052 158568
rect 262864 158516 262916 158568
rect 367744 158516 367796 158568
rect 213368 158448 213420 158500
rect 234712 158448 234764 158500
rect 259552 158448 259604 158500
rect 364800 158448 364852 158500
rect 219072 158380 219124 158432
rect 242992 158380 243044 158432
rect 263600 158380 263652 158432
rect 362316 158380 362368 158432
rect 214564 158312 214616 158364
rect 242900 158312 242952 158364
rect 268752 158312 268804 158364
rect 357716 158312 357768 158364
rect 214932 158244 214984 158296
rect 245660 158244 245712 158296
rect 269856 158244 269908 158296
rect 357532 158244 357584 158296
rect 216220 158176 216272 158228
rect 247040 158176 247092 158228
rect 271144 158176 271196 158228
rect 357624 158176 357676 158228
rect 217968 158108 218020 158160
rect 251180 158108 251232 158160
rect 303528 158108 303580 158160
rect 310428 158108 310480 158160
rect 321008 158108 321060 158160
rect 360568 158108 360620 158160
rect 219164 158040 219216 158092
rect 252560 158040 252612 158092
rect 313464 158040 313516 158092
rect 359096 158040 359148 158092
rect 216312 157972 216364 158024
rect 249800 157972 249852 158024
rect 315856 157972 315908 158024
rect 359280 157972 359332 158024
rect 216128 157904 216180 157956
rect 233240 157904 233292 157956
rect 318616 157904 318668 157956
rect 359188 157904 359240 157956
rect 218980 157836 219032 157888
rect 234620 157836 234672 157888
rect 272248 157836 272300 157888
rect 322940 157836 322992 157888
rect 323400 157836 323452 157888
rect 360384 157836 360436 157888
rect 214656 157768 214708 157820
rect 229100 157768 229152 157820
rect 325976 157768 326028 157820
rect 360476 157768 360528 157820
rect 240692 157700 240744 157752
rect 372988 157700 373040 157752
rect 261484 157632 261536 157684
rect 366456 157632 366508 157684
rect 248328 157292 248380 157344
rect 370412 157292 370464 157344
rect 252376 157224 252428 157276
rect 369124 157224 369176 157276
rect 250444 157156 250496 157208
rect 366364 157156 366416 157208
rect 254952 157088 255004 157140
rect 363512 157088 363564 157140
rect 257252 157020 257304 157072
rect 366180 157020 366232 157072
rect 259092 156952 259144 157004
rect 366272 156952 366324 157004
rect 255872 156884 255924 156936
rect 360936 156884 360988 156936
rect 271052 156816 271104 156868
rect 374184 156816 374236 156868
rect 276112 156748 276164 156800
rect 369032 156748 369084 156800
rect 281356 156680 281408 156732
rect 371700 156680 371752 156732
rect 286324 156612 286376 156664
rect 371792 156612 371844 156664
rect 274456 156544 274508 156596
rect 358912 156544 358964 156596
rect 293684 156476 293736 156528
rect 371608 156476 371660 156528
rect 311072 156408 311124 156460
rect 359004 156408 359056 156460
rect 248696 155864 248748 155916
rect 368848 155864 368900 155916
rect 211988 155796 212040 155848
rect 237380 155796 237432 155848
rect 252284 155796 252336 155848
rect 370228 155796 370280 155848
rect 213552 155728 213604 155780
rect 241520 155728 241572 155780
rect 253572 155728 253624 155780
rect 363604 155728 363656 155780
rect 216036 155660 216088 155712
rect 248420 155660 248472 155712
rect 260656 155660 260708 155712
rect 367284 155660 367336 155712
rect 213460 155592 213512 155644
rect 253940 155592 253992 155644
rect 261760 155592 261812 155644
rect 367468 155592 367520 155644
rect 210700 155524 210752 155576
rect 267832 155524 267884 155576
rect 268936 155524 268988 155576
rect 372804 155524 372856 155576
rect 210884 155456 210936 155508
rect 255320 155456 255372 155508
rect 264520 155456 264572 155508
rect 367560 155456 367612 155508
rect 219256 155388 219308 155440
rect 264980 155388 265032 155440
rect 266912 155388 266964 155440
rect 370044 155388 370096 155440
rect 214472 155320 214524 155372
rect 260840 155320 260892 155372
rect 265992 155320 266044 155372
rect 367376 155320 367428 155372
rect 218796 155252 218848 155304
rect 266360 155252 266412 155304
rect 267648 155252 267700 155304
rect 368572 155252 368624 155304
rect 212172 155184 212224 155236
rect 273260 155184 273312 155236
rect 274548 155184 274600 155236
rect 368756 155184 368808 155236
rect 217692 155116 217744 155168
rect 277400 155116 277452 155168
rect 278688 155116 278740 155168
rect 368940 155116 368992 155168
rect 217416 155048 217468 155100
rect 278780 155048 278832 155100
rect 283932 155048 283984 155100
rect 371516 155048 371568 155100
rect 217876 154980 217928 155032
rect 274640 154980 274692 155032
rect 291016 154980 291068 155032
rect 372068 154980 372120 155032
rect 253664 154504 253716 154556
rect 371424 154504 371476 154556
rect 256240 154436 256292 154488
rect 359556 154436 359608 154488
rect 345756 154232 345808 154284
rect 366548 154232 366600 154284
rect 295340 154164 295392 154216
rect 362224 154164 362276 154216
rect 299572 154096 299624 154148
rect 370504 154096 370556 154148
rect 288440 154028 288492 154080
rect 361028 154028 361080 154080
rect 298100 153960 298152 154012
rect 372896 153960 372948 154012
rect 293960 153892 294012 153944
rect 369308 153892 369360 153944
rect 285680 153824 285732 153876
rect 367836 153824 367888 153876
rect 3516 150356 3568 150408
rect 199384 150356 199436 150408
rect 3516 137912 3568 137964
rect 203524 137912 203576 137964
rect 3424 97928 3476 97980
rect 198004 97928 198056 97980
rect 3148 85484 3200 85536
rect 206284 85484 206336 85536
rect 3424 71680 3476 71732
rect 207664 71680 207716 71732
rect 378784 60664 378836 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 25504 59304 25556 59356
rect 3424 45500 3476 45552
rect 82084 45500 82136 45552
rect 3516 33056 3568 33108
rect 88984 33056 89036 33108
rect 3424 20612 3476 20664
rect 192576 20612 192628 20664
rect 160100 11704 160152 11756
rect 161296 11704 161348 11756
rect 176660 11704 176712 11756
rect 177856 11704 177908 11756
rect 184940 11704 184992 11756
rect 186136 11704 186188 11756
rect 201500 11704 201552 11756
rect 202696 11704 202748 11756
rect 234620 11704 234672 11756
rect 235816 11704 235868 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 319720 9392 319772 9444
rect 365812 9392 365864 9444
rect 316224 9324 316276 9376
rect 364708 9324 364760 9376
rect 322112 9256 322164 9308
rect 372712 9256 372764 9308
rect 303160 9188 303212 9240
rect 358268 9188 358320 9240
rect 306748 9120 306800 9172
rect 368480 9120 368532 9172
rect 309048 9052 309100 9104
rect 369952 9052 370004 9104
rect 305552 8984 305604 9036
rect 367192 8984 367244 9036
rect 304356 8916 304408 8968
rect 366088 8916 366140 8968
rect 3424 6808 3476 6860
rect 200764 6808 200816 6860
rect 337476 6808 337528 6860
rect 363144 6808 363196 6860
rect 333888 6740 333940 6792
rect 363236 6740 363288 6792
rect 577504 6740 577556 6792
rect 580264 6740 580316 6792
rect 330392 6672 330444 6724
rect 363328 6672 363380 6724
rect 318524 6604 318576 6656
rect 364340 6604 364392 6656
rect 313832 6536 313884 6588
rect 360292 6536 360344 6588
rect 317328 6468 317380 6520
rect 363420 6468 363472 6520
rect 315028 6400 315080 6452
rect 362040 6400 362092 6452
rect 312636 6332 312688 6384
rect 360200 6332 360252 6384
rect 311440 6264 311492 6316
rect 358820 6264 358872 6316
rect 307944 6196 307996 6248
rect 369860 6196 369912 6248
rect 310244 6128 310296 6180
rect 371332 6128 371384 6180
rect 340972 6060 341024 6112
rect 365904 6060 365956 6112
rect 344560 5992 344612 6044
rect 365996 5992 366048 6044
rect 350448 5924 350500 5976
rect 364616 5924 364668 5976
rect 6460 4088 6512 4140
rect 8944 4088 8996 4140
rect 44272 4088 44324 4140
rect 46204 4088 46256 4140
rect 180248 4088 180300 4140
rect 181444 4088 181496 4140
rect 216404 4088 216456 4140
rect 240508 4088 240560 4140
rect 336280 4088 336332 4140
rect 364432 4088 364484 4140
rect 428556 4088 428608 4140
rect 434444 4088 434496 4140
rect 460204 4088 460256 4140
rect 462780 4088 462832 4140
rect 468484 4088 468536 4140
rect 471060 4088 471112 4140
rect 478236 4088 478288 4140
rect 482836 4088 482888 4140
rect 536196 4088 536248 4140
rect 538404 4088 538456 4140
rect 51356 4020 51408 4072
rect 57244 4020 57296 4072
rect 212356 4020 212408 4072
rect 245200 4020 245252 4072
rect 332692 4020 332744 4072
rect 363052 4020 363104 4072
rect 213736 3952 213788 4004
rect 258264 3952 258316 4004
rect 329196 3952 329248 4004
rect 362960 3952 363012 4004
rect 213828 3884 213880 3936
rect 260656 3884 260708 3936
rect 301964 3884 302016 3936
rect 352564 3884 352616 3936
rect 4068 3816 4120 3868
rect 7564 3816 7616 3868
rect 215024 3816 215076 3868
rect 262956 3816 263008 3868
rect 291384 3816 291436 3868
rect 345756 3816 345808 3868
rect 354036 3816 354088 3868
rect 363788 3816 363840 3868
rect 440884 3816 440936 3868
rect 443828 3816 443880 3868
rect 516784 3816 516836 3868
rect 519544 3816 519596 3868
rect 566464 3816 566516 3868
rect 569132 3816 569184 3868
rect 211068 3748 211120 3800
rect 268844 3748 268896 3800
rect 292580 3748 292632 3800
rect 348424 3748 348476 3800
rect 349252 3748 349304 3800
rect 361856 3748 361908 3800
rect 30104 3680 30156 3732
rect 39396 3680 39448 3732
rect 69112 3680 69164 3732
rect 71044 3680 71096 3732
rect 135260 3680 135312 3732
rect 136456 3680 136508 3732
rect 212264 3680 212316 3732
rect 272432 3680 272484 3732
rect 299572 3680 299624 3732
rect 300768 3680 300820 3732
rect 301780 3680 301832 3732
rect 353944 3680 353996 3732
rect 445024 3680 445076 3732
rect 458088 3680 458140 3732
rect 489184 3680 489236 3732
rect 491116 3680 491168 3732
rect 1676 3612 1728 3664
rect 32404 3612 32456 3664
rect 37188 3612 37240 3664
rect 43444 3612 43496 3664
rect 46664 3612 46716 3664
rect 170496 3612 170548 3664
rect 187332 3612 187384 3664
rect 196624 3612 196676 3664
rect 215944 3612 215996 3664
rect 276020 3612 276072 3664
rect 285404 3612 285456 3664
rect 345664 3612 345716 3664
rect 346952 3612 347004 3664
rect 363880 3612 363932 3664
rect 427084 3612 427136 3664
rect 440332 3612 440384 3664
rect 476764 3612 476816 3664
rect 20628 3544 20680 3596
rect 21364 3544 21416 3596
rect 25320 3544 25372 3596
rect 171784 3544 171836 3596
rect 183744 3544 183796 3596
rect 188344 3544 188396 3596
rect 195612 3544 195664 3596
rect 203616 3544 203668 3596
rect 216588 3544 216640 3596
rect 284300 3544 284352 3596
rect 287796 3544 287848 3596
rect 354128 3544 354180 3596
rect 355232 3544 355284 3596
rect 365720 3544 365772 3596
rect 377404 3544 377456 3596
rect 411904 3544 411956 3596
rect 421564 3544 421616 3596
rect 427268 3544 427320 3596
rect 442264 3544 442316 3596
rect 445024 3544 445076 3596
rect 458824 3544 458876 3596
rect 465172 3544 465224 3596
rect 467104 3544 467156 3596
rect 469864 3544 469916 3596
rect 12348 3476 12400 3528
rect 13084 3476 13136 3528
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 15936 3476 15988 3528
rect 170404 3476 170456 3528
rect 219348 3476 219400 3528
rect 280712 3476 280764 3528
rect 281908 3476 281960 3528
rect 357440 3476 357492 3528
rect 374092 3476 374144 3528
rect 375288 3476 375340 3528
rect 381544 3476 381596 3528
rect 572 3408 624 3460
rect 171140 3408 171192 3460
rect 190828 3408 190880 3460
rect 199476 3408 199528 3460
rect 215116 3408 215168 3460
rect 277124 3408 277176 3460
rect 283104 3408 283156 3460
rect 367100 3408 367152 3460
rect 373264 3408 373316 3460
rect 384764 3408 384816 3460
rect 387064 3408 387116 3460
rect 388260 3408 388312 3460
rect 390560 3408 390612 3460
rect 391848 3408 391900 3460
rect 33600 3340 33652 3392
rect 35164 3340 35216 3392
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 56048 3340 56100 3392
rect 57336 3340 57388 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 212448 3340 212500 3392
rect 227536 3340 227588 3392
rect 297272 3340 297324 3392
rect 301780 3340 301832 3392
rect 338672 3340 338724 3392
rect 361948 3340 362000 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 388444 3340 388496 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 57244 3272 57296 3324
rect 58624 3272 58676 3324
rect 208584 3272 208636 3324
rect 211804 3272 211856 3324
rect 215208 3272 215260 3324
rect 222752 3272 222804 3324
rect 343364 3272 343416 3324
rect 364524 3272 364576 3324
rect 414664 3408 414716 3460
rect 416688 3408 416740 3460
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 431960 3476 432012 3528
rect 433248 3476 433300 3528
rect 439504 3476 439556 3528
rect 441528 3476 441580 3528
rect 448520 3476 448572 3528
rect 449808 3476 449860 3528
rect 454684 3476 454736 3528
rect 456892 3476 456944 3528
rect 462964 3476 463016 3528
rect 471244 3476 471296 3528
rect 473452 3476 473504 3528
rect 475384 3544 475436 3596
rect 476948 3544 477000 3596
rect 484032 3544 484084 3596
rect 500224 3544 500276 3596
rect 501788 3544 501840 3596
rect 511264 3544 511316 3596
rect 513564 3544 513616 3596
rect 525064 3544 525116 3596
rect 527732 3544 527784 3596
rect 479340 3476 479392 3528
rect 496084 3476 496136 3528
rect 497096 3476 497148 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 520924 3476 520976 3528
rect 523040 3476 523092 3528
rect 527824 3476 527876 3528
rect 533712 3544 533764 3596
rect 549904 3544 549956 3596
rect 551468 3544 551520 3596
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 545764 3476 545816 3528
rect 546684 3476 546736 3528
rect 570604 3476 570656 3528
rect 572720 3476 572772 3528
rect 429660 3340 429712 3392
rect 581000 3408 581052 3460
rect 493324 3340 493376 3392
rect 499396 3340 499448 3392
rect 543004 3340 543056 3392
rect 549076 3340 549128 3392
rect 446404 3272 446456 3324
rect 452108 3272 452160 3324
rect 509884 3272 509936 3324
rect 514760 3272 514812 3324
rect 216496 3204 216548 3256
rect 226340 3204 226392 3256
rect 342168 3204 342220 3256
rect 361672 3204 361724 3256
rect 405004 3204 405056 3256
rect 408408 3204 408460 3256
rect 554044 3204 554096 3256
rect 557356 3204 557408 3256
rect 345756 3136 345808 3188
rect 361764 3136 361816 3188
rect 371884 3136 371936 3188
rect 376484 3136 376536 3188
rect 435364 3136 435416 3188
rect 437940 3136 437992 3188
rect 485044 3136 485096 3188
rect 487620 3136 487672 3188
rect 534724 3136 534776 3188
rect 537208 3136 537260 3188
rect 560944 3136 560996 3188
rect 563244 3136 563296 3188
rect 352840 3068 352892 3120
rect 362500 3068 362552 3120
rect 445116 3068 445168 3120
rect 447416 3068 447468 3120
rect 19432 3000 19484 3052
rect 25596 3000 25648 3052
rect 413284 3000 413336 3052
rect 415492 3000 415544 3052
rect 417516 3000 417568 3052
rect 420184 3000 420236 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 486516 3000 486568 3052
rect 488816 3000 488868 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 522304 3000 522356 3052
rect 524236 3000 524288 3052
rect 538864 3000 538916 3052
rect 540796 3000 540848 3052
rect 563704 3000 563756 3052
rect 565636 3000 565688 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 396724 2932 396776 2984
rect 402520 2932 402572 2984
rect 540244 2932 540296 2984
rect 541992 2932 542044 2984
rect 552756 2932 552808 2984
rect 554964 2932 555016 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 21364 683188 21416 683194
rect 21364 683130 21416 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3422 606112 3478 606121
rect 3422 606047 3424 606056
rect 3476 606047 3478 606056
rect 3424 606018 3476 606024
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553722 3464 553823
rect 3424 553716 3476 553722
rect 3424 553658 3476 553664
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 4816 467158 4844 632062
rect 7564 606076 7616 606082
rect 7564 606018 7616 606024
rect 7576 478174 7604 606018
rect 8944 553716 8996 553722
rect 8944 553658 8996 553664
rect 7564 478168 7616 478174
rect 7564 478110 7616 478116
rect 8956 472666 8984 553658
rect 13084 501016 13136 501022
rect 13084 500958 13136 500964
rect 8944 472660 8996 472666
rect 8944 472602 8996 472608
rect 13096 471306 13124 500958
rect 13084 471300 13136 471306
rect 13084 471242 13136 471248
rect 4804 467152 4856 467158
rect 4804 467094 4856 467100
rect 21376 465730 21404 683130
rect 21364 465724 21416 465730
rect 21364 465666 21416 465672
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 25516 450566 25544 699654
rect 28264 656940 28316 656946
rect 28264 656882 28316 656888
rect 28276 457502 28304 656882
rect 35164 527196 35216 527202
rect 35164 527138 35216 527144
rect 35176 469878 35204 527138
rect 35164 469872 35216 469878
rect 35164 469814 35216 469820
rect 28264 457496 28316 457502
rect 28264 457438 28316 457444
rect 40052 454714 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 57244 579692 57296 579698
rect 57244 579634 57296 579640
rect 57256 468518 57284 579634
rect 57244 468512 57296 468518
rect 57244 468454 57296 468460
rect 71792 461650 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 71780 461644 71832 461650
rect 71780 461586 71832 461592
rect 88352 456074 88380 702406
rect 98644 700324 98696 700330
rect 98644 700266 98696 700272
rect 98656 460222 98684 700266
rect 105464 699786 105492 703520
rect 105452 699780 105504 699786
rect 105452 699722 105504 699728
rect 108304 699780 108356 699786
rect 108304 699722 108356 699728
rect 98644 460216 98696 460222
rect 98644 460158 98696 460164
rect 88340 456068 88392 456074
rect 88340 456010 88392 456016
rect 40040 454708 40092 454714
rect 40040 454650 40092 454656
rect 108316 451926 108344 699722
rect 137848 699718 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 140044 699712 140096 699718
rect 140044 699654 140096 699660
rect 140056 458930 140084 699654
rect 153212 474026 153240 702406
rect 153200 474020 153252 474026
rect 153200 473962 153252 473968
rect 140044 458924 140096 458930
rect 140044 458866 140096 458872
rect 169772 453422 169800 702406
rect 201512 456278 201540 702986
rect 217968 700392 218020 700398
rect 217968 700334 218020 700340
rect 217876 700324 217928 700330
rect 217876 700266 217928 700272
rect 215944 670744 215996 670750
rect 215944 670686 215996 670692
rect 214564 618316 214616 618322
rect 214564 618258 214616 618264
rect 211804 565888 211856 565894
rect 211804 565830 211856 565836
rect 210424 514820 210476 514826
rect 210424 514762 210476 514768
rect 201500 456272 201552 456278
rect 201500 456214 201552 456220
rect 169760 453416 169812 453422
rect 169760 453358 169812 453364
rect 210436 452130 210464 514762
rect 211816 461854 211844 565830
rect 211804 461848 211856 461854
rect 211804 461790 211856 461796
rect 214576 453626 214604 618258
rect 215956 459066 215984 670686
rect 217784 565140 217836 565146
rect 217784 565082 217836 565088
rect 217598 516896 217654 516905
rect 217598 516831 217654 516840
rect 217506 513768 217562 513777
rect 217506 513703 217562 513712
rect 217414 489968 217470 489977
rect 217414 489903 217470 489912
rect 217322 488064 217378 488073
rect 217322 487999 217378 488008
rect 215944 459060 215996 459066
rect 215944 459002 215996 459008
rect 214564 453620 214616 453626
rect 214564 453562 214616 453568
rect 210424 452124 210476 452130
rect 210424 452066 210476 452072
rect 108304 451920 108356 451926
rect 108304 451862 108356 451868
rect 25504 450560 25556 450566
rect 25504 450502 25556 450508
rect 4066 449576 4122 449585
rect 4122 449534 4200 449562
rect 4066 449511 4122 449520
rect 4172 446486 4200 449534
rect 217336 447846 217364 487999
rect 217428 478378 217456 489903
rect 217416 478372 217468 478378
rect 217416 478314 217468 478320
rect 217520 472802 217548 513703
rect 217508 472796 217560 472802
rect 217508 472738 217560 472744
rect 217612 471374 217640 516831
rect 217690 515944 217746 515953
rect 217690 515879 217746 515888
rect 217600 471368 217652 471374
rect 217600 471310 217652 471316
rect 217704 467294 217732 515879
rect 217692 467288 217744 467294
rect 217692 467230 217744 467236
rect 217324 447840 217376 447846
rect 217324 447782 217376 447788
rect 4160 446480 4212 446486
rect 4160 446422 4212 446428
rect 203524 446208 203576 446214
rect 203524 446150 203576 446156
rect 199384 446140 199436 446146
rect 199384 446082 199436 446088
rect 82084 445800 82136 445806
rect 82084 445742 82136 445748
rect 7564 444508 7616 444514
rect 7564 444450 7616 444456
rect 3516 442604 3568 442610
rect 3516 442546 3568 442552
rect 3424 440904 3476 440910
rect 3424 440846 3476 440852
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2780 284980 2832 284986
rect 2780 284922 2832 284928
rect 2792 16574 2820 284922
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3332 254788 3384 254794
rect 3332 254730 3384 254736
rect 3344 254153 3372 254730
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 110673 3464 440846
rect 3528 241097 3556 442546
rect 3608 442536 3660 442542
rect 3608 442478 3660 442484
rect 3620 345409 3648 442478
rect 7576 423638 7604 444450
rect 8944 441720 8996 441726
rect 8944 441662 8996 441668
rect 7564 423632 7616 423638
rect 7564 423574 7616 423580
rect 3700 376032 3752 376038
rect 3700 375974 3752 375980
rect 3712 358465 3740 375974
rect 3698 358456 3754 358465
rect 3698 358391 3754 358400
rect 3606 345400 3662 345409
rect 3606 345335 3662 345344
rect 8300 286340 8352 286346
rect 8300 286282 8352 286288
rect 7564 268388 7616 268394
rect 7564 268330 7616 268336
rect 4160 260160 4212 260166
rect 4160 260102 4212 260108
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 260102
rect 6920 246356 6972 246362
rect 6920 246298 6972 246304
rect 6932 16574 6960 246298
rect 2792 16546 2912 16574
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3606
rect 2884 480 2912 16546
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 3868 4120 3874
rect 4068 3810 4120 3816
rect 4080 480 4108 3810
rect 5276 480 5304 16546
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6472 480 6500 4082
rect 7484 3482 7512 16546
rect 7576 3874 7604 268330
rect 8312 16574 8340 286282
rect 8956 254794 8984 441662
rect 25504 440360 25556 440366
rect 25504 440302 25556 440308
rect 16580 295996 16632 296002
rect 16580 295938 16632 295944
rect 13084 290488 13136 290494
rect 13084 290430 13136 290436
rect 9680 289128 9732 289134
rect 9680 289070 9732 289076
rect 8944 254788 8996 254794
rect 8944 254730 8996 254736
rect 8944 247716 8996 247722
rect 8944 247658 8996 247664
rect 8312 16546 8800 16574
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 8956 4146 8984 247658
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 289070
rect 11060 275324 11112 275330
rect 11060 275266 11112 275272
rect 11072 16574 11100 275266
rect 11072 16546 11192 16574
rect 11164 480 11192 16546
rect 13096 3534 13124 290430
rect 14464 269816 14516 269822
rect 14464 269758 14516 269764
rect 13820 261520 13872 261526
rect 13820 261462 13872 261468
rect 13832 16574 13860 261462
rect 13832 16546 14320 16574
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 12360 480 12388 3470
rect 13556 480 13584 3470
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 3534 14504 269758
rect 16592 16574 16620 295938
rect 22100 291848 22152 291854
rect 22100 291790 22152 291796
rect 20720 283620 20772 283626
rect 20720 283562 20772 283568
rect 17960 256012 18012 256018
rect 17960 255954 18012 255960
rect 16592 16546 17080 16574
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 480 15976 3470
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 255954
rect 20732 16574 20760 283562
rect 21364 279472 21416 279478
rect 21364 279414 21416 279420
rect 20732 16546 21312 16574
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 20640 480 20668 3538
rect 21284 3482 21312 16546
rect 21376 3602 21404 279414
rect 22112 16574 22140 291790
rect 23480 257440 23532 257446
rect 23480 257382 23532 257388
rect 23492 16574 23520 257382
rect 25516 59362 25544 440302
rect 32404 373108 32456 373114
rect 32404 373050 32456 373056
rect 27620 287700 27672 287706
rect 27620 287642 27672 287648
rect 26240 280832 26292 280838
rect 26240 280774 26292 280780
rect 25596 257372 25648 257378
rect 25596 257314 25648 257320
rect 25504 59356 25556 59362
rect 25504 59298 25556 59304
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21284 3454 21864 3482
rect 21836 480 21864 3454
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 480 25360 3538
rect 25608 3058 25636 257314
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 280774
rect 27632 6914 27660 287642
rect 31760 265668 31812 265674
rect 31760 265610 31812 265616
rect 30380 260228 30432 260234
rect 30380 260170 30432 260176
rect 27712 244928 27764 244934
rect 27712 244870 27764 244876
rect 27724 16574 27752 244870
rect 30392 16574 30420 260170
rect 31772 16574 31800 265610
rect 27724 16546 28488 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30116 480 30144 3674
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3670 32444 373050
rect 34518 300112 34574 300121
rect 34518 300047 34574 300056
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 480 33640 3334
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 300047
rect 63500 296064 63552 296070
rect 63500 296006 63552 296012
rect 43444 294636 43496 294642
rect 43444 294578 43496 294584
rect 40040 285048 40092 285054
rect 40040 284990 40092 284996
rect 39304 282192 39356 282198
rect 39304 282134 39356 282140
rect 35900 276684 35952 276690
rect 35900 276626 35952 276632
rect 35164 247784 35216 247790
rect 35164 247726 35216 247732
rect 35176 3398 35204 247726
rect 35912 16574 35940 276626
rect 38660 246424 38712 246430
rect 38660 246366 38712 246372
rect 38672 16574 38700 246366
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36004 480 36032 16546
rect 37188 3664 37240 3670
rect 37188 3606 37240 3612
rect 37200 480 37228 3606
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 38396 480 38424 3334
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3398 39344 282134
rect 39396 260296 39448 260302
rect 39396 260238 39448 260244
rect 39408 3738 39436 260238
rect 40052 16574 40080 284990
rect 42800 278044 42852 278050
rect 42800 277986 42852 277992
rect 41420 247852 41472 247858
rect 41420 247794 41472 247800
rect 41432 16574 41460 247794
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 277986
rect 43456 3670 43484 294578
rect 52460 293276 52512 293282
rect 52460 293218 52512 293224
rect 44180 290556 44232 290562
rect 44180 290498 44232 290504
rect 44192 16574 44220 290498
rect 46940 286408 46992 286414
rect 46940 286350 46992 286356
rect 46204 251864 46256 251870
rect 46204 251806 46256 251812
rect 44192 16546 45048 16574
rect 44272 4140 44324 4146
rect 44272 4082 44324 4088
rect 43444 3664 43496 3670
rect 43444 3606 43496 3612
rect 44284 480 44312 4082
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46216 4146 46244 251806
rect 46952 16574 46980 286350
rect 48320 267028 48372 267034
rect 48320 266970 48372 266976
rect 48332 16574 48360 266970
rect 49700 251932 49752 251938
rect 49700 251874 49752 251880
rect 49712 16574 49740 251874
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 46664 3664 46716 3670
rect 46664 3606 46716 3612
rect 46676 480 46704 3606
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 4072 51408 4078
rect 51356 4014 51408 4020
rect 51368 480 51396 4014
rect 52472 3398 52500 293218
rect 58624 283688 58676 283694
rect 58624 283630 58676 283636
rect 57244 279540 57296 279546
rect 57244 279482 57296 279488
rect 53840 271176 53892 271182
rect 53840 271118 53892 271124
rect 52552 250504 52604 250510
rect 52552 250446 52604 250452
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52564 480 52592 250446
rect 53852 16574 53880 271118
rect 53852 16546 54984 16574
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54956 480 54984 16546
rect 57256 4078 57284 279482
rect 57980 272536 58032 272542
rect 57980 272478 58032 272484
rect 57336 249076 57388 249082
rect 57336 249018 57388 249024
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57348 3398 57376 249018
rect 57992 16574 58020 272478
rect 57992 16546 58480 16574
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 57336 3392 57388 3398
rect 57336 3334 57388 3340
rect 56060 480 56088 3334
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57256 480 57284 3266
rect 58452 480 58480 16546
rect 58636 3330 58664 283630
rect 60740 252000 60792 252006
rect 60740 251942 60792 251948
rect 59360 249144 59412 249150
rect 59360 249086 59412 249092
rect 58624 3324 58676 3330
rect 58624 3266 58676 3272
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59372 354 59400 249086
rect 60752 6914 60780 251942
rect 62120 250572 62172 250578
rect 62120 250514 62172 250520
rect 60832 244996 60884 245002
rect 60832 244938 60884 244944
rect 60844 16574 60872 244938
rect 62132 16574 62160 250514
rect 63512 16574 63540 296006
rect 71044 293344 71096 293350
rect 71044 293286 71096 293292
rect 67640 267096 67692 267102
rect 67640 267038 67692 267044
rect 66260 250640 66312 250646
rect 66260 250582 66312 250588
rect 64880 246492 64932 246498
rect 64880 246434 64932 246440
rect 64892 16574 64920 246434
rect 66272 16574 66300 250582
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 267038
rect 69020 261588 69072 261594
rect 69020 261530 69072 261536
rect 69032 16574 69060 261530
rect 70400 250708 70452 250714
rect 70400 250650 70452 250656
rect 70412 16574 70440 250650
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3732 69164 3738
rect 69112 3674 69164 3680
rect 69124 480 69152 3674
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3738 71084 293286
rect 81440 285116 81492 285122
rect 81440 285058 81492 285064
rect 71780 278112 71832 278118
rect 71780 278054 71832 278060
rect 71792 16574 71820 278054
rect 78680 276752 78732 276758
rect 78680 276694 78732 276700
rect 77300 271244 77352 271250
rect 77300 271186 77352 271192
rect 75920 269884 75972 269890
rect 75920 269826 75972 269832
rect 74540 268456 74592 268462
rect 74540 268398 74592 268404
rect 73160 253224 73212 253230
rect 73160 253166 73212 253172
rect 73172 16574 73200 253166
rect 74552 16574 74580 268398
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 71044 3732 71096 3738
rect 71044 3674 71096 3680
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 269826
rect 77312 6914 77340 271186
rect 77392 256080 77444 256086
rect 77392 256022 77444 256028
rect 77404 16574 77432 256022
rect 78692 16574 78720 276694
rect 80060 272604 80112 272610
rect 80060 272546 80112 272552
rect 80072 16574 80100 272546
rect 81452 16574 81480 285058
rect 82096 45558 82124 445742
rect 100024 444644 100076 444650
rect 100024 444586 100076 444592
rect 95884 444576 95936 444582
rect 95884 444518 95936 444524
rect 94504 443896 94556 443902
rect 94504 443838 94556 443844
rect 88984 440428 89036 440434
rect 88984 440370 89036 440376
rect 84200 264240 84252 264246
rect 84200 264182 84252 264188
rect 82820 249212 82872 249218
rect 82820 249154 82872 249160
rect 82084 45552 82136 45558
rect 82084 45494 82136 45500
rect 82832 16574 82860 249154
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 264182
rect 88340 254720 88392 254726
rect 88340 254662 88392 254668
rect 86960 254584 87012 254590
rect 86960 254526 87012 254532
rect 85580 249280 85632 249286
rect 85580 249222 85632 249228
rect 85592 6914 85620 249222
rect 85672 246560 85724 246566
rect 85672 246502 85724 246508
rect 85684 16574 85712 246502
rect 86972 16574 87000 254526
rect 88352 16574 88380 254662
rect 88996 33114 89024 440370
rect 94516 306338 94544 443838
rect 95896 320142 95924 444518
rect 97632 438184 97684 438190
rect 97632 438126 97684 438132
rect 97644 351121 97672 438126
rect 100036 372570 100064 444586
rect 196716 443284 196768 443290
rect 196716 443226 196768 443232
rect 192576 441992 192628 441998
rect 192576 441934 192628 441940
rect 140780 441856 140832 441862
rect 140780 441798 140832 441804
rect 140792 383654 140820 441798
rect 140792 383626 141464 383654
rect 116124 374876 116176 374882
rect 116124 374818 116176 374824
rect 103244 374808 103296 374814
rect 103244 374750 103296 374756
rect 100668 374740 100720 374746
rect 100668 374682 100720 374688
rect 100024 372564 100076 372570
rect 100024 372506 100076 372512
rect 100680 372028 100708 374682
rect 103256 372028 103284 374750
rect 108396 374332 108448 374338
rect 108396 374274 108448 374280
rect 105820 372904 105872 372910
rect 105820 372846 105872 372852
rect 105832 372028 105860 372846
rect 108408 372028 108436 374274
rect 110972 372700 111024 372706
rect 110972 372642 111024 372648
rect 110984 372028 111012 372642
rect 116136 372028 116164 374818
rect 139308 374604 139360 374610
rect 139308 374546 139360 374552
rect 121276 374536 121328 374542
rect 121276 374478 121328 374484
rect 118700 372972 118752 372978
rect 118700 372914 118752 372920
rect 118712 372028 118740 372914
rect 121288 372028 121316 374478
rect 131580 374264 131632 374270
rect 131580 374206 131632 374212
rect 126428 374196 126480 374202
rect 126428 374138 126480 374144
rect 123852 373040 123904 373046
rect 123852 372982 123904 372988
rect 123864 372028 123892 372982
rect 126440 372028 126468 374138
rect 131592 372028 131620 374206
rect 136732 372768 136784 372774
rect 134154 372736 134210 372745
rect 136732 372710 136784 372716
rect 134154 372671 134210 372680
rect 134168 372028 134196 372671
rect 136744 372028 136772 372710
rect 139320 372028 139348 374546
rect 141436 372042 141464 383626
rect 154764 374944 154816 374950
rect 154764 374886 154816 374892
rect 170404 374944 170456 374950
rect 170404 374886 170456 374892
rect 147036 374672 147088 374678
rect 147036 374614 147088 374620
rect 141436 372014 141910 372042
rect 147048 372028 147076 374614
rect 149612 372836 149664 372842
rect 149612 372778 149664 372784
rect 149624 372028 149652 372778
rect 154776 372028 154804 374886
rect 165528 374468 165580 374474
rect 165528 374410 165580 374416
rect 159914 374096 159970 374105
rect 159914 374031 159970 374040
rect 162492 374060 162544 374066
rect 157340 372632 157392 372638
rect 157340 372574 157392 372580
rect 157352 372028 157380 372574
rect 159928 372028 159956 374031
rect 162492 374002 162544 374008
rect 162504 372028 162532 374002
rect 165540 373114 165568 374410
rect 167644 374400 167696 374406
rect 167644 374342 167696 374348
rect 165068 373108 165120 373114
rect 165068 373050 165120 373056
rect 165528 373108 165580 373114
rect 165528 373050 165580 373056
rect 165080 372028 165108 373050
rect 167656 372028 167684 374342
rect 134064 371816 134116 371822
rect 133846 371764 134064 371770
rect 133846 371758 134116 371764
rect 133846 371754 134104 371758
rect 97816 371748 97868 371754
rect 97816 371690 97868 371696
rect 113456 371748 113508 371754
rect 113456 371690 113508 371696
rect 115756 371748 115808 371754
rect 115756 371690 115808 371696
rect 133834 371748 134104 371754
rect 133886 371742 134104 371748
rect 143172 371748 143224 371754
rect 133834 371690 133886 371696
rect 143172 371690 143224 371696
rect 144368 371748 144420 371754
rect 144368 371690 144420 371696
rect 97724 371680 97776 371686
rect 97724 371622 97776 371628
rect 97736 362001 97764 371622
rect 97828 364721 97856 371690
rect 113468 371618 113496 371690
rect 113574 371618 113864 371634
rect 115768 371618 115796 371690
rect 135168 371680 135220 371686
rect 133878 371648 133934 371657
rect 129030 371618 129228 371634
rect 133846 371618 133878 371634
rect 99840 371612 99892 371618
rect 99840 371554 99892 371560
rect 113456 371612 113508 371618
rect 113574 371612 113876 371618
rect 113574 371606 113824 371612
rect 113456 371554 113508 371560
rect 113824 371554 113876 371560
rect 115756 371612 115808 371618
rect 129030 371612 129240 371618
rect 129030 371606 129188 371612
rect 115756 371554 115808 371560
rect 129188 371554 129240 371560
rect 133834 371612 133878 371618
rect 133886 371583 133934 371592
rect 135166 371648 135168 371657
rect 135220 371648 135222 371657
rect 143184 371618 143212 371690
rect 143262 371648 143318 371657
rect 135166 371583 135222 371592
rect 143172 371612 143224 371618
rect 133834 371554 133886 371560
rect 144380 371618 144408 371690
rect 145012 371680 145064 371686
rect 144486 371618 144776 371634
rect 144932 371628 145012 371634
rect 153016 371680 153068 371686
rect 153014 371648 153016 371657
rect 153068 371648 153070 371657
rect 144932 371622 145064 371628
rect 144932 371618 145052 371622
rect 143262 371583 143264 371592
rect 143172 371554 143224 371560
rect 143316 371583 143318 371592
rect 144368 371612 144420 371618
rect 143264 371554 143316 371560
rect 144486 371612 144788 371618
rect 144486 371606 144736 371612
rect 144368 371554 144420 371560
rect 144736 371554 144788 371560
rect 144920 371612 145052 371618
rect 144972 371606 145052 371612
rect 152214 371618 152596 371634
rect 152214 371612 152608 371618
rect 152214 371606 152556 371612
rect 144920 371554 144972 371560
rect 153014 371583 153070 371592
rect 152556 371554 152608 371560
rect 97908 371544 97960 371550
rect 97908 371486 97960 371492
rect 97920 367441 97948 371486
rect 99852 370705 99880 371554
rect 169602 371470 169984 371498
rect 99838 370696 99894 370705
rect 99838 370631 99894 370640
rect 169956 367946 169984 371470
rect 169944 367940 169996 367946
rect 169944 367882 169996 367888
rect 97906 367432 97962 367441
rect 97906 367367 97962 367376
rect 97814 364712 97870 364721
rect 97814 364647 97870 364656
rect 97722 361992 97778 362001
rect 97722 361927 97778 361936
rect 99286 359272 99342 359281
rect 99286 359207 99342 359216
rect 99194 356552 99250 356561
rect 99194 356487 99250 356496
rect 97906 353832 97962 353841
rect 97906 353767 97962 353776
rect 97630 351112 97686 351121
rect 97630 351047 97686 351056
rect 97814 345672 97870 345681
rect 97814 345607 97870 345616
rect 97722 340232 97778 340241
rect 97722 340167 97778 340176
rect 97630 334792 97686 334801
rect 97630 334727 97686 334736
rect 97538 332072 97594 332081
rect 97538 332007 97594 332016
rect 97446 326632 97502 326641
rect 97446 326567 97502 326576
rect 97354 323912 97410 323921
rect 97354 323847 97410 323856
rect 95884 320136 95936 320142
rect 95884 320078 95936 320084
rect 97262 310312 97318 310321
rect 97262 310247 97318 310256
rect 94504 306332 94556 306338
rect 94504 306274 94556 306280
rect 97276 305538 97304 310247
rect 97092 305510 97304 305538
rect 97092 300694 97120 305510
rect 97368 305402 97396 323847
rect 97276 305374 97396 305402
rect 97460 305386 97488 326567
rect 97448 305380 97500 305386
rect 97080 300688 97132 300694
rect 97080 300630 97132 300636
rect 97276 299169 97304 305374
rect 97448 305322 97500 305328
rect 97552 305266 97580 332007
rect 97368 305238 97580 305266
rect 97262 299160 97318 299169
rect 97262 299095 97318 299104
rect 97368 298081 97396 305238
rect 97448 305176 97500 305182
rect 97644 305130 97672 334727
rect 97448 305118 97500 305124
rect 97460 300830 97488 305118
rect 97552 305102 97672 305130
rect 97448 300824 97500 300830
rect 97448 300766 97500 300772
rect 97552 299441 97580 305102
rect 97632 304972 97684 304978
rect 97632 304914 97684 304920
rect 97644 300150 97672 304914
rect 97736 300354 97764 340167
rect 97828 300626 97856 345607
rect 97920 304978 97948 353767
rect 99102 348392 99158 348401
rect 99102 348327 99158 348336
rect 99010 342952 99066 342961
rect 99010 342887 99066 342896
rect 98918 337512 98974 337521
rect 98918 337447 98974 337456
rect 98826 329352 98882 329361
rect 98826 329287 98882 329296
rect 98734 321192 98790 321201
rect 98734 321127 98790 321136
rect 98642 315752 98698 315761
rect 98642 315687 98698 315696
rect 98550 307592 98606 307601
rect 98550 307527 98606 307536
rect 97908 304972 97960 304978
rect 97908 304914 97960 304920
rect 97906 304872 97962 304881
rect 97906 304807 97962 304816
rect 97816 300620 97868 300626
rect 97816 300562 97868 300568
rect 97920 300490 97948 304807
rect 97908 300484 97960 300490
rect 97908 300426 97960 300432
rect 97724 300348 97776 300354
rect 97724 300290 97776 300296
rect 97632 300144 97684 300150
rect 97632 300086 97684 300092
rect 97538 299432 97594 299441
rect 97538 299367 97594 299376
rect 98564 299334 98592 307527
rect 98656 299402 98684 315687
rect 98644 299396 98696 299402
rect 98644 299338 98696 299344
rect 98552 299328 98604 299334
rect 98552 299270 98604 299276
rect 97354 298072 97410 298081
rect 97354 298007 97410 298016
rect 98748 297158 98776 321127
rect 98840 300082 98868 329287
rect 98932 300422 98960 337447
rect 98920 300416 98972 300422
rect 98920 300358 98972 300364
rect 98828 300076 98880 300082
rect 98828 300018 98880 300024
rect 99024 299470 99052 342887
rect 99116 300762 99144 348327
rect 99104 300756 99156 300762
rect 99104 300698 99156 300704
rect 99012 299464 99064 299470
rect 99012 299406 99064 299412
rect 99208 299305 99236 356487
rect 99300 300801 99328 359207
rect 99378 318472 99434 318481
rect 99378 318407 99434 318416
rect 99286 300792 99342 300801
rect 99286 300727 99342 300736
rect 99392 300558 99420 318407
rect 99470 313032 99526 313041
rect 99470 312967 99526 312976
rect 99380 300552 99432 300558
rect 99380 300494 99432 300500
rect 99484 300218 99512 312967
rect 170416 307018 170444 374886
rect 170956 374876 171008 374882
rect 170956 374818 171008 374824
rect 170772 374536 170824 374542
rect 170772 374478 170824 374484
rect 170496 374060 170548 374066
rect 170496 374002 170548 374008
rect 170508 307222 170536 374002
rect 170588 373040 170640 373046
rect 170588 372982 170640 372988
rect 170600 308582 170628 372982
rect 170680 367940 170732 367946
rect 170680 367882 170732 367888
rect 170692 309194 170720 367882
rect 170784 309505 170812 374478
rect 170770 309496 170826 309505
rect 170770 309431 170826 309440
rect 170968 309369 170996 374818
rect 174728 374672 174780 374678
rect 174728 374614 174780 374620
rect 171784 374604 171836 374610
rect 171784 374546 171836 374552
rect 171690 358592 171746 358601
rect 171690 358527 171746 358536
rect 171704 357474 171732 358527
rect 171692 357468 171744 357474
rect 171692 357410 171744 357416
rect 171796 354674 171824 374546
rect 174544 372972 174596 372978
rect 174544 372914 174596 372920
rect 173164 372632 173216 372638
rect 173164 372574 173216 372580
rect 172334 369472 172390 369481
rect 172334 369407 172390 369416
rect 172348 368558 172376 369407
rect 172336 368552 172388 368558
rect 172336 368494 172388 368500
rect 172426 366752 172482 366761
rect 172426 366687 172482 366696
rect 172440 365770 172468 366687
rect 172428 365764 172480 365770
rect 172428 365706 172480 365712
rect 171874 364032 171930 364041
rect 171874 363967 171930 363976
rect 171704 354646 171824 354674
rect 171704 350690 171732 354646
rect 171612 350662 171732 350690
rect 171140 349172 171192 349178
rect 171140 349114 171192 349120
rect 170954 309360 171010 309369
rect 170954 309295 171010 309304
rect 170680 309188 170732 309194
rect 170680 309130 170732 309136
rect 170588 308576 170640 308582
rect 170588 308518 170640 308524
rect 170496 307216 170548 307222
rect 170496 307158 170548 307164
rect 170588 307148 170640 307154
rect 170588 307090 170640 307096
rect 170404 307012 170456 307018
rect 170404 306954 170456 306960
rect 170404 305788 170456 305794
rect 170404 305730 170456 305736
rect 169944 304632 169996 304638
rect 169944 304574 169996 304580
rect 169852 304564 169904 304570
rect 169852 304506 169904 304512
rect 169760 303068 169812 303074
rect 169760 303010 169812 303016
rect 99838 302152 99894 302161
rect 99838 302087 99894 302096
rect 99852 300286 99880 302087
rect 169772 300778 169800 303010
rect 169680 300750 169800 300778
rect 169680 300642 169708 300750
rect 168958 300614 169708 300642
rect 164238 300384 164294 300393
rect 164238 300319 164294 300328
rect 99840 300280 99892 300286
rect 99840 300222 99892 300228
rect 160098 300248 160154 300257
rect 99472 300212 99524 300218
rect 160098 300183 160154 300192
rect 99472 300154 99524 300160
rect 99194 299296 99250 299305
rect 99194 299231 99250 299240
rect 100036 297702 100064 300084
rect 100024 297696 100076 297702
rect 100024 297638 100076 297644
rect 101968 297634 101996 300084
rect 104544 299266 104572 300084
rect 104532 299260 104584 299266
rect 104532 299202 104584 299208
rect 101956 297628 102008 297634
rect 101956 297570 102008 297576
rect 107120 297566 107148 300084
rect 109696 297945 109724 300084
rect 109682 297936 109738 297945
rect 109682 297871 109738 297880
rect 107108 297560 107160 297566
rect 107108 297502 107160 297508
rect 98736 297152 98788 297158
rect 98736 297094 98788 297100
rect 112272 297090 112300 300084
rect 114848 299198 114876 300084
rect 114836 299192 114888 299198
rect 114836 299134 114888 299140
rect 117424 299062 117452 300084
rect 120000 299130 120028 300084
rect 119988 299124 120040 299130
rect 119988 299066 120040 299072
rect 117412 299056 117464 299062
rect 117412 298998 117464 299004
rect 122576 297906 122604 300084
rect 125152 298926 125180 300084
rect 126992 300070 127742 300098
rect 125140 298920 125192 298926
rect 125140 298862 125192 298868
rect 122564 297900 122616 297906
rect 122564 297842 122616 297848
rect 112260 297084 112312 297090
rect 112260 297026 112312 297032
rect 126992 296682 127020 300070
rect 130304 298994 130332 300084
rect 130292 298988 130344 298994
rect 130292 298930 130344 298936
rect 132880 297974 132908 300084
rect 132868 297968 132920 297974
rect 132868 297910 132920 297916
rect 135456 297498 135484 300084
rect 138032 297838 138060 300084
rect 140608 298858 140636 300084
rect 140596 298852 140648 298858
rect 140596 298794 140648 298800
rect 138020 297832 138072 297838
rect 138020 297774 138072 297780
rect 135444 297492 135496 297498
rect 135444 297434 135496 297440
rect 143184 297430 143212 300084
rect 145760 298722 145788 300084
rect 145748 298716 145800 298722
rect 145748 298658 145800 298664
rect 148336 297770 148364 300084
rect 150912 297809 150940 300084
rect 153212 300070 153502 300098
rect 150898 297800 150954 297809
rect 148324 297764 148376 297770
rect 150898 297735 150954 297744
rect 148324 297706 148376 297712
rect 143172 297424 143224 297430
rect 143172 297366 143224 297372
rect 126980 296676 127032 296682
rect 126980 296618 127032 296624
rect 153212 296614 153240 300070
rect 156064 298790 156092 300084
rect 156052 298784 156104 298790
rect 156052 298726 156104 298732
rect 158640 298110 158668 300084
rect 158628 298104 158680 298110
rect 158628 298046 158680 298052
rect 153200 296608 153252 296614
rect 153200 296550 153252 296556
rect 129740 296200 129792 296206
rect 129740 296142 129792 296148
rect 125600 296132 125652 296138
rect 125600 296074 125652 296080
rect 103520 289196 103572 289202
rect 103520 289138 103572 289144
rect 98000 278180 98052 278186
rect 98000 278122 98052 278128
rect 93860 275392 93912 275398
rect 93860 275334 93912 275340
rect 92480 269952 92532 269958
rect 92480 269894 92532 269900
rect 91100 254652 91152 254658
rect 91100 254594 91152 254600
rect 89720 247920 89772 247926
rect 89720 247862 89772 247868
rect 88984 33108 89036 33114
rect 88984 33050 89036 33056
rect 89732 16574 89760 247862
rect 91112 16574 91140 254594
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 269894
rect 93872 6914 93900 275334
rect 93952 273964 94004 273970
rect 93952 273906 94004 273912
rect 93964 16574 93992 273906
rect 96620 264308 96672 264314
rect 96620 264250 96672 264256
rect 95240 253292 95292 253298
rect 95240 253234 95292 253240
rect 95252 16574 95280 253234
rect 96632 16574 96660 264250
rect 98012 16574 98040 278122
rect 102140 276820 102192 276826
rect 102140 276762 102192 276768
rect 99380 271312 99432 271318
rect 99380 271254 99432 271260
rect 99392 16574 99420 271254
rect 100760 245064 100812 245070
rect 100760 245006 100812 245012
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 245006
rect 102152 6914 102180 276762
rect 102232 272672 102284 272678
rect 102232 272614 102284 272620
rect 102244 16574 102272 272614
rect 103532 16574 103560 289138
rect 107660 282260 107712 282266
rect 107660 282202 107712 282208
rect 106280 257508 106332 257514
rect 106280 257450 106332 257456
rect 104900 245132 104952 245138
rect 104900 245074 104952 245080
rect 104912 16574 104940 245074
rect 106292 16574 106320 257450
rect 107672 16574 107700 282202
rect 111800 275460 111852 275466
rect 111800 275402 111852 275408
rect 110420 254788 110472 254794
rect 110420 254730 110472 254736
rect 109040 246628 109092 246634
rect 109040 246570 109092 246576
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 246570
rect 110432 6914 110460 254730
rect 110512 253360 110564 253366
rect 110512 253302 110564 253308
rect 110524 16574 110552 253302
rect 111812 16574 111840 275402
rect 120080 274032 120132 274038
rect 120080 273974 120132 273980
rect 115940 265804 115992 265810
rect 115940 265746 115992 265752
rect 114560 265736 114612 265742
rect 114560 265678 114612 265684
rect 113180 264376 113232 264382
rect 113180 264318 113232 264324
rect 113192 16574 113220 264318
rect 114572 16574 114600 265678
rect 115952 16574 115980 265746
rect 117320 257576 117372 257582
rect 117320 257518 117372 257524
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 257518
rect 118700 256148 118752 256154
rect 118700 256090 118752 256096
rect 118712 3398 118740 256090
rect 118792 253428 118844 253434
rect 118792 253370 118844 253376
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 253370
rect 120092 16574 120120 273974
rect 124220 260364 124272 260370
rect 124220 260306 124272 260312
rect 122840 256216 122892 256222
rect 122840 256158 122892 256164
rect 121460 246696 121512 246702
rect 121460 246638 121512 246644
rect 121472 16574 121500 246638
rect 122852 16574 122880 256158
rect 124232 16574 124260 260306
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 296074
rect 128360 291916 128412 291922
rect 128360 291858 128412 291864
rect 126980 280900 127032 280906
rect 126980 280842 127032 280848
rect 126992 480 127020 280842
rect 127072 275528 127124 275534
rect 127072 275470 127124 275476
rect 127084 16574 127112 275470
rect 128372 16574 128400 291858
rect 129752 16574 129780 296142
rect 135260 294704 135312 294710
rect 135260 294646 135312 294652
rect 132500 289264 132552 289270
rect 132500 289206 132552 289212
rect 131120 282328 131172 282334
rect 131120 282270 131172 282276
rect 131132 16574 131160 282270
rect 132512 16574 132540 289206
rect 133880 265872 133932 265878
rect 133880 265814 133932 265820
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 265814
rect 135272 3738 135300 294646
rect 151820 290760 151872 290766
rect 151820 290702 151872 290708
rect 143540 290624 143592 290630
rect 143540 290566 143592 290572
rect 139400 287768 139452 287774
rect 139400 287710 139452 287716
rect 138020 283756 138072 283762
rect 138020 283698 138072 283704
rect 136640 276888 136692 276894
rect 136640 276830 136692 276836
rect 135352 250776 135404 250782
rect 135352 250718 135404 250724
rect 135260 3732 135312 3738
rect 135260 3674 135312 3680
rect 135364 3482 135392 250718
rect 136652 16574 136680 276830
rect 138032 16574 138060 283698
rect 139412 16574 139440 287710
rect 142160 280968 142212 280974
rect 142160 280910 142212 280916
rect 140780 247988 140832 247994
rect 140780 247930 140832 247936
rect 140792 16574 140820 247930
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 3732 136508 3738
rect 136456 3674 136508 3680
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3674
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 280910
rect 143552 480 143580 290566
rect 146300 286476 146352 286482
rect 146300 286418 146352 286424
rect 144920 268524 144972 268530
rect 144920 268466 144972 268472
rect 143632 264444 143684 264450
rect 143632 264386 143684 264392
rect 143644 16574 143672 264386
rect 144932 16574 144960 268466
rect 146312 16574 146340 286418
rect 150440 285184 150492 285190
rect 150440 285126 150492 285132
rect 147680 278248 147732 278254
rect 147680 278190 147732 278196
rect 147692 16574 147720 278190
rect 149060 261724 149112 261730
rect 149060 261666 149112 261672
rect 149072 16574 149100 261666
rect 150452 16574 150480 285126
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 290702
rect 153200 283892 153252 283898
rect 153200 283834 153252 283840
rect 151912 262880 151964 262886
rect 151912 262822 151964 262828
rect 151924 16574 151952 262822
rect 153212 16574 153240 283834
rect 157340 282396 157392 282402
rect 157340 282338 157392 282344
rect 154580 262948 154632 262954
rect 154580 262890 154632 262896
rect 154592 16574 154620 262890
rect 155960 252136 156012 252142
rect 155960 252078 156012 252084
rect 155972 16574 156000 252078
rect 157352 16574 157380 282338
rect 158720 261792 158772 261798
rect 158720 261734 158772 261740
rect 158732 16574 158760 261734
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11762 160140 300183
rect 161216 298654 161244 300084
rect 161204 298648 161256 298654
rect 161204 298590 161256 298596
rect 163792 298586 163820 300084
rect 163780 298580 163832 298586
rect 163780 298522 163832 298528
rect 161480 291984 161532 291990
rect 161480 291926 161532 291932
rect 160192 252204 160244 252210
rect 160192 252146 160244 252152
rect 160100 11756 160152 11762
rect 160100 11698 160152 11704
rect 160204 6914 160232 252146
rect 161492 16574 161520 291926
rect 162860 274100 162912 274106
rect 162860 274042 162912 274048
rect 162872 16574 162900 274042
rect 164252 16574 164280 300319
rect 166368 298110 166396 300084
rect 166356 298104 166408 298110
rect 166356 298046 166408 298052
rect 169864 298042 169892 304506
rect 169852 298036 169904 298042
rect 169852 297978 169904 297984
rect 169956 297566 169984 304574
rect 169944 297560 169996 297566
rect 169944 297502 169996 297508
rect 168380 294772 168432 294778
rect 168380 294714 168432 294720
rect 165620 279608 165672 279614
rect 165620 279550 165672 279556
rect 165632 16574 165660 279550
rect 167000 270020 167052 270026
rect 167000 269962 167052 269968
rect 167012 16574 167040 269962
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11756 161348 11762
rect 161296 11698 161348 11704
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11698
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 294714
rect 169760 254856 169812 254862
rect 169760 254798 169812 254804
rect 168472 245200 168524 245206
rect 168472 245142 168524 245148
rect 168484 16574 168512 245142
rect 169772 16574 169800 254798
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 169588 480 169616 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 170416 3534 170444 305730
rect 170494 302968 170550 302977
rect 170494 302903 170550 302912
rect 170508 3670 170536 302903
rect 170600 298110 170628 307090
rect 170588 298104 170640 298110
rect 170588 298046 170640 298052
rect 170496 3664 170548 3670
rect 170496 3606 170548 3612
rect 170404 3528 170456 3534
rect 170404 3470 170456 3476
rect 171152 3466 171180 349114
rect 171612 345014 171640 350662
rect 171888 350538 171916 363967
rect 171966 361312 172022 361321
rect 171966 361247 172022 361256
rect 171692 350532 171744 350538
rect 171692 350474 171744 350480
rect 171876 350532 171928 350538
rect 171876 350474 171928 350480
rect 171704 349058 171732 350474
rect 171874 350432 171930 350441
rect 171874 350367 171930 350376
rect 171888 349178 171916 350367
rect 171876 349172 171928 349178
rect 171876 349114 171928 349120
rect 171704 349030 171916 349058
rect 171612 344986 171824 345014
rect 171414 325952 171470 325961
rect 171414 325887 171470 325896
rect 171428 325718 171456 325887
rect 171416 325712 171468 325718
rect 171416 325654 171468 325660
rect 171796 311302 171824 344986
rect 171784 311296 171836 311302
rect 171784 311238 171836 311244
rect 171888 310622 171916 349030
rect 171980 311234 172008 361247
rect 172426 355872 172482 355881
rect 172426 355807 172482 355816
rect 172440 354754 172468 355807
rect 172428 354748 172480 354754
rect 172428 354690 172480 354696
rect 172426 353152 172482 353161
rect 172426 353087 172482 353096
rect 172440 351966 172468 353087
rect 172428 351960 172480 351966
rect 172428 351902 172480 351908
rect 172426 347712 172482 347721
rect 172426 347647 172482 347656
rect 172440 346458 172468 347647
rect 172428 346452 172480 346458
rect 172428 346394 172480 346400
rect 172058 344992 172114 345001
rect 172058 344927 172114 344936
rect 171968 311228 172020 311234
rect 171968 311170 172020 311176
rect 172072 310865 172100 344927
rect 172428 342304 172480 342310
rect 172426 342272 172428 342281
rect 172480 342272 172482 342281
rect 172426 342207 172482 342216
rect 172150 339552 172206 339561
rect 172150 339487 172206 339496
rect 172164 311370 172192 339487
rect 172426 336832 172482 336841
rect 172426 336767 172428 336776
rect 172480 336767 172482 336776
rect 172428 336738 172480 336744
rect 172426 334112 172482 334121
rect 172426 334047 172482 334056
rect 172440 334014 172468 334047
rect 172428 334008 172480 334014
rect 172428 333950 172480 333956
rect 172426 331392 172482 331401
rect 172426 331327 172482 331336
rect 172440 331294 172468 331327
rect 172428 331288 172480 331294
rect 172428 331230 172480 331236
rect 172426 328672 172482 328681
rect 172426 328607 172482 328616
rect 172440 328506 172468 328607
rect 172428 328500 172480 328506
rect 172428 328442 172480 328448
rect 172242 323232 172298 323241
rect 172242 323167 172298 323176
rect 172152 311364 172204 311370
rect 172152 311306 172204 311312
rect 172058 310856 172114 310865
rect 172058 310791 172114 310800
rect 171876 310616 171928 310622
rect 171876 310558 171928 310564
rect 172256 310010 172284 323167
rect 172426 320512 172482 320521
rect 172426 320447 172482 320456
rect 172440 320210 172468 320447
rect 172428 320204 172480 320210
rect 172428 320146 172480 320152
rect 172426 317792 172482 317801
rect 172426 317727 172482 317736
rect 172440 317490 172468 317727
rect 172428 317484 172480 317490
rect 172428 317426 172480 317432
rect 172426 315072 172482 315081
rect 172426 315007 172482 315016
rect 172440 314702 172468 315007
rect 172428 314696 172480 314702
rect 172428 314638 172480 314644
rect 172426 312352 172482 312361
rect 172426 312287 172482 312296
rect 172440 311914 172468 312287
rect 172428 311908 172480 311914
rect 172428 311850 172480 311856
rect 172428 310072 172480 310078
rect 172428 310014 172480 310020
rect 172244 310004 172296 310010
rect 172244 309946 172296 309952
rect 172440 309641 172468 310014
rect 172426 309632 172482 309641
rect 172426 309567 172482 309576
rect 173176 308718 173204 372574
rect 173256 371748 173308 371754
rect 173256 371690 173308 371696
rect 173164 308712 173216 308718
rect 173164 308654 173216 308660
rect 173268 308281 173296 371690
rect 174556 308378 174584 372914
rect 174636 372904 174688 372910
rect 174636 372846 174688 372852
rect 174648 308961 174676 372846
rect 174740 309233 174768 374614
rect 175924 374332 175976 374338
rect 175924 374274 175976 374280
rect 174726 309224 174782 309233
rect 174726 309159 174782 309168
rect 174634 308952 174690 308961
rect 174634 308887 174690 308896
rect 174544 308372 174596 308378
rect 174544 308314 174596 308320
rect 173254 308272 173310 308281
rect 173254 308207 173310 308216
rect 175936 307562 175964 374274
rect 192484 349172 192536 349178
rect 192484 349114 192536 349120
rect 192496 311166 192524 349114
rect 192484 311160 192536 311166
rect 192484 311102 192536 311108
rect 175924 307556 175976 307562
rect 175924 307498 175976 307504
rect 172428 307284 172480 307290
rect 172428 307226 172480 307232
rect 172440 306921 172468 307226
rect 172426 306912 172482 306921
rect 172426 306847 172482 306856
rect 171692 306196 171744 306202
rect 171692 306138 171744 306144
rect 171416 304428 171468 304434
rect 171416 304370 171468 304376
rect 171428 297634 171456 304370
rect 171416 297628 171468 297634
rect 171416 297570 171468 297576
rect 171704 297498 171732 306138
rect 178040 305652 178092 305658
rect 178040 305594 178092 305600
rect 172152 305448 172204 305454
rect 172152 305390 172204 305396
rect 171784 301572 171836 301578
rect 171784 301514 171836 301520
rect 171692 297492 171744 297498
rect 171692 297434 171744 297440
rect 171232 245268 171284 245274
rect 171232 245210 171284 245216
rect 171244 16574 171272 245210
rect 171244 16546 171732 16574
rect 171704 3482 171732 16546
rect 171796 3602 171824 301514
rect 172164 297362 172192 305390
rect 172336 304972 172388 304978
rect 172336 304914 172388 304920
rect 172244 304496 172296 304502
rect 172244 304438 172296 304444
rect 172256 297702 172284 304438
rect 172348 304201 172376 304914
rect 172334 304192 172390 304201
rect 172334 304127 172390 304136
rect 172428 302184 172480 302190
rect 172428 302126 172480 302132
rect 172440 301481 172468 302126
rect 172426 301472 172482 301481
rect 172426 301407 172482 301416
rect 172244 297696 172296 297702
rect 172244 297638 172296 297644
rect 172152 297356 172204 297362
rect 172152 297298 172204 297304
rect 176660 258868 176712 258874
rect 176660 258810 176712 258816
rect 173900 258800 173952 258806
rect 173900 258742 173952 258748
rect 172520 252272 172572 252278
rect 172520 252214 172572 252220
rect 172532 16574 172560 252214
rect 172532 16546 172744 16574
rect 171784 3596 171836 3602
rect 171784 3538 171836 3544
rect 171140 3460 171192 3466
rect 171704 3454 172008 3482
rect 171140 3402 171192 3408
rect 171980 480 172008 3454
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 258742
rect 175280 248056 175332 248062
rect 175280 247998 175332 248004
rect 175292 16574 175320 247998
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 11762 176700 258810
rect 176752 253564 176804 253570
rect 176752 253506 176804 253512
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 176764 6914 176792 253506
rect 178052 16574 178080 305594
rect 189080 304292 189132 304298
rect 189080 304234 189132 304240
rect 184940 302932 184992 302938
rect 184940 302874 184992 302880
rect 182178 302832 182234 302841
rect 182178 302767 182234 302776
rect 181444 287836 181496 287842
rect 181444 287778 181496 287784
rect 180800 271380 180852 271386
rect 180800 271322 180852 271328
rect 180812 16574 180840 271322
rect 178052 16546 178632 16574
rect 180812 16546 181024 16574
rect 177856 11756 177908 11762
rect 177856 11698 177908 11704
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11698
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180248 4140 180300 4146
rect 180248 4082 180300 4088
rect 180260 480 180288 4082
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 4146 181484 287778
rect 181444 4140 181496 4146
rect 181444 4082 181496 4088
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 302767
rect 184952 11762 184980 302874
rect 188344 278316 188396 278322
rect 188344 278258 188396 278264
rect 187700 272740 187752 272746
rect 187700 272682 187752 272688
rect 185032 249348 185084 249354
rect 185032 249290 185084 249296
rect 184940 11756 184992 11762
rect 184940 11698 184992 11704
rect 185044 6914 185072 249290
rect 187712 16574 187740 272682
rect 187712 16546 188292 16574
rect 186136 11756 186188 11762
rect 186136 11698 186188 11704
rect 184952 6886 185072 6914
rect 183744 3596 183796 3602
rect 183744 3538 183796 3544
rect 183756 480 183784 3538
rect 184952 480 184980 6886
rect 186148 480 186176 11698
rect 187332 3664 187384 3670
rect 187332 3606 187384 3612
rect 187344 480 187372 3606
rect 188264 3482 188292 16546
rect 188356 3602 188384 278258
rect 189092 16574 189120 304234
rect 191840 265940 191892 265946
rect 191840 265882 191892 265888
rect 191852 16574 191880 265882
rect 192588 20670 192616 441934
rect 195980 305720 196032 305726
rect 195980 305662 196032 305668
rect 193220 301504 193272 301510
rect 193220 301446 193272 301452
rect 192576 20664 192628 20670
rect 192576 20606 192628 20612
rect 189092 16546 189304 16574
rect 191852 16546 192064 16574
rect 188344 3596 188396 3602
rect 188344 3538 188396 3544
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 190828 3460 190880 3466
rect 190828 3402 190880 3408
rect 190840 480 190868 3402
rect 192036 480 192064 16546
rect 193232 480 193260 301446
rect 193312 275596 193364 275602
rect 193312 275538 193364 275544
rect 193324 16574 193352 275538
rect 195992 16574 196020 305662
rect 196624 276956 196676 276962
rect 196624 276898 196676 276904
rect 193324 16546 194456 16574
rect 195992 16546 196572 16574
rect 194428 480 194456 16546
rect 195612 3596 195664 3602
rect 195612 3538 195664 3544
rect 195624 480 195652 3538
rect 196544 3482 196572 16546
rect 196636 3670 196664 276898
rect 196728 202842 196756 443226
rect 198004 442060 198056 442066
rect 198004 442002 198056 442008
rect 197360 274168 197412 274174
rect 197360 274110 197412 274116
rect 196716 202836 196768 202842
rect 196716 202778 196768 202784
rect 197372 16574 197400 274110
rect 198016 97986 198044 442002
rect 198740 248124 198792 248130
rect 198740 248066 198792 248072
rect 198004 97980 198056 97986
rect 198004 97922 198056 97928
rect 197372 16546 197952 16574
rect 196624 3664 196676 3670
rect 196624 3606 196676 3612
rect 196544 3454 196848 3482
rect 196820 480 196848 3454
rect 197924 480 197952 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 248066
rect 199396 150414 199424 446082
rect 200764 446072 200816 446078
rect 200764 446014 200816 446020
rect 200120 307080 200172 307086
rect 200120 307022 200172 307028
rect 199476 286544 199528 286550
rect 199476 286486 199528 286492
rect 199384 150408 199436 150414
rect 199384 150350 199436 150356
rect 199488 3466 199516 286486
rect 200132 16574 200160 307022
rect 200132 16546 200344 16574
rect 199476 3460 199528 3466
rect 199476 3402 199528 3408
rect 200316 480 200344 16546
rect 200776 6866 200804 446014
rect 202880 293412 202932 293418
rect 202880 293354 202932 293360
rect 201500 289332 201552 289338
rect 201500 289274 201552 289280
rect 201512 11762 201540 289274
rect 201592 272808 201644 272814
rect 201592 272750 201644 272756
rect 201500 11756 201552 11762
rect 201500 11698 201552 11704
rect 201604 6914 201632 272750
rect 202892 16574 202920 293354
rect 203536 137970 203564 446150
rect 215944 444848 215996 444854
rect 215944 444790 215996 444796
rect 206284 442128 206336 442134
rect 206284 442070 206336 442076
rect 205640 300008 205692 300014
rect 205640 299950 205692 299956
rect 203616 245336 203668 245342
rect 203616 245278 203668 245284
rect 203524 137964 203576 137970
rect 203524 137906 203576 137912
rect 202892 16546 203472 16574
rect 202696 11756 202748 11762
rect 202696 11698 202748 11704
rect 201512 6886 201632 6914
rect 200764 6860 200816 6866
rect 200764 6802 200816 6808
rect 201512 480 201540 6886
rect 202708 480 202736 11698
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 203628 3602 203656 245278
rect 205652 16574 205680 299950
rect 206296 85542 206324 442070
rect 207664 440700 207716 440706
rect 207664 440642 207716 440648
rect 207020 304360 207072 304366
rect 207020 304302 207072 304308
rect 206284 85536 206336 85542
rect 206284 85478 206336 85484
rect 205652 16546 206232 16574
rect 203616 3596 203668 3602
rect 203616 3538 203668 3544
rect 205086 3360 205142 3369
rect 205086 3295 205142 3304
rect 205100 480 205128 3295
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 304302
rect 207676 71738 207704 440642
rect 215208 306128 215260 306134
rect 215208 306070 215260 306076
rect 214932 305992 214984 305998
rect 214932 305934 214984 305940
rect 213828 305856 213880 305862
rect 213828 305798 213880 305804
rect 212448 303408 212500 303414
rect 212448 303350 212500 303356
rect 212080 303136 212132 303142
rect 212080 303078 212132 303084
rect 210976 301776 211028 301782
rect 210976 301718 211028 301724
rect 210884 297492 210936 297498
rect 210884 297434 210936 297440
rect 209780 296268 209832 296274
rect 209780 296210 209832 296216
rect 207664 71732 207716 71738
rect 207664 71674 207716 71680
rect 209792 9674 209820 296210
rect 210700 294908 210752 294914
rect 210700 294850 210752 294856
rect 209872 250844 209924 250850
rect 209872 250786 209924 250792
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 250786
rect 210712 155582 210740 294850
rect 210792 294840 210844 294846
rect 210792 294782 210844 294788
rect 210700 155576 210752 155582
rect 210700 155518 210752 155524
rect 210804 155281 210832 294782
rect 210896 155514 210924 297434
rect 210884 155508 210936 155514
rect 210884 155450 210936 155456
rect 210988 155417 211016 301718
rect 211896 301640 211948 301646
rect 211896 301582 211948 301588
rect 211712 297424 211764 297430
rect 211712 297366 211764 297372
rect 211068 294976 211120 294982
rect 211068 294918 211120 294924
rect 210974 155408 211030 155417
rect 210974 155343 211030 155352
rect 210790 155272 210846 155281
rect 210790 155207 210846 155216
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 208584 3324 208636 3330
rect 208584 3266 208636 3272
rect 208596 480 208624 3266
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 211080 3806 211108 294918
rect 211724 159458 211752 297366
rect 211804 271448 211856 271454
rect 211804 271390 211856 271396
rect 211712 159452 211764 159458
rect 211712 159394 211764 159400
rect 211068 3800 211120 3806
rect 211068 3742 211120 3748
rect 211816 3330 211844 271390
rect 211908 158778 211936 301582
rect 211986 297528 212042 297537
rect 211986 297463 212042 297472
rect 211896 158772 211948 158778
rect 211896 158714 211948 158720
rect 212000 155854 212028 297463
rect 212092 158642 212120 303078
rect 212172 301708 212224 301714
rect 212172 301650 212224 301656
rect 212080 158636 212132 158642
rect 212080 158578 212132 158584
rect 211988 155848 212040 155854
rect 211988 155790 212040 155796
rect 212184 155242 212212 301650
rect 212354 297392 212410 297401
rect 212354 297327 212410 297336
rect 212264 295044 212316 295050
rect 212264 294986 212316 294992
rect 212172 155236 212224 155242
rect 212172 155178 212224 155184
rect 212276 3738 212304 294986
rect 212368 4078 212396 297327
rect 212356 4072 212408 4078
rect 212356 4014 212408 4020
rect 212264 3732 212316 3738
rect 212264 3674 212316 3680
rect 212170 3632 212226 3641
rect 212170 3567 212226 3576
rect 211804 3324 211856 3330
rect 211804 3266 211856 3272
rect 212184 480 212212 3567
rect 212460 3398 212488 303350
rect 213644 303000 213696 303006
rect 213644 302942 213696 302948
rect 213368 299940 213420 299946
rect 213368 299882 213420 299888
rect 213276 297560 213328 297566
rect 213276 297502 213328 297508
rect 212540 261860 212592 261866
rect 212540 261802 212592 261808
rect 212552 16574 212580 261802
rect 213288 158710 213316 297502
rect 213276 158704 213328 158710
rect 213276 158646 213328 158652
rect 213380 158506 213408 299882
rect 213550 297664 213606 297673
rect 213550 297599 213606 297608
rect 213460 297356 213512 297362
rect 213460 297298 213512 297304
rect 213368 158500 213420 158506
rect 213368 158442 213420 158448
rect 213472 155650 213500 297298
rect 213564 155786 213592 297599
rect 213656 159526 213684 302942
rect 213736 297628 213788 297634
rect 213736 297570 213788 297576
rect 213644 159520 213696 159526
rect 213644 159462 213696 159468
rect 213552 155780 213604 155786
rect 213552 155722 213604 155728
rect 213460 155644 213512 155650
rect 213460 155586 213512 155592
rect 212552 16546 213408 16574
rect 212448 3392 212500 3398
rect 212448 3334 212500 3340
rect 213380 480 213408 16546
rect 213748 4010 213776 297570
rect 213736 4004 213788 4010
rect 213736 3946 213788 3952
rect 213840 3942 213868 305798
rect 214840 303476 214892 303482
rect 214840 303418 214892 303424
rect 214564 303204 214616 303210
rect 214564 303146 214616 303152
rect 214472 297696 214524 297702
rect 214472 297638 214524 297644
rect 214380 295112 214432 295118
rect 214380 295054 214432 295060
rect 214392 213926 214420 295054
rect 214380 213920 214432 213926
rect 214380 213862 214432 213868
rect 214484 155378 214512 297638
rect 214576 158370 214604 303146
rect 214656 302864 214708 302870
rect 214656 302806 214708 302812
rect 214564 158364 214616 158370
rect 214564 158306 214616 158312
rect 214668 157826 214696 302806
rect 214748 302728 214800 302734
rect 214748 302670 214800 302676
rect 214760 157865 214788 302670
rect 214852 158574 214880 303418
rect 214840 158568 214892 158574
rect 214840 158510 214892 158516
rect 214944 158302 214972 305934
rect 215116 295180 215168 295186
rect 215116 295122 215168 295128
rect 215024 294568 215076 294574
rect 215024 294510 215076 294516
rect 214932 158296 214984 158302
rect 214932 158238 214984 158244
rect 214746 157856 214802 157865
rect 214656 157820 214708 157826
rect 214746 157791 214802 157800
rect 214656 157762 214708 157768
rect 214472 155372 214524 155378
rect 214472 155314 214524 155320
rect 213828 3936 213880 3942
rect 213828 3878 213880 3884
rect 215036 3874 215064 294510
rect 215024 3868 215076 3874
rect 215024 3810 215076 3816
rect 214470 3496 214526 3505
rect 215128 3466 215156 295122
rect 214470 3431 214526 3440
rect 215116 3460 215168 3466
rect 214484 480 214512 3431
rect 215116 3402 215168 3408
rect 215220 3330 215248 306070
rect 215852 297288 215904 297294
rect 215852 297230 215904 297236
rect 215760 295248 215812 295254
rect 215760 295190 215812 295196
rect 215772 195430 215800 295190
rect 215760 195424 215812 195430
rect 215760 195366 215812 195372
rect 215864 159390 215892 297230
rect 215956 215286 215984 444790
rect 217796 443698 217824 565082
rect 217888 478650 217916 700266
rect 217876 478644 217928 478650
rect 217876 478586 217928 478592
rect 217980 478582 218008 700334
rect 217968 478576 218020 478582
rect 217968 478518 218020 478524
rect 218072 464438 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 219348 700460 219400 700466
rect 219348 700402 219400 700408
rect 219162 512816 219218 512825
rect 219162 512751 219218 512760
rect 219070 509960 219126 509969
rect 219070 509895 219126 509904
rect 218978 508192 219034 508201
rect 218978 508127 219034 508136
rect 218886 488336 218942 488345
rect 218886 488271 218942 488280
rect 218900 465866 218928 488271
rect 218992 478310 219020 508127
rect 218980 478304 219032 478310
rect 218980 478246 219032 478252
rect 219084 474162 219112 509895
rect 219176 475454 219204 512751
rect 219254 511048 219310 511057
rect 219254 510983 219310 510992
rect 219164 475448 219216 475454
rect 219164 475390 219216 475396
rect 219072 474156 219124 474162
rect 219072 474098 219124 474104
rect 219268 468654 219296 510983
rect 219256 468648 219308 468654
rect 219256 468590 219308 468596
rect 218888 465860 218940 465866
rect 218888 465802 218940 465808
rect 218060 464432 218112 464438
rect 218060 464374 218112 464380
rect 219360 443766 219388 700402
rect 234632 565146 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700466 267688 703520
rect 267648 700460 267700 700466
rect 267648 700402 267700 700408
rect 283852 700398 283880 703520
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 300136 700330 300164 703520
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 358820 700392 358872 700398
rect 358820 700334 358872 700340
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 357440 700324 357492 700330
rect 357440 700266 357492 700272
rect 234620 565140 234672 565146
rect 234620 565082 234672 565088
rect 269948 478644 270000 478650
rect 269948 478586 270000 478592
rect 268660 478508 268712 478514
rect 268660 478450 268712 478456
rect 256884 478236 256936 478242
rect 256884 478178 256936 478184
rect 238482 477320 238538 477329
rect 238482 477255 238538 477264
rect 238496 476814 238524 477255
rect 242806 477184 242862 477193
rect 242806 477119 242862 477128
rect 240046 476912 240102 476921
rect 240046 476847 240102 476856
rect 241426 476912 241482 476921
rect 241426 476847 241428 476856
rect 238484 476808 238536 476814
rect 237286 476776 237342 476785
rect 238484 476750 238536 476756
rect 237286 476711 237288 476720
rect 237340 476711 237342 476720
rect 239404 476740 239456 476746
rect 237288 476682 237340 476688
rect 239404 476682 239456 476688
rect 237194 476232 237250 476241
rect 237194 476167 237250 476176
rect 237208 447982 237236 476167
rect 239416 460426 239444 476682
rect 240060 476134 240088 476847
rect 241480 476847 241482 476856
rect 241428 476818 241480 476824
rect 242820 476678 242848 477119
rect 256606 477048 256662 477057
rect 256606 476983 256662 476992
rect 242808 476672 242860 476678
rect 242808 476614 242860 476620
rect 253754 476504 253810 476513
rect 256620 476474 256648 476983
rect 253754 476439 253810 476448
rect 256608 476468 256660 476474
rect 245474 476368 245530 476377
rect 245474 476303 245530 476312
rect 248326 476368 248382 476377
rect 248326 476303 248382 476312
rect 251086 476368 251142 476377
rect 251086 476303 251142 476312
rect 252374 476368 252430 476377
rect 252374 476303 252430 476312
rect 244186 476232 244242 476241
rect 244186 476167 244242 476176
rect 240048 476128 240100 476134
rect 240048 476070 240100 476076
rect 239404 460420 239456 460426
rect 239404 460362 239456 460368
rect 244200 454850 244228 476167
rect 244188 454844 244240 454850
rect 244188 454786 244240 454792
rect 245488 449750 245516 476303
rect 245566 476232 245622 476241
rect 245566 476167 245622 476176
rect 246946 476232 247002 476241
rect 246946 476167 247002 476176
rect 248234 476232 248290 476241
rect 248234 476167 248290 476176
rect 245476 449744 245528 449750
rect 245476 449686 245528 449692
rect 245580 449682 245608 476167
rect 246960 464506 246988 476167
rect 248248 470082 248276 476167
rect 248236 470076 248288 470082
rect 248236 470018 248288 470024
rect 248340 467362 248368 476303
rect 249706 476232 249762 476241
rect 249706 476167 249762 476176
rect 250994 476232 251050 476241
rect 250994 476167 251050 476176
rect 248328 467356 248380 467362
rect 248328 467298 248380 467304
rect 246948 464500 247000 464506
rect 246948 464442 247000 464448
rect 249720 457638 249748 476167
rect 251008 460494 251036 476167
rect 250996 460488 251048 460494
rect 250996 460430 251048 460436
rect 249708 457632 249760 457638
rect 249708 457574 249760 457580
rect 251100 453558 251128 476303
rect 252388 463146 252416 476303
rect 252466 476232 252522 476241
rect 252466 476167 252522 476176
rect 252376 463140 252428 463146
rect 252376 463082 252428 463088
rect 252284 456816 252336 456822
rect 252284 456758 252336 456764
rect 251088 453552 251140 453558
rect 251088 453494 251140 453500
rect 245568 449676 245620 449682
rect 245568 449618 245620 449624
rect 237196 447976 237248 447982
rect 237196 447918 237248 447924
rect 250996 446004 251048 446010
rect 250996 445946 251048 445952
rect 249708 445936 249760 445942
rect 241794 445904 241850 445913
rect 235908 445868 235960 445874
rect 249708 445878 249760 445884
rect 241794 445839 241850 445848
rect 235908 445810 235960 445816
rect 231124 444984 231176 444990
rect 231124 444926 231176 444932
rect 225604 444916 225656 444922
rect 225604 444858 225656 444864
rect 219348 443760 219400 443766
rect 219348 443702 219400 443708
rect 217784 443692 217836 443698
rect 217784 443634 217836 443640
rect 224224 372768 224276 372774
rect 224224 372710 224276 372716
rect 220084 346452 220136 346458
rect 220084 346394 220136 346400
rect 216586 308408 216642 308417
rect 216586 308343 216642 308352
rect 216496 306264 216548 306270
rect 216496 306206 216548 306212
rect 216312 305924 216364 305930
rect 216312 305866 216364 305872
rect 216220 303272 216272 303278
rect 216220 303214 216272 303220
rect 216128 302796 216180 302802
rect 216128 302738 216180 302744
rect 216036 297220 216088 297226
rect 216036 297162 216088 297168
rect 215944 215280 215996 215286
rect 215944 215222 215996 215228
rect 215944 213920 215996 213926
rect 215944 213862 215996 213868
rect 215852 159384 215904 159390
rect 215852 159326 215904 159332
rect 215956 3670 215984 213862
rect 216048 155718 216076 297162
rect 216140 157962 216168 302738
rect 216232 158234 216260 303214
rect 216220 158228 216272 158234
rect 216220 158170 216272 158176
rect 216324 158030 216352 305866
rect 216404 303544 216456 303550
rect 216404 303486 216456 303492
rect 216312 158024 216364 158030
rect 216312 157966 216364 157972
rect 216128 157956 216180 157962
rect 216128 157898 216180 157904
rect 216036 155712 216088 155718
rect 216036 155654 216088 155660
rect 216416 4146 216444 303486
rect 216404 4140 216456 4146
rect 216404 4082 216456 4088
rect 215944 3664 215996 3670
rect 215944 3606 215996 3612
rect 215666 3496 215722 3505
rect 215666 3431 215722 3440
rect 215208 3324 215260 3330
rect 215208 3266 215260 3272
rect 215680 480 215708 3431
rect 216508 3262 216536 306206
rect 216600 3602 216628 308343
rect 220096 307494 220124 346394
rect 224236 308446 224264 372710
rect 224224 308440 224276 308446
rect 224224 308382 224276 308388
rect 220084 307488 220136 307494
rect 220084 307430 220136 307436
rect 219072 306332 219124 306338
rect 219072 306274 219124 306280
rect 218980 305584 219032 305590
rect 218980 305526 219032 305532
rect 218888 305516 218940 305522
rect 218888 305458 218940 305464
rect 217968 303612 218020 303618
rect 217968 303554 218020 303560
rect 217876 295316 217928 295322
rect 217876 295258 217928 295264
rect 217692 290692 217744 290698
rect 217692 290634 217744 290640
rect 217600 283824 217652 283830
rect 217600 283766 217652 283772
rect 217508 258732 217560 258738
rect 217508 258674 217560 258680
rect 217232 256284 217284 256290
rect 217232 256226 217284 256232
rect 217140 253496 217192 253502
rect 217140 253438 217192 253444
rect 217152 192817 217180 253438
rect 217244 195945 217272 256226
rect 217324 246764 217376 246770
rect 217324 246706 217376 246712
rect 217230 195936 217286 195945
rect 217230 195871 217286 195880
rect 217138 192808 217194 192817
rect 217138 192743 217194 192752
rect 217336 168065 217364 246706
rect 217416 243568 217468 243574
rect 217416 243510 217468 243516
rect 217322 168056 217378 168065
rect 217322 167991 217378 168000
rect 217428 155106 217456 243510
rect 217520 169969 217548 258674
rect 217612 193769 217640 283766
rect 217704 196897 217732 290634
rect 217784 261656 217836 261662
rect 217784 261598 217836 261604
rect 217690 196888 217746 196897
rect 217690 196823 217746 196832
rect 217692 195424 217744 195430
rect 217692 195366 217744 195372
rect 217598 193760 217654 193769
rect 217598 193695 217654 193704
rect 217506 169960 217562 169969
rect 217506 169895 217562 169904
rect 217704 155174 217732 195366
rect 217796 168337 217824 261598
rect 217782 168328 217838 168337
rect 217782 168263 217838 168272
rect 217692 155168 217744 155174
rect 217692 155110 217744 155116
rect 217416 155100 217468 155106
rect 217416 155042 217468 155048
rect 217888 155038 217916 295258
rect 217980 158166 218008 303554
rect 218796 294500 218848 294506
rect 218796 294442 218848 294448
rect 218704 293480 218756 293486
rect 218704 293422 218756 293428
rect 218612 267232 218664 267238
rect 218612 267174 218664 267180
rect 218428 256352 218480 256358
rect 218428 256294 218480 256300
rect 218440 243545 218468 256294
rect 218520 252068 218572 252074
rect 218520 252010 218572 252016
rect 218426 243536 218482 243545
rect 218426 243471 218482 243480
rect 218532 189961 218560 252010
rect 218518 189952 218574 189961
rect 218518 189887 218574 189896
rect 218624 188193 218652 267174
rect 218716 191049 218744 293422
rect 218702 191040 218758 191049
rect 218702 190975 218758 190984
rect 218610 188184 218666 188193
rect 218610 188119 218666 188128
rect 217968 158160 218020 158166
rect 217968 158102 218020 158108
rect 218808 155310 218836 294442
rect 218900 158273 218928 305458
rect 218886 158264 218942 158273
rect 218886 158199 218942 158208
rect 218992 157894 219020 305526
rect 219084 158438 219112 306274
rect 219164 306060 219216 306066
rect 219164 306002 219216 306008
rect 219072 158432 219124 158438
rect 219072 158374 219124 158380
rect 219176 158098 219204 306002
rect 219256 303340 219308 303346
rect 219256 303282 219308 303288
rect 219164 158092 219216 158098
rect 219164 158034 219216 158040
rect 218980 157888 219032 157894
rect 218980 157830 219032 157836
rect 219268 155446 219296 303282
rect 225616 267714 225644 444858
rect 230480 443828 230532 443834
rect 230480 443770 230532 443776
rect 229744 443488 229796 443494
rect 229744 443430 229796 443436
rect 228364 443420 228416 443426
rect 228364 443362 228416 443368
rect 225696 374808 225748 374814
rect 225696 374750 225748 374756
rect 225708 310593 225736 374750
rect 226984 374468 227036 374474
rect 226984 374410 227036 374416
rect 225788 328500 225840 328506
rect 225788 328442 225840 328448
rect 225694 310584 225750 310593
rect 225694 310519 225750 310528
rect 225800 307698 225828 328442
rect 226996 310554 227024 374410
rect 227076 368552 227128 368558
rect 227076 368494 227128 368500
rect 226984 310548 227036 310554
rect 226984 310490 227036 310496
rect 227088 309641 227116 368494
rect 227168 351960 227220 351966
rect 227168 351902 227220 351908
rect 227074 309632 227130 309641
rect 227074 309567 227130 309576
rect 227180 307766 227208 351902
rect 227168 307760 227220 307766
rect 227168 307702 227220 307708
rect 225788 307692 225840 307698
rect 225788 307634 225840 307640
rect 228376 293962 228404 443362
rect 229756 376038 229784 443430
rect 230492 438190 230520 443770
rect 230480 438184 230532 438190
rect 230480 438126 230532 438132
rect 231136 398818 231164 444926
rect 234618 444680 234674 444689
rect 234618 444615 234674 444624
rect 233974 443456 234030 443465
rect 233974 443391 234030 443400
rect 232686 443184 232742 443193
rect 232686 443119 232742 443128
rect 231216 442196 231268 442202
rect 231216 442138 231268 442144
rect 231228 411262 231256 442138
rect 232700 441524 232728 443119
rect 233330 443048 233386 443057
rect 233330 442983 233386 442992
rect 233344 441524 233372 442983
rect 233988 441524 234016 443391
rect 234632 441524 234660 444615
rect 235264 443012 235316 443018
rect 235264 442954 235316 442960
rect 235276 441524 235304 442954
rect 235920 441524 235948 445810
rect 237838 445768 237894 445777
rect 237838 445703 237894 445712
rect 236550 444408 236606 444417
rect 236550 444343 236606 444352
rect 236564 441524 236592 444343
rect 237196 443148 237248 443154
rect 237196 443090 237248 443096
rect 237208 441524 237236 443090
rect 237852 441524 237880 445703
rect 240508 444712 240560 444718
rect 240508 444654 240560 444660
rect 238574 444544 238630 444553
rect 238574 444479 238630 444488
rect 238588 441524 238616 444479
rect 239220 443352 239272 443358
rect 239220 443294 239272 443300
rect 239862 443320 239918 443329
rect 239232 441524 239260 443294
rect 239862 443255 239918 443264
rect 239876 441524 239904 443255
rect 240520 441524 240548 444654
rect 241152 441652 241204 441658
rect 241152 441594 241204 441600
rect 241164 441524 241192 441594
rect 241808 441524 241836 445839
rect 245752 444780 245804 444786
rect 245752 444722 245804 444728
rect 244464 444440 244516 444446
rect 244464 444382 244516 444388
rect 243084 443964 243136 443970
rect 243084 443906 243136 443912
rect 242900 443012 242952 443018
rect 242900 442954 242952 442960
rect 242912 442270 242940 442954
rect 242900 442264 242952 442270
rect 242900 442206 242952 442212
rect 243096 441524 243124 443906
rect 243728 443624 243780 443630
rect 243728 443566 243780 443572
rect 243740 441524 243768 443566
rect 244476 441524 244504 444382
rect 245108 444100 245160 444106
rect 245108 444042 245160 444048
rect 245120 441524 245148 444042
rect 245568 443148 245620 443154
rect 245568 443090 245620 443096
rect 245580 442338 245608 443090
rect 245568 442332 245620 442338
rect 245568 442274 245620 442280
rect 245764 441524 245792 444722
rect 248328 444168 248380 444174
rect 248328 444110 248380 444116
rect 246396 443012 246448 443018
rect 246396 442954 246448 442960
rect 246408 441524 246436 442954
rect 247040 441788 247092 441794
rect 247040 441730 247092 441736
rect 247052 441524 247080 441730
rect 248340 441524 248368 444110
rect 248972 441924 249024 441930
rect 248972 441866 249024 441872
rect 248984 441524 249012 441866
rect 249720 441524 249748 445878
rect 250352 443216 250404 443222
rect 250352 443158 250404 443164
rect 250364 441524 250392 443158
rect 251008 441524 251036 445946
rect 251180 443964 251232 443970
rect 251180 443906 251232 443912
rect 251192 442406 251220 443906
rect 251272 443556 251324 443562
rect 251272 443498 251324 443504
rect 251180 442400 251232 442406
rect 251180 442342 251232 442348
rect 242348 441176 242400 441182
rect 242348 441118 242400 441124
rect 248052 441176 248104 441182
rect 248052 441118 248104 441124
rect 242360 441046 242388 441118
rect 248064 441046 248092 441118
rect 251284 441114 251312 443498
rect 252296 441524 252324 456758
rect 252480 452198 252508 476167
rect 252928 474088 252980 474094
rect 252928 474030 252980 474036
rect 252468 452192 252520 452198
rect 252468 452134 252520 452140
rect 252940 441524 252968 474030
rect 253768 472870 253796 476439
rect 256608 476410 256660 476416
rect 253846 476232 253902 476241
rect 253846 476167 253902 476176
rect 255226 476232 255282 476241
rect 255226 476167 255282 476176
rect 256514 476232 256570 476241
rect 256514 476167 256570 476176
rect 253756 472864 253808 472870
rect 253756 472806 253808 472812
rect 253572 470620 253624 470626
rect 253572 470562 253624 470568
rect 253584 441524 253612 470562
rect 253860 468790 253888 476167
rect 254860 472728 254912 472734
rect 254860 472670 254912 472676
rect 253848 468784 253900 468790
rect 253848 468726 253900 468732
rect 254216 450696 254268 450702
rect 254216 450638 254268 450644
rect 254228 441524 254256 450638
rect 254872 441524 254900 472670
rect 255240 463078 255268 476167
rect 255596 475380 255648 475386
rect 255596 475322 255648 475328
rect 255228 463072 255280 463078
rect 255228 463014 255280 463020
rect 255608 441524 255636 475322
rect 256528 457570 256556 476167
rect 256516 457564 256568 457570
rect 256516 457506 256568 457512
rect 255964 451988 256016 451994
rect 255964 451930 256016 451936
rect 255976 441862 256004 451930
rect 255964 441856 256016 441862
rect 255964 441798 256016 441804
rect 255976 441538 256004 441798
rect 255976 441510 256266 441538
rect 256896 441524 256924 478178
rect 259366 476776 259422 476785
rect 259366 476711 259422 476720
rect 264794 476776 264850 476785
rect 264794 476711 264850 476720
rect 257986 476232 258042 476241
rect 257986 476167 258042 476176
rect 259274 476232 259330 476241
rect 259274 476167 259330 476176
rect 258000 470014 258028 476167
rect 259288 471442 259316 476167
rect 259276 471436 259328 471442
rect 259276 471378 259328 471384
rect 257988 470008 258040 470014
rect 257988 469950 258040 469956
rect 257528 469940 257580 469946
rect 257528 469882 257580 469888
rect 257540 441524 257568 469882
rect 258816 465792 258868 465798
rect 258816 465734 258868 465740
rect 258172 453348 258224 453354
rect 258172 453290 258224 453296
rect 258184 441524 258212 453290
rect 258828 441524 258856 465734
rect 259380 456210 259408 476711
rect 262126 476504 262182 476513
rect 262126 476439 262182 476448
rect 262140 476406 262168 476439
rect 262128 476400 262180 476406
rect 260746 476368 260802 476377
rect 262128 476342 262180 476348
rect 260746 476303 260802 476312
rect 260654 476232 260710 476241
rect 260654 476167 260710 476176
rect 260668 458998 260696 476167
rect 260656 458992 260708 458998
rect 260656 458934 260708 458940
rect 259368 456204 259420 456210
rect 259368 456146 259420 456152
rect 260104 454776 260156 454782
rect 260104 454718 260156 454724
rect 259460 446412 259512 446418
rect 259460 446354 259512 446360
rect 259472 443834 259500 446354
rect 259460 443828 259512 443834
rect 259460 443770 259512 443776
rect 259472 441524 259500 443770
rect 260116 441524 260144 454718
rect 260760 447914 260788 476303
rect 262034 476232 262090 476241
rect 262034 476167 262090 476176
rect 263506 476232 263562 476241
rect 263506 476167 263562 476176
rect 260840 463004 260892 463010
rect 260840 462946 260892 462952
rect 260748 447908 260800 447914
rect 260748 447850 260800 447856
rect 260852 441524 260880 462946
rect 262048 461786 262076 476167
rect 262772 467220 262824 467226
rect 262772 467162 262824 467168
rect 262036 461780 262088 461786
rect 262036 461722 262088 461728
rect 262128 456136 262180 456142
rect 262128 456078 262180 456084
rect 261484 450628 261536 450634
rect 261484 450570 261536 450576
rect 261496 441524 261524 450570
rect 262140 441524 262168 456078
rect 262784 441524 262812 467162
rect 263520 449478 263548 476167
rect 264808 474298 264836 476711
rect 266266 476640 266322 476649
rect 266266 476575 266322 476584
rect 266280 476542 266308 476575
rect 266268 476536 266320 476542
rect 266268 476478 266320 476484
rect 267646 476368 267702 476377
rect 267646 476303 267702 476312
rect 264886 476232 264942 476241
rect 264886 476167 264942 476176
rect 266174 476232 266230 476241
rect 266174 476167 266230 476176
rect 267554 476232 267610 476241
rect 267554 476167 267610 476176
rect 264796 474292 264848 474298
rect 264796 474234 264848 474240
rect 264704 468580 264756 468586
rect 264704 468522 264756 468528
rect 264060 458856 264112 458862
rect 264060 458798 264112 458804
rect 263508 449472 263560 449478
rect 263508 449414 263560 449420
rect 263416 446548 263468 446554
rect 263416 446490 263468 446496
rect 263428 441524 263456 446490
rect 264072 441524 264100 458798
rect 264716 441524 264744 468522
rect 264900 449410 264928 476167
rect 265992 460284 266044 460290
rect 265992 460226 266044 460232
rect 264888 449404 264940 449410
rect 264888 449346 264940 449352
rect 265348 446616 265400 446622
rect 265348 446558 265400 446564
rect 265360 441524 265388 446558
rect 266004 441524 266032 460226
rect 266188 449546 266216 476167
rect 266728 464364 266780 464370
rect 266728 464306 266780 464312
rect 266176 449540 266228 449546
rect 266176 449482 266228 449488
rect 266740 441524 266768 464306
rect 267568 449206 267596 476167
rect 267660 449614 267688 476303
rect 268016 461712 268068 461718
rect 268016 461654 268068 461660
rect 267648 449608 267700 449614
rect 267648 449550 267700 449556
rect 267556 449200 267608 449206
rect 267556 449142 267608 449148
rect 267372 446684 267424 446690
rect 267372 446626 267424 446632
rect 267384 441524 267412 446626
rect 268028 441524 268056 461654
rect 268672 441524 268700 478450
rect 269304 478440 269356 478446
rect 269304 478382 269356 478388
rect 268934 476368 268990 476377
rect 268934 476303 268990 476312
rect 268948 454918 268976 476303
rect 269026 476232 269082 476241
rect 269026 476167 269082 476176
rect 268936 454912 268988 454918
rect 268936 454854 268988 454860
rect 269040 449342 269068 476167
rect 269028 449336 269080 449342
rect 269028 449278 269080 449284
rect 269316 441524 269344 478382
rect 269960 441524 269988 478586
rect 271236 478576 271288 478582
rect 271236 478518 271288 478524
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 270420 449274 270448 476167
rect 270408 449268 270460 449274
rect 270408 449210 270460 449216
rect 270592 443760 270644 443766
rect 270592 443702 270644 443708
rect 270604 441524 270632 443702
rect 271248 441524 271276 478518
rect 357452 478514 357480 700266
rect 358084 510672 358136 510678
rect 358084 510614 358136 510620
rect 357440 478508 357492 478514
rect 357440 478450 357492 478456
rect 308588 478372 308640 478378
rect 308588 478314 308640 478320
rect 282368 478168 282420 478174
rect 282368 478110 282420 478116
rect 271786 476640 271842 476649
rect 271786 476575 271788 476584
rect 271840 476575 271842 476584
rect 271788 476546 271840 476552
rect 274454 476504 274510 476513
rect 274454 476439 274510 476448
rect 271694 476232 271750 476241
rect 271694 476167 271750 476176
rect 273166 476232 273222 476241
rect 273166 476167 273222 476176
rect 274362 476232 274418 476241
rect 274362 476167 274418 476176
rect 271708 453490 271736 476167
rect 272616 456272 272668 456278
rect 272616 456214 272668 456220
rect 271696 453484 271748 453490
rect 271696 453426 271748 453432
rect 271972 443692 272024 443698
rect 271972 443634 272024 443640
rect 271984 441524 272012 443634
rect 272628 441524 272656 456214
rect 273180 452062 273208 476167
rect 274376 464438 274404 476167
rect 274468 474230 274496 476439
rect 274546 476368 274602 476377
rect 274546 476303 274602 476312
rect 277306 476368 277362 476377
rect 277306 476303 277362 476312
rect 278594 476368 278650 476377
rect 278594 476303 278650 476312
rect 274560 475522 274588 476303
rect 275926 476232 275982 476241
rect 275926 476167 275982 476176
rect 277214 476232 277270 476241
rect 277214 476167 277270 476176
rect 274548 475516 274600 475522
rect 274548 475458 274600 475464
rect 274456 474224 274508 474230
rect 274456 474166 274508 474172
rect 275192 474020 275244 474026
rect 275192 473962 275244 473968
rect 273260 464432 273312 464438
rect 273260 464374 273312 464380
rect 274364 464432 274416 464438
rect 274364 464374 274416 464380
rect 273168 452056 273220 452062
rect 273168 451998 273220 452004
rect 273272 441524 273300 464374
rect 274548 458924 274600 458930
rect 274548 458866 274600 458872
rect 273904 453416 273956 453422
rect 273904 453358 273956 453364
rect 273916 441524 273944 453358
rect 274560 441524 274588 458866
rect 275204 441524 275232 473962
rect 275940 465934 275968 476167
rect 275928 465928 275980 465934
rect 275928 465870 275980 465876
rect 276480 461644 276532 461650
rect 276480 461586 276532 461592
rect 275836 451920 275888 451926
rect 275836 451862 275888 451868
rect 275848 441524 275876 451862
rect 276112 443624 276164 443630
rect 276112 443566 276164 443572
rect 276020 443080 276072 443086
rect 276020 443022 276072 443028
rect 276032 442542 276060 443022
rect 276020 442536 276072 442542
rect 276020 442478 276072 442484
rect 276124 442474 276152 443566
rect 276112 442468 276164 442474
rect 276112 442410 276164 442416
rect 276492 441524 276520 461586
rect 277228 460358 277256 476167
rect 277216 460352 277268 460358
rect 277216 460294 277268 460300
rect 277320 456074 277348 476303
rect 278504 460216 278556 460222
rect 278504 460158 278556 460164
rect 277124 456068 277176 456074
rect 277124 456010 277176 456016
rect 277308 456068 277360 456074
rect 277308 456010 277360 456016
rect 277136 441524 277164 456010
rect 277860 454708 277912 454714
rect 277860 454650 277912 454656
rect 277400 443012 277452 443018
rect 277400 442954 277452 442960
rect 251272 441108 251324 441114
rect 251272 441050 251324 441056
rect 277412 441046 277440 442954
rect 277872 441524 277900 454650
rect 278516 441524 278544 460158
rect 278608 454714 278636 476303
rect 278686 476232 278742 476241
rect 278686 476167 278742 476176
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 281446 476232 281502 476241
rect 281446 476167 281502 476176
rect 278596 454708 278648 454714
rect 278596 454650 278648 454656
rect 278700 450770 278728 476167
rect 280080 468722 280108 476167
rect 280068 468716 280120 468722
rect 280068 468658 280120 468664
rect 279792 465724 279844 465730
rect 279792 465666 279844 465672
rect 278688 450764 278740 450770
rect 278688 450706 278740 450712
rect 279148 450560 279200 450566
rect 279148 450502 279200 450508
rect 279160 441524 279188 450502
rect 279804 441524 279832 465666
rect 281080 459060 281132 459066
rect 281080 459002 281132 459008
rect 280436 457496 280488 457502
rect 280436 457438 280488 457444
rect 279974 443456 280030 443465
rect 279974 443391 280030 443400
rect 279988 442542 280016 443391
rect 280068 443012 280120 443018
rect 280068 442954 280120 442960
rect 280080 442610 280108 442954
rect 280068 442604 280120 442610
rect 280068 442546 280120 442552
rect 279976 442536 280028 442542
rect 279976 442478 280028 442484
rect 280448 441524 280476 457438
rect 281092 441524 281120 459002
rect 281460 458930 281488 476167
rect 281724 467152 281776 467158
rect 281724 467094 281776 467100
rect 281448 458924 281500 458930
rect 281448 458866 281500 458872
rect 281736 441524 281764 467094
rect 282380 441524 282408 478110
rect 284206 476232 284262 476241
rect 284206 476167 284262 476176
rect 286506 476232 286562 476241
rect 286506 476167 286562 476176
rect 288346 476232 288402 476241
rect 288346 476167 288402 476176
rect 291106 476232 291162 476241
rect 291106 476167 291162 476176
rect 293866 476232 293922 476241
rect 293866 476167 293922 476176
rect 296626 476232 296682 476241
rect 296626 476167 296682 476176
rect 299386 476232 299442 476241
rect 299386 476167 299442 476176
rect 302146 476232 302202 476241
rect 302146 476167 302202 476176
rect 303526 476232 303582 476241
rect 303526 476167 303582 476176
rect 306286 476232 306342 476241
rect 306286 476167 306342 476176
rect 283748 468512 283800 468518
rect 283748 468454 283800 468460
rect 283012 453620 283064 453626
rect 283012 453562 283064 453568
rect 283024 441524 283052 453562
rect 283760 441524 283788 468454
rect 284220 448050 284248 476167
rect 284392 472660 284444 472666
rect 284392 472602 284444 472608
rect 284208 448044 284260 448050
rect 284208 447986 284260 447992
rect 284404 441524 284432 472602
rect 286520 471306 286548 476167
rect 287612 474768 287664 474774
rect 287612 474710 287664 474716
rect 286324 471300 286376 471306
rect 286324 471242 286376 471248
rect 286508 471300 286560 471306
rect 286508 471242 286560 471248
rect 285680 469872 285732 469878
rect 285680 469814 285732 469820
rect 285036 461848 285088 461854
rect 285036 461790 285088 461796
rect 285048 441524 285076 461790
rect 285692 441524 285720 469814
rect 286336 441524 286364 471242
rect 286968 452124 287020 452130
rect 286968 452066 287020 452072
rect 286980 441524 287008 452066
rect 287624 441524 287652 474710
rect 288360 461650 288388 476167
rect 291120 465730 291148 476167
rect 293880 469878 293908 476167
rect 294604 471436 294656 471442
rect 294604 471378 294656 471384
rect 293868 469872 293920 469878
rect 293868 469814 293920 469820
rect 291108 465724 291160 465730
rect 291108 465666 291160 465672
rect 288992 462392 289044 462398
rect 288992 462334 289044 462340
rect 288348 461644 288400 461650
rect 288348 461586 288400 461592
rect 288256 446480 288308 446486
rect 288256 446422 288308 446428
rect 288268 441524 288296 446422
rect 289004 441524 289032 462334
rect 293224 454912 293276 454918
rect 293224 454854 293276 454860
rect 290280 444984 290332 444990
rect 290280 444926 290332 444932
rect 289636 444508 289688 444514
rect 289636 444450 289688 444456
rect 289648 441524 289676 444450
rect 290292 441524 290320 444926
rect 291568 444644 291620 444650
rect 291568 444586 291620 444592
rect 290924 442196 290976 442202
rect 290924 442138 290976 442144
rect 290936 441524 290964 442138
rect 291580 441524 291608 444586
rect 293236 443698 293264 454854
rect 293500 444576 293552 444582
rect 293500 444518 293552 444524
rect 293224 443692 293276 443698
rect 293224 443634 293276 443640
rect 292856 443488 292908 443494
rect 292856 443430 292908 443436
rect 292212 443080 292264 443086
rect 292212 443022 292264 443028
rect 292224 441524 292252 443022
rect 292868 441524 292896 443430
rect 293512 441524 293540 444518
rect 294616 443834 294644 471378
rect 296640 454918 296668 476167
rect 297364 474292 297416 474298
rect 297364 474234 297416 474240
rect 296628 454912 296680 454918
rect 296628 454854 296680 454860
rect 295524 444916 295576 444922
rect 295524 444858 295576 444864
rect 294880 443896 294932 443902
rect 294880 443838 294932 443844
rect 294604 443828 294656 443834
rect 294604 443770 294656 443776
rect 294144 443420 294196 443426
rect 294144 443362 294196 443368
rect 294156 441524 294184 443362
rect 294892 441524 294920 443838
rect 295536 441524 295564 444858
rect 297376 443766 297404 474234
rect 299400 467158 299428 476167
rect 302160 472666 302188 476167
rect 302148 472660 302200 472666
rect 302148 472602 302200 472608
rect 301504 468784 301556 468790
rect 301504 468726 301556 468732
rect 299388 467152 299440 467158
rect 299388 467094 299440 467100
rect 300124 446208 300176 446214
rect 300124 446150 300176 446156
rect 297456 444848 297508 444854
rect 297456 444790 297508 444796
rect 299386 444816 299442 444825
rect 297364 443760 297416 443766
rect 297364 443702 297416 443708
rect 296168 443012 296220 443018
rect 296168 442954 296220 442960
rect 296180 441524 296208 442954
rect 296812 441720 296864 441726
rect 296812 441662 296864 441668
rect 296824 441524 296852 441662
rect 297468 441524 297496 444790
rect 299386 444751 299442 444760
rect 298744 443284 298796 443290
rect 298744 443226 298796 443232
rect 298098 441688 298154 441697
rect 298098 441623 298154 441632
rect 298112 441524 298140 441623
rect 298756 441524 298784 443226
rect 299400 441524 299428 444751
rect 300136 441524 300164 446150
rect 300768 446140 300820 446146
rect 300768 446082 300820 446088
rect 300780 441524 300808 446082
rect 301516 443902 301544 468726
rect 303540 448118 303568 476167
rect 306300 457502 306328 476167
rect 307300 465860 307352 465866
rect 307300 465802 307352 465808
rect 306288 457496 306340 457502
rect 306288 457438 306340 457444
rect 303528 448112 303580 448118
rect 303528 448054 303580 448060
rect 306012 446072 306064 446078
rect 306012 446014 306064 446020
rect 303988 445800 304040 445806
rect 303988 445742 304040 445748
rect 301504 443896 301556 443902
rect 301504 443838 301556 443844
rect 301412 443556 301464 443562
rect 301412 443498 301464 443504
rect 300858 443320 300914 443329
rect 300858 443255 300914 443264
rect 300872 442610 300900 443255
rect 300860 442604 300912 442610
rect 300860 442546 300912 442552
rect 301424 441524 301452 443498
rect 302056 442128 302108 442134
rect 302056 442070 302108 442076
rect 302068 441524 302096 442070
rect 302700 442060 302752 442066
rect 302700 442002 302752 442008
rect 302712 441524 302740 442002
rect 304000 441524 304028 445742
rect 306024 441524 306052 446014
rect 306656 441992 306708 441998
rect 306656 441934 306708 441940
rect 306668 441524 306696 441934
rect 307312 441524 307340 465802
rect 307944 447840 307996 447846
rect 307944 447782 307996 447788
rect 307956 441524 307984 447782
rect 308600 441524 308628 478314
rect 314476 478304 314528 478310
rect 314476 478246 314528 478252
rect 309046 476776 309102 476785
rect 309046 476711 309102 476720
rect 311256 476740 311308 476746
rect 309060 476338 309088 476711
rect 311256 476682 311308 476688
rect 309048 476332 309100 476338
rect 309048 476274 309100 476280
rect 310520 470076 310572 470082
rect 310520 470018 310572 470024
rect 309232 460420 309284 460426
rect 309232 460362 309284 460368
rect 309244 441524 309272 460362
rect 309876 454844 309928 454850
rect 309876 454786 309928 454792
rect 309888 441524 309916 454786
rect 310532 441524 310560 470018
rect 311268 441524 311296 476682
rect 311806 476368 311862 476377
rect 311806 476303 311862 476312
rect 311820 476270 311848 476303
rect 311808 476264 311860 476270
rect 311808 476206 311860 476212
rect 313832 476128 313884 476134
rect 313832 476070 313884 476076
rect 313188 460488 313240 460494
rect 313188 460430 313240 460436
rect 312544 449744 312596 449750
rect 312544 449686 312596 449692
rect 311900 447976 311952 447982
rect 311900 447918 311952 447924
rect 311912 441524 311940 447918
rect 312556 441524 312584 449686
rect 313200 441524 313228 460430
rect 313844 441524 313872 476070
rect 314488 441524 314516 478246
rect 316408 476808 316460 476814
rect 314566 476776 314622 476785
rect 316408 476750 316460 476756
rect 314566 476711 314622 476720
rect 314580 476134 314608 476711
rect 315946 476232 316002 476241
rect 315946 476167 315948 476176
rect 316000 476167 316002 476176
rect 315948 476138 316000 476144
rect 314568 476128 314620 476134
rect 314568 476070 314620 476076
rect 315120 449676 315172 449682
rect 315120 449618 315172 449624
rect 315132 441524 315160 449618
rect 315764 443896 315816 443902
rect 315764 443838 315816 443844
rect 315776 441524 315804 443838
rect 316420 441524 316448 476750
rect 319076 476672 319128 476678
rect 319076 476614 319128 476620
rect 318706 476504 318762 476513
rect 318432 476468 318484 476474
rect 318706 476439 318708 476448
rect 318432 476410 318484 476416
rect 318760 476439 318762 476448
rect 318708 476410 318760 476416
rect 317144 474156 317196 474162
rect 317144 474098 317196 474104
rect 317156 441524 317184 474098
rect 317788 464500 317840 464506
rect 317788 464442 317840 464448
rect 317800 441524 317828 464442
rect 318444 441524 318472 476410
rect 319088 441524 319116 476614
rect 330208 476604 330260 476610
rect 330208 476546 330260 476552
rect 326896 476536 326948 476542
rect 326896 476478 326948 476484
rect 326986 476504 327042 476513
rect 323032 476400 323084 476406
rect 323032 476342 323084 476348
rect 321466 476232 321522 476241
rect 321466 476167 321522 476176
rect 321480 475590 321508 476167
rect 321468 475584 321520 475590
rect 321468 475526 321520 475532
rect 321652 475448 321704 475454
rect 321652 475390 321704 475396
rect 319720 468648 319772 468654
rect 319720 468590 319772 468596
rect 319732 441524 319760 468590
rect 320364 467356 320416 467362
rect 320364 467298 320416 467304
rect 320376 441524 320404 467298
rect 321008 443828 321060 443834
rect 321008 443770 321060 443776
rect 321020 441524 321048 443770
rect 321664 441524 321692 475390
rect 322296 457632 322348 457638
rect 322296 457574 322348 457580
rect 322308 441524 322336 457574
rect 323044 441524 323072 476342
rect 324226 476232 324282 476241
rect 324226 476167 324282 476176
rect 323676 472796 323728 472802
rect 323676 472738 323728 472744
rect 323688 441524 323716 472738
rect 324240 463214 324268 476167
rect 325608 467288 325660 467294
rect 325608 467230 325660 467236
rect 324228 463208 324280 463214
rect 324228 463150 324280 463156
rect 324320 453552 324372 453558
rect 324320 453494 324372 453500
rect 324332 441524 324360 453494
rect 324964 443760 325016 443766
rect 324964 443702 325016 443708
rect 324976 441524 325004 443702
rect 325620 441524 325648 467230
rect 326252 463140 326304 463146
rect 326252 463082 326304 463088
rect 326264 441524 326292 463082
rect 326908 441524 326936 476478
rect 326986 476439 327042 476448
rect 327000 476406 327028 476439
rect 326988 476400 327040 476406
rect 326988 476342 327040 476348
rect 329104 476332 329156 476338
rect 329104 476274 329156 476280
rect 327540 471368 327592 471374
rect 327540 471310 327592 471316
rect 327552 441524 327580 471310
rect 328276 452192 328328 452198
rect 328276 452134 328328 452140
rect 328288 441524 328316 452134
rect 329116 443766 329144 476274
rect 329564 472864 329616 472870
rect 329564 472806 329616 472812
rect 329104 443760 329156 443766
rect 329104 443702 329156 443708
rect 328920 443692 328972 443698
rect 328920 443634 328972 443640
rect 328932 441524 328960 443634
rect 329576 441524 329604 472806
rect 329748 443352 329800 443358
rect 329748 443294 329800 443300
rect 329760 442678 329788 443294
rect 329748 442672 329800 442678
rect 329748 442614 329800 442620
rect 330220 441524 330248 476546
rect 336004 476468 336056 476474
rect 336004 476410 336056 476416
rect 331864 476264 331916 476270
rect 331864 476206 331916 476212
rect 331496 475516 331548 475522
rect 331496 475458 331548 475464
rect 330852 463072 330904 463078
rect 330852 463014 330904 463020
rect 330864 441524 330892 463014
rect 331508 441524 331536 475458
rect 331876 443902 331904 476206
rect 334624 476196 334676 476202
rect 334624 476138 334676 476144
rect 333244 476128 333296 476134
rect 333244 476070 333296 476076
rect 332140 457564 332192 457570
rect 332140 457506 332192 457512
rect 331864 443896 331916 443902
rect 331864 443838 331916 443844
rect 332152 441524 332180 457506
rect 332784 456068 332836 456074
rect 332784 456010 332836 456016
rect 332796 441524 332824 456010
rect 333256 443970 333284 476070
rect 333428 470008 333480 470014
rect 333428 469950 333480 469956
rect 333244 443964 333296 443970
rect 333244 443906 333296 443912
rect 333440 441524 333468 469950
rect 334164 450764 334216 450770
rect 334164 450706 334216 450712
rect 334176 441524 334204 450706
rect 334636 444038 334664 476138
rect 335452 458924 335504 458930
rect 335452 458866 335504 458872
rect 334808 456204 334860 456210
rect 334808 456146 334860 456152
rect 334624 444032 334676 444038
rect 334624 443974 334676 443980
rect 334820 441524 334848 456146
rect 335464 441524 335492 458866
rect 336016 443834 336044 476410
rect 338764 476400 338816 476406
rect 338764 476342 338816 476348
rect 338028 471300 338080 471306
rect 338028 471242 338080 471248
rect 337384 458992 337436 458998
rect 337384 458934 337436 458940
rect 336740 448044 336792 448050
rect 336740 447986 336792 447992
rect 336096 447908 336148 447914
rect 336096 447850 336148 447856
rect 336004 443828 336056 443834
rect 336004 443770 336056 443776
rect 336108 441524 336136 447850
rect 336752 441524 336780 447986
rect 337396 441524 337424 458934
rect 338040 441524 338068 471242
rect 338672 461780 338724 461786
rect 338672 461722 338724 461728
rect 338684 441524 338712 461722
rect 338776 443698 338804 476342
rect 355324 475584 355376 475590
rect 355324 475526 355376 475532
rect 353116 474224 353168 474230
rect 353116 474166 353168 474172
rect 345940 472660 345992 472666
rect 345940 472602 345992 472608
rect 341984 469872 342036 469878
rect 341984 469814 342036 469820
rect 340696 465724 340748 465730
rect 340696 465666 340748 465672
rect 339408 461644 339460 461650
rect 339408 461586 339460 461592
rect 338764 443692 338816 443698
rect 338764 443634 338816 443640
rect 339420 441524 339448 461586
rect 340052 449472 340104 449478
rect 340052 449414 340104 449420
rect 340064 441524 340092 449414
rect 340708 441524 340736 465666
rect 341340 449404 341392 449410
rect 341340 449346 341392 449352
rect 341352 441524 341380 449346
rect 341996 441524 342024 469814
rect 344560 467152 344612 467158
rect 344560 467094 344612 467100
rect 343272 454912 343324 454918
rect 343272 454854 343324 454860
rect 342628 449540 342680 449546
rect 342628 449482 342680 449488
rect 342640 441524 342668 449482
rect 343284 441524 343312 454854
rect 343916 449608 343968 449614
rect 343916 449550 343968 449556
rect 343928 441524 343956 449550
rect 344572 441524 344600 467094
rect 345296 449200 345348 449206
rect 345296 449142 345348 449148
rect 345308 441524 345336 449142
rect 345952 441524 345980 472602
rect 351828 464432 351880 464438
rect 351828 464374 351880 464380
rect 348516 457496 348568 457502
rect 348516 457438 348568 457444
rect 346584 449336 346636 449342
rect 346584 449278 346636 449284
rect 346596 441524 346624 449278
rect 347872 449268 347924 449274
rect 347872 449210 347924 449216
rect 347228 448112 347280 448118
rect 347228 448054 347280 448060
rect 347240 441524 347268 448054
rect 347884 441524 347912 449210
rect 348528 441524 348556 457438
rect 349160 453484 349212 453490
rect 349160 453426 349212 453432
rect 349172 441524 349200 453426
rect 350540 452056 350592 452062
rect 350540 451998 350592 452004
rect 349804 443760 349856 443766
rect 349804 443702 349856 443708
rect 349816 441524 349844 443702
rect 350552 441524 350580 451998
rect 351184 443896 351236 443902
rect 351184 443838 351236 443844
rect 351196 441524 351224 443838
rect 351840 441524 351868 464374
rect 352472 443964 352524 443970
rect 352472 443906 352524 443912
rect 352484 441524 352512 443906
rect 353128 441524 353156 474166
rect 354404 465928 354456 465934
rect 354404 465870 354456 465876
rect 353760 444032 353812 444038
rect 353760 443974 353812 443980
rect 353772 441524 353800 443974
rect 354416 441524 354444 465870
rect 355336 444378 355364 475526
rect 356704 468716 356756 468722
rect 356704 468658 356756 468664
rect 355692 460352 355744 460358
rect 355692 460294 355744 460300
rect 355324 444372 355376 444378
rect 355324 444314 355376 444320
rect 355048 443828 355100 443834
rect 355048 443770 355100 443776
rect 355060 441524 355088 443770
rect 355704 441524 355732 460294
rect 356716 444378 356744 468658
rect 357716 463208 357768 463214
rect 357716 463150 357768 463156
rect 357072 454708 357124 454714
rect 357072 454650 357124 454656
rect 356428 444372 356480 444378
rect 356428 444314 356480 444320
rect 356704 444372 356756 444378
rect 356704 444314 356756 444320
rect 356440 441524 356468 444314
rect 357084 441524 357112 454650
rect 357728 441524 357756 463150
rect 358096 450702 358124 510614
rect 358832 478446 358860 700334
rect 359464 700324 359516 700330
rect 359464 700266 359516 700272
rect 358820 478440 358872 478446
rect 358820 478382 358872 478388
rect 359476 460290 359504 700266
rect 363604 616888 363656 616894
rect 363604 616830 363656 616836
rect 360844 484424 360896 484430
rect 360844 484366 360896 484372
rect 360856 474094 360884 484366
rect 360844 474088 360896 474094
rect 360844 474030 360896 474036
rect 359464 460284 359516 460290
rect 359464 460226 359516 460232
rect 363616 453354 363644 616830
rect 364352 461718 364380 702406
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 391204 696992 391256 696998
rect 391204 696934 391256 696940
rect 381544 683188 381596 683194
rect 381544 683130 381596 683136
rect 377404 670744 377456 670750
rect 377404 670686 377456 670692
rect 373264 643136 373316 643142
rect 373264 643078 373316 643084
rect 367744 563100 367796 563106
rect 367744 563042 367796 563048
rect 364340 461712 364392 461718
rect 364340 461654 364392 461660
rect 363604 453348 363656 453354
rect 363604 453290 363656 453296
rect 367756 451994 367784 563042
rect 369124 536852 369176 536858
rect 369124 536794 369176 536800
rect 369136 472734 369164 536794
rect 371884 524476 371936 524482
rect 371884 524418 371936 524424
rect 371896 475386 371924 524418
rect 371884 475380 371936 475386
rect 371884 475322 371936 475328
rect 369124 472728 369176 472734
rect 369124 472670 369176 472676
rect 373276 465798 373304 643078
rect 374644 590708 374696 590714
rect 374644 590650 374696 590656
rect 374656 478242 374684 590650
rect 374644 478236 374696 478242
rect 374644 478178 374696 478184
rect 373264 465792 373316 465798
rect 373264 465734 373316 465740
rect 377416 454782 377444 670686
rect 378784 576904 378836 576910
rect 378784 576846 378836 576852
rect 378796 469946 378824 576846
rect 378784 469940 378836 469946
rect 378784 469882 378836 469888
rect 377404 454776 377456 454782
rect 377404 454718 377456 454724
rect 367744 451988 367796 451994
rect 367744 451930 367796 451936
rect 358084 450696 358136 450702
rect 358084 450638 358136 450644
rect 381556 450634 381584 683130
rect 391216 463010 391244 696934
rect 396736 464370 396764 699654
rect 396724 464364 396776 464370
rect 396724 464306 396776 464312
rect 391204 463004 391256 463010
rect 391204 462946 391256 462952
rect 381544 450628 381596 450634
rect 381544 450570 381596 450576
rect 412652 446690 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 442264 700324 442316 700330
rect 442264 700266 442316 700272
rect 442276 456142 442304 700266
rect 462332 468586 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 468580 462372 468586
rect 462320 468522 462372 468528
rect 442264 456136 442316 456142
rect 442264 456078 442316 456084
rect 412640 446684 412692 446690
rect 412640 446626 412692 446632
rect 477512 446622 477540 702406
rect 494072 458862 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 467226 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 467220 527232 467226
rect 527180 467162 527232 467168
rect 494060 458856 494112 458862
rect 494060 458798 494112 458804
rect 477500 446616 477552 446622
rect 477500 446558 477552 446564
rect 542372 446554 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 542360 446548 542412 446554
rect 542360 446490 542412 446496
rect 580276 446418 580304 630799
rect 580264 446412 580316 446418
rect 580264 446354 580316 446360
rect 362592 446004 362644 446010
rect 362592 445946 362644 445952
rect 358360 444372 358412 444378
rect 358360 444314 358412 444320
rect 358372 441524 358400 444314
rect 362408 444168 362460 444174
rect 362408 444110 362460 444116
rect 362224 444100 362276 444106
rect 362224 444042 362276 444048
rect 359004 443692 359056 443698
rect 359004 443634 359056 443640
rect 359016 441524 359044 443634
rect 359648 443148 359700 443154
rect 359648 443090 359700 443096
rect 359660 441524 359688 443090
rect 360292 443080 360344 443086
rect 360292 443022 360344 443028
rect 360304 441524 360332 443022
rect 360936 443012 360988 443018
rect 360936 442954 360988 442960
rect 360948 441524 360976 442954
rect 289268 441448 289320 441454
rect 289268 441390 289320 441396
rect 284576 441380 284628 441386
rect 284576 441322 284628 441328
rect 283852 441250 284064 441266
rect 283840 441244 284076 441250
rect 283892 441238 284024 441244
rect 283840 441186 283892 441192
rect 284024 441186 284076 441192
rect 283562 441144 283618 441153
rect 283852 441114 284064 441130
rect 283562 441079 283618 441088
rect 283840 441108 284076 441114
rect 283576 441046 283604 441079
rect 283892 441102 284024 441108
rect 283840 441050 283892 441056
rect 284024 441050 284076 441056
rect 284588 441046 284616 441322
rect 284852 441312 284904 441318
rect 284852 441254 284904 441260
rect 288900 441312 288952 441318
rect 288900 441254 288952 441260
rect 284864 441046 284892 441254
rect 288912 441182 288940 441254
rect 288900 441176 288952 441182
rect 288900 441118 288952 441124
rect 289280 441046 289308 441390
rect 304920 441386 305302 441402
rect 304908 441380 305302 441386
rect 304960 441374 305302 441380
rect 304908 441322 304960 441328
rect 303068 441312 303120 441318
rect 303120 441260 303370 441266
rect 303068 441254 303370 441260
rect 298652 441244 298704 441250
rect 303080 441238 303370 441254
rect 298652 441186 298704 441192
rect 242348 441040 242400 441046
rect 242716 441040 242768 441046
rect 242348 440982 242400 440988
rect 242466 440988 242716 440994
rect 247868 441040 247920 441046
rect 242466 440982 242768 440988
rect 247710 440988 247868 440994
rect 247710 440982 247920 440988
rect 248052 441040 248104 441046
rect 252008 441040 252060 441046
rect 248052 440982 248104 440988
rect 251666 440988 252008 440994
rect 251666 440982 252060 440988
rect 277400 441040 277452 441046
rect 283104 441040 283156 441046
rect 277400 440982 277452 440988
rect 283102 441008 283104 441017
rect 283564 441040 283616 441046
rect 283156 441008 283158 441017
rect 242466 440966 242756 440982
rect 247710 440966 247908 440982
rect 251666 440966 252048 440982
rect 283564 440982 283616 440988
rect 284576 441040 284628 441046
rect 284576 440982 284628 440988
rect 284852 441040 284904 441046
rect 284852 440982 284904 440988
rect 289268 441040 289320 441046
rect 298664 441017 298692 441186
rect 304998 441144 305054 441153
rect 304998 441079 305054 441088
rect 305012 441046 305040 441079
rect 304356 441040 304408 441046
rect 289268 440982 289320 440988
rect 298650 441008 298706 441017
rect 283102 440943 283158 440952
rect 305000 441040 305052 441046
rect 304408 440988 304658 440994
rect 304356 440982 304658 440988
rect 305000 440982 305052 440988
rect 304368 440966 304658 440982
rect 298650 440943 298706 440952
rect 231216 411256 231268 411262
rect 231216 411198 231268 411204
rect 231124 398812 231176 398818
rect 231124 398754 231176 398760
rect 229744 376032 229796 376038
rect 229744 375974 229796 375980
rect 229836 374740 229888 374746
rect 229836 374682 229888 374688
rect 229744 374400 229796 374406
rect 229744 374342 229796 374348
rect 228456 374264 228508 374270
rect 228456 374206 228508 374212
rect 228468 307358 228496 374206
rect 228548 372836 228600 372842
rect 228548 372778 228600 372784
rect 228560 308310 228588 372778
rect 228640 372700 228692 372706
rect 228640 372642 228692 372648
rect 228652 308825 228680 372642
rect 228732 357468 228784 357474
rect 228732 357410 228784 357416
rect 228744 309534 228772 357410
rect 228824 334008 228876 334014
rect 228824 333950 228876 333956
rect 228836 310690 228864 333950
rect 228824 310684 228876 310690
rect 228824 310626 228876 310632
rect 228732 309528 228784 309534
rect 228732 309470 228784 309476
rect 228638 308816 228694 308825
rect 228638 308751 228694 308760
rect 228548 308304 228600 308310
rect 228548 308246 228600 308252
rect 229756 307426 229784 374342
rect 229848 307630 229876 374682
rect 231124 374196 231176 374202
rect 231124 374138 231176 374144
rect 229928 371680 229980 371686
rect 229928 371622 229980 371628
rect 229940 309126 229968 371622
rect 230020 371408 230072 371414
rect 230020 371350 230072 371356
rect 229928 309120 229980 309126
rect 229928 309062 229980 309068
rect 230032 308922 230060 371350
rect 230112 371340 230164 371346
rect 230112 371282 230164 371288
rect 230020 308916 230072 308922
rect 230020 308858 230072 308864
rect 230124 308242 230152 371282
rect 230204 354748 230256 354754
rect 230204 354690 230256 354696
rect 230216 309874 230244 354690
rect 230296 336796 230348 336802
rect 230296 336738 230348 336744
rect 230308 310214 230336 336738
rect 230388 331288 230440 331294
rect 230388 331230 230440 331236
rect 230296 310208 230348 310214
rect 230296 310150 230348 310156
rect 230204 309868 230256 309874
rect 230204 309810 230256 309816
rect 230400 309670 230428 331230
rect 230940 312996 230992 313002
rect 230940 312938 230992 312944
rect 230388 309664 230440 309670
rect 230388 309606 230440 309612
rect 230952 308650 230980 312938
rect 231032 311364 231084 311370
rect 231032 311306 231084 311312
rect 231044 310078 231072 311306
rect 231032 310072 231084 310078
rect 231032 310014 231084 310020
rect 231136 309913 231164 374138
rect 231216 371612 231268 371618
rect 231216 371554 231268 371560
rect 231122 309904 231178 309913
rect 231122 309839 231178 309848
rect 231228 308990 231256 371554
rect 231400 371544 231452 371550
rect 231400 371486 231452 371492
rect 231308 371476 231360 371482
rect 231308 371418 231360 371424
rect 231320 313002 231348 371418
rect 231308 312996 231360 313002
rect 231308 312938 231360 312944
rect 231412 312882 231440 371486
rect 231492 371272 231544 371278
rect 231492 371214 231544 371220
rect 231320 312854 231440 312882
rect 231320 309097 231348 312854
rect 231400 312724 231452 312730
rect 231400 312666 231452 312672
rect 231412 309262 231440 312666
rect 231400 309256 231452 309262
rect 231400 309198 231452 309204
rect 231306 309088 231362 309097
rect 231504 309058 231532 371214
rect 231584 365764 231636 365770
rect 231584 365706 231636 365712
rect 231596 309466 231624 365706
rect 231676 342304 231728 342310
rect 231676 342246 231728 342252
rect 231688 312730 231716 342246
rect 232228 325712 232280 325718
rect 232280 325666 232360 325694
rect 232228 325654 232280 325660
rect 231768 320204 231820 320210
rect 231768 320146 231820 320152
rect 231676 312724 231728 312730
rect 231676 312666 231728 312672
rect 231780 312610 231808 320146
rect 231860 317484 231912 317490
rect 231860 317426 231912 317432
rect 231688 312582 231808 312610
rect 231584 309460 231636 309466
rect 231584 309402 231636 309408
rect 231688 309330 231716 312582
rect 231872 312066 231900 317426
rect 231952 314696 232004 314702
rect 231952 314638 232004 314644
rect 231780 312038 231900 312066
rect 231780 311846 231808 312038
rect 231860 311908 231912 311914
rect 231860 311850 231912 311856
rect 231768 311840 231820 311846
rect 231768 311782 231820 311788
rect 231768 311228 231820 311234
rect 231768 311170 231820 311176
rect 231780 310162 231808 311170
rect 231872 310282 231900 311850
rect 231964 310350 231992 314638
rect 232044 311840 232096 311846
rect 232044 311782 232096 311788
rect 231952 310344 232004 310350
rect 231952 310286 232004 310292
rect 231860 310276 231912 310282
rect 231860 310218 231912 310224
rect 231780 310134 231900 310162
rect 231676 309324 231728 309330
rect 231676 309266 231728 309272
rect 231306 309023 231362 309032
rect 231492 309052 231544 309058
rect 231492 308994 231544 309000
rect 231216 308984 231268 308990
rect 231216 308926 231268 308932
rect 231872 308854 231900 310134
rect 231952 310072 232004 310078
rect 231952 310014 232004 310020
rect 231860 308848 231912 308854
rect 231860 308790 231912 308796
rect 231964 308786 231992 310014
rect 232056 309398 232084 311782
rect 232136 311296 232188 311302
rect 232136 311238 232188 311244
rect 232148 310554 232176 311238
rect 232228 311160 232280 311166
rect 232228 311102 232280 311108
rect 232136 310548 232188 310554
rect 232136 310490 232188 310496
rect 232240 310332 232268 311102
rect 232332 310729 232360 325666
rect 232318 310720 232374 310729
rect 232318 310655 232374 310664
rect 233148 310616 233200 310622
rect 233148 310558 233200 310564
rect 234434 310584 234490 310593
rect 232780 310548 232832 310554
rect 232780 310490 232832 310496
rect 232516 310332 232544 310420
rect 232596 310412 232648 310418
rect 232596 310354 232648 310360
rect 232240 310304 232544 310332
rect 232608 310298 232636 310354
rect 232700 310298 232728 310420
rect 232608 310270 232728 310298
rect 232792 310298 232820 310490
rect 232962 310448 233018 310457
rect 232884 310298 232912 310420
rect 232962 310383 233018 310392
rect 232792 310270 232912 310298
rect 232976 309942 233004 310383
rect 233160 310298 233188 310558
rect 233700 310548 233752 310554
rect 234434 310519 234490 310528
rect 235814 310584 235870 310593
rect 255608 310554 255806 310570
rect 273732 310554 273930 310570
rect 235814 310519 235870 310528
rect 255412 310548 255464 310554
rect 233700 310490 233752 310496
rect 233252 310298 233280 310420
rect 233160 310270 233280 310298
rect 232964 309936 233016 309942
rect 232964 309878 233016 309884
rect 232044 309392 232096 309398
rect 232044 309334 232096 309340
rect 233620 309126 233648 310420
rect 233712 310298 233740 310490
rect 233804 310298 233832 310420
rect 233712 310270 233832 310298
rect 233608 309120 233660 309126
rect 233608 309062 233660 309068
rect 231952 308780 232004 308786
rect 231952 308722 232004 308728
rect 230940 308644 230992 308650
rect 230940 308586 230992 308592
rect 230112 308236 230164 308242
rect 230112 308178 230164 308184
rect 229836 307624 229888 307630
rect 229836 307566 229888 307572
rect 229744 307420 229796 307426
rect 229744 307362 229796 307368
rect 228456 307352 228508 307358
rect 228456 307294 228508 307300
rect 233988 302234 234016 310420
rect 234172 309194 234200 310420
rect 234160 309188 234212 309194
rect 234160 309130 234212 309136
rect 233344 302206 234016 302234
rect 233344 300082 233372 302206
rect 233332 300076 233384 300082
rect 233332 300018 233384 300024
rect 234356 299305 234384 310420
rect 234448 310298 234476 310519
rect 234540 310298 234568 310420
rect 234448 310270 234568 310298
rect 234342 299296 234398 299305
rect 234342 299231 234398 299240
rect 234724 298586 234752 310420
rect 234922 310406 235028 310434
rect 235000 299266 235028 310406
rect 235184 305454 235212 310420
rect 235368 309058 235396 310420
rect 235552 310350 235580 310420
rect 235540 310344 235592 310350
rect 235540 310286 235592 310292
rect 235356 309052 235408 309058
rect 235356 308994 235408 309000
rect 235736 308990 235764 310420
rect 235828 309126 235856 310519
rect 255412 310490 255464 310496
rect 255596 310548 255806 310554
rect 255648 310542 255806 310548
rect 273536 310548 273588 310554
rect 255596 310490 255648 310496
rect 273536 310490 273588 310496
rect 273720 310548 273930 310554
rect 273772 310542 273930 310548
rect 273720 310490 273772 310496
rect 235920 310146 235948 310420
rect 235908 310140 235960 310146
rect 235908 310082 235960 310088
rect 235816 309120 235868 309126
rect 235816 309062 235868 309068
rect 235724 308984 235776 308990
rect 235724 308926 235776 308932
rect 236104 306218 236132 310420
rect 236288 310282 236316 310420
rect 236276 310276 236328 310282
rect 236276 310218 236328 310224
rect 236104 306190 236316 306218
rect 235172 305448 235224 305454
rect 235172 305390 235224 305396
rect 235908 305448 235960 305454
rect 235908 305390 235960 305396
rect 234988 299260 235040 299266
rect 234988 299202 235040 299208
rect 234712 298580 234764 298586
rect 234712 298522 234764 298528
rect 235920 297090 235948 305390
rect 236184 302252 236236 302258
rect 236184 302194 236236 302200
rect 236196 298722 236224 302194
rect 236184 298716 236236 298722
rect 236184 298658 236236 298664
rect 236288 297770 236316 306190
rect 236472 302326 236500 310420
rect 236552 309324 236604 309330
rect 236552 309266 236604 309272
rect 236564 309194 236592 309266
rect 236552 309188 236604 309194
rect 236552 309130 236604 309136
rect 236656 305454 236684 310420
rect 236644 305448 236696 305454
rect 236644 305390 236696 305396
rect 236460 302320 236512 302326
rect 236460 302262 236512 302268
rect 236840 302234 236868 310420
rect 237024 308446 237052 310420
rect 237012 308440 237064 308446
rect 237012 308382 237064 308388
rect 237208 304638 237236 310420
rect 237392 306406 237420 310420
rect 237380 306400 237432 306406
rect 237380 306342 237432 306348
rect 237196 304632 237248 304638
rect 237196 304574 237248 304580
rect 236380 302206 236868 302234
rect 236276 297764 236328 297770
rect 236276 297706 236328 297712
rect 236380 297158 236408 302206
rect 237576 300150 237604 310420
rect 237668 310406 237866 310434
rect 237564 300144 237616 300150
rect 237564 300086 237616 300092
rect 237668 298081 237696 310406
rect 238036 308553 238064 310420
rect 238220 308922 238248 310420
rect 238208 308916 238260 308922
rect 238208 308858 238260 308864
rect 238022 308544 238078 308553
rect 238022 308479 238078 308488
rect 238404 307154 238432 310420
rect 238588 309126 238616 310420
rect 238772 309874 238800 310420
rect 238956 310214 238984 310420
rect 238944 310208 238996 310214
rect 238944 310150 238996 310156
rect 238760 309868 238812 309874
rect 238760 309810 238812 309816
rect 238576 309120 238628 309126
rect 238576 309062 238628 309068
rect 238392 307148 238444 307154
rect 238392 307090 238444 307096
rect 238944 306536 238996 306542
rect 238944 306478 238996 306484
rect 237932 306400 237984 306406
rect 237932 306342 237984 306348
rect 238852 306400 238904 306406
rect 238852 306342 238904 306348
rect 237654 298072 237710 298081
rect 237654 298007 237710 298016
rect 237944 297906 237972 306342
rect 238864 298926 238892 306342
rect 238956 299334 238984 306478
rect 239036 306468 239088 306474
rect 239036 306410 239088 306416
rect 239048 301617 239076 306410
rect 239034 301608 239090 301617
rect 239034 301543 239090 301552
rect 238944 299328 238996 299334
rect 238944 299270 238996 299276
rect 238852 298920 238904 298926
rect 238852 298862 238904 298868
rect 237932 297900 237984 297906
rect 237932 297842 237984 297848
rect 239140 297838 239168 310420
rect 239324 306406 239352 310420
rect 239508 310010 239536 310420
rect 239496 310004 239548 310010
rect 239496 309946 239548 309952
rect 239692 307018 239720 310420
rect 239680 307012 239732 307018
rect 239680 306954 239732 306960
rect 239876 306542 239904 310420
rect 239864 306536 239916 306542
rect 239864 306478 239916 306484
rect 240060 306474 240088 310420
rect 240336 308650 240364 310420
rect 240324 308644 240376 308650
rect 240324 308586 240376 308592
rect 240520 307000 240548 310420
rect 240152 306972 240548 307000
rect 240048 306468 240100 306474
rect 240048 306410 240100 306416
rect 239312 306400 239364 306406
rect 239312 306342 239364 306348
rect 240152 302190 240180 306972
rect 240232 306400 240284 306406
rect 240232 306342 240284 306348
rect 240140 302184 240192 302190
rect 240140 302126 240192 302132
rect 240244 299402 240272 306342
rect 240704 302308 240732 310420
rect 240428 302280 240732 302308
rect 240428 300286 240456 302280
rect 240888 302234 240916 310420
rect 240520 302206 240916 302234
rect 240416 300280 240468 300286
rect 240416 300222 240468 300228
rect 240520 299470 240548 302206
rect 241072 300218 241100 310420
rect 241256 309505 241284 310420
rect 241242 309496 241298 309505
rect 241242 309431 241298 309440
rect 241440 306406 241468 310420
rect 241624 308922 241652 310420
rect 241808 309670 241836 310420
rect 241796 309664 241848 309670
rect 241796 309606 241848 309612
rect 241612 308916 241664 308922
rect 241612 308858 241664 308864
rect 241992 307698 242020 310420
rect 242176 308242 242204 310420
rect 242360 308582 242388 310420
rect 242348 308576 242400 308582
rect 242348 308518 242400 308524
rect 242164 308236 242216 308242
rect 242164 308178 242216 308184
rect 241980 307692 242032 307698
rect 241980 307634 242032 307640
rect 242544 307494 242572 310420
rect 242532 307488 242584 307494
rect 242532 307430 242584 307436
rect 241428 306400 241480 306406
rect 241428 306342 241480 306348
rect 242728 300354 242756 310420
rect 243004 309534 243032 310420
rect 242992 309528 243044 309534
rect 242992 309470 243044 309476
rect 242808 307828 242860 307834
rect 242808 307770 242860 307776
rect 242820 300490 242848 307770
rect 243084 306400 243136 306406
rect 243084 306342 243136 306348
rect 242808 300484 242860 300490
rect 242808 300426 242860 300432
rect 242716 300348 242768 300354
rect 242716 300290 242768 300296
rect 241060 300212 241112 300218
rect 241060 300154 241112 300160
rect 240508 299464 240560 299470
rect 240508 299406 240560 299412
rect 240232 299396 240284 299402
rect 240232 299338 240284 299344
rect 243096 299062 243124 306342
rect 243188 304570 243216 310420
rect 243372 308689 243400 310420
rect 243358 308680 243414 308689
rect 243358 308615 243414 308624
rect 243556 307834 243584 310420
rect 243544 307828 243596 307834
rect 243544 307770 243596 307776
rect 243740 307766 243768 310420
rect 243728 307760 243780 307766
rect 243728 307702 243780 307708
rect 243924 306354 243952 310420
rect 244004 307896 244056 307902
rect 244004 307838 244056 307844
rect 243372 306326 243952 306354
rect 243176 304564 243228 304570
rect 243176 304506 243228 304512
rect 243372 300422 243400 306326
rect 244016 302234 244044 307838
rect 244108 306406 244136 310420
rect 244292 308961 244320 310420
rect 244476 309942 244504 310420
rect 244464 309936 244516 309942
rect 244660 309913 244688 310420
rect 244464 309878 244516 309884
rect 244646 309904 244702 309913
rect 244646 309839 244702 309848
rect 244278 308952 244334 308961
rect 244278 308887 244334 308896
rect 244844 307562 244872 310420
rect 244832 307556 244884 307562
rect 244832 307498 244884 307504
rect 244096 306400 244148 306406
rect 244096 306342 244148 306348
rect 245028 302234 245056 310420
rect 245212 304978 245240 310420
rect 245488 306202 245516 310420
rect 245672 308122 245700 310420
rect 245856 308854 245884 310420
rect 245844 308848 245896 308854
rect 245844 308790 245896 308796
rect 245672 308094 245884 308122
rect 245752 308032 245804 308038
rect 245752 307974 245804 307980
rect 245476 306196 245528 306202
rect 245476 306138 245528 306144
rect 245200 304972 245252 304978
rect 245200 304914 245252 304920
rect 243556 302206 244044 302234
rect 244476 302206 245056 302234
rect 243360 300416 243412 300422
rect 243360 300358 243412 300364
rect 243084 299056 243136 299062
rect 243084 298998 243136 299004
rect 239128 297832 239180 297838
rect 239128 297774 239180 297780
rect 236368 297152 236420 297158
rect 236368 297094 236420 297100
rect 235908 297084 235960 297090
rect 235908 297026 235960 297032
rect 243556 296682 243584 302206
rect 244476 299198 244504 302206
rect 245764 300694 245792 307974
rect 245856 300801 245884 308094
rect 246040 304502 246068 310420
rect 246028 304496 246080 304502
rect 246028 304438 246080 304444
rect 245842 300792 245898 300801
rect 245842 300727 245898 300736
rect 245752 300688 245804 300694
rect 245752 300630 245804 300636
rect 246224 300626 246252 310420
rect 246408 309369 246436 310420
rect 246394 309360 246450 309369
rect 246394 309295 246450 309304
rect 246592 308825 246620 310420
rect 246578 308816 246634 308825
rect 246578 308751 246634 308760
rect 246776 308242 246804 310420
rect 246764 308236 246816 308242
rect 246764 308178 246816 308184
rect 246304 308168 246356 308174
rect 246304 308110 246356 308116
rect 246212 300620 246264 300626
rect 246212 300562 246264 300568
rect 244464 299192 244516 299198
rect 244464 299134 244516 299140
rect 243544 296676 243596 296682
rect 243544 296618 243596 296624
rect 228364 293956 228416 293962
rect 228364 293898 228416 293904
rect 225604 267708 225656 267714
rect 225604 267650 225656 267656
rect 246316 260166 246344 308110
rect 246960 307290 246988 310420
rect 247144 307358 247172 310420
rect 247328 309777 247356 310420
rect 247314 309768 247370 309777
rect 247314 309703 247370 309712
rect 247512 309466 247540 310420
rect 247500 309460 247552 309466
rect 247500 309402 247552 309408
rect 247132 307352 247184 307358
rect 247132 307294 247184 307300
rect 246948 307284 247000 307290
rect 246948 307226 247000 307232
rect 247696 306354 247724 310420
rect 247776 307828 247828 307834
rect 247776 307770 247828 307776
rect 247144 306326 247724 306354
rect 247144 300558 247172 306326
rect 247224 306196 247276 306202
rect 247224 306138 247276 306144
rect 247132 300552 247184 300558
rect 247132 300494 247184 300500
rect 247236 299130 247264 306138
rect 247684 305448 247736 305454
rect 247684 305390 247736 305396
rect 247224 299124 247276 299130
rect 247224 299066 247276 299072
rect 247696 275330 247724 305390
rect 247788 298654 247816 307770
rect 247880 306202 247908 310420
rect 248156 308786 248184 310420
rect 248340 309097 248368 310420
rect 248326 309088 248382 309097
rect 248326 309023 248382 309032
rect 248144 308780 248196 308786
rect 248144 308722 248196 308728
rect 247960 308712 248012 308718
rect 247960 308654 248012 308660
rect 247868 306196 247920 306202
rect 247868 306138 247920 306144
rect 247972 305454 248000 308654
rect 248524 307834 248552 310420
rect 248512 307828 248564 307834
rect 248512 307770 248564 307776
rect 248512 306400 248564 306406
rect 248512 306342 248564 306348
rect 247960 305448 248012 305454
rect 247960 305390 248012 305396
rect 248524 301209 248552 306342
rect 248708 302234 248736 310420
rect 248892 306406 248920 310420
rect 249076 309641 249104 310420
rect 249062 309632 249118 309641
rect 249062 309567 249118 309576
rect 249260 307902 249288 310420
rect 249248 307896 249300 307902
rect 249248 307838 249300 307844
rect 248880 306400 248932 306406
rect 248880 306342 248932 306348
rect 249444 304434 249472 310420
rect 249628 309398 249656 310420
rect 249616 309392 249668 309398
rect 249616 309334 249668 309340
rect 249812 309194 249840 310420
rect 249800 309188 249852 309194
rect 249800 309130 249852 309136
rect 249996 307222 250024 310420
rect 249984 307216 250036 307222
rect 249984 307158 250036 307164
rect 249892 306400 249944 306406
rect 249892 306342 249944 306348
rect 249432 304428 249484 304434
rect 249432 304370 249484 304376
rect 248616 302206 248736 302234
rect 248510 301200 248566 301209
rect 248510 301135 248566 301144
rect 247776 298648 247828 298654
rect 247776 298590 247828 298596
rect 248616 296614 248644 302206
rect 249904 299441 249932 306342
rect 250180 302234 250208 310420
rect 250364 308378 250392 310420
rect 250640 309233 250668 310420
rect 250626 309224 250682 309233
rect 250626 309159 250682 309168
rect 250444 308576 250496 308582
rect 250444 308518 250496 308524
rect 250352 308372 250404 308378
rect 250352 308314 250404 308320
rect 250352 304428 250404 304434
rect 250352 304370 250404 304376
rect 249996 302206 250208 302234
rect 249996 300830 250024 302206
rect 249984 300824 250036 300830
rect 249984 300766 250036 300772
rect 249890 299432 249946 299441
rect 249890 299367 249946 299376
rect 250364 298994 250392 304370
rect 250352 298988 250404 298994
rect 250352 298930 250404 298936
rect 248604 296608 248656 296614
rect 248604 296550 248656 296556
rect 247684 275324 247736 275330
rect 247684 275266 247736 275272
rect 246304 260160 246356 260166
rect 246304 260102 246356 260108
rect 250456 246430 250484 308518
rect 250536 307896 250588 307902
rect 250536 307838 250588 307844
rect 250548 265674 250576 307838
rect 250824 304434 250852 310420
rect 250904 307828 250956 307834
rect 250904 307770 250956 307776
rect 250812 304428 250864 304434
rect 250812 304370 250864 304376
rect 250916 302234 250944 307770
rect 251008 306406 251036 310420
rect 250996 306400 251048 306406
rect 250996 306342 251048 306348
rect 251192 306354 251220 310420
rect 251376 307834 251404 310420
rect 251364 307828 251416 307834
rect 251364 307770 251416 307776
rect 251192 306326 251496 306354
rect 251364 306196 251416 306202
rect 251364 306138 251416 306144
rect 250640 302206 250944 302234
rect 250640 298858 250668 302206
rect 251376 300762 251404 306138
rect 251364 300756 251416 300762
rect 251364 300698 251416 300704
rect 250628 298852 250680 298858
rect 250628 298794 250680 298800
rect 251468 297974 251496 306326
rect 251560 303074 251588 310420
rect 251744 307426 251772 310420
rect 251928 308038 251956 310420
rect 251916 308032 251968 308038
rect 251916 307974 251968 307980
rect 251824 307964 251876 307970
rect 251824 307906 251876 307912
rect 251732 307420 251784 307426
rect 251732 307362 251784 307368
rect 251732 306400 251784 306406
rect 251732 306342 251784 306348
rect 251548 303068 251600 303074
rect 251548 303010 251600 303016
rect 251744 298790 251772 306342
rect 251732 298784 251784 298790
rect 251732 298726 251784 298732
rect 251456 297968 251508 297974
rect 251456 297910 251508 297916
rect 250536 265668 250588 265674
rect 250536 265610 250588 265616
rect 251836 257446 251864 307906
rect 252112 306406 252140 310420
rect 252192 308100 252244 308106
rect 252192 308042 252244 308048
rect 252100 306400 252152 306406
rect 252100 306342 252152 306348
rect 252204 302234 252232 308042
rect 252296 307630 252324 310420
rect 252284 307624 252336 307630
rect 252284 307566 252336 307572
rect 252480 306202 252508 310420
rect 252664 308281 252692 310420
rect 252848 309262 252876 310420
rect 252836 309256 252888 309262
rect 252836 309198 252888 309204
rect 253032 309134 253060 310420
rect 252940 309106 253060 309134
rect 253124 310406 253322 310434
rect 252650 308272 252706 308281
rect 252650 308207 252706 308216
rect 252652 306400 252704 306406
rect 252652 306342 252704 306348
rect 252468 306196 252520 306202
rect 252468 306138 252520 306144
rect 251928 302206 252232 302234
rect 251928 260370 251956 302206
rect 251916 260364 251968 260370
rect 251916 260306 251968 260312
rect 251824 257440 251876 257446
rect 251824 257382 251876 257388
rect 252664 247722 252692 306342
rect 252940 304314 252968 309106
rect 252848 304286 252968 304314
rect 252744 304224 252796 304230
rect 252744 304166 252796 304172
rect 252756 268394 252784 304166
rect 252848 284986 252876 304286
rect 253124 304230 253152 310406
rect 253204 308644 253256 308650
rect 253204 308586 253256 308592
rect 253112 304224 253164 304230
rect 253112 304166 253164 304172
rect 252928 303884 252980 303890
rect 252928 303826 252980 303832
rect 252836 284980 252888 284986
rect 252836 284922 252888 284928
rect 252744 268388 252796 268394
rect 252744 268330 252796 268336
rect 252652 247716 252704 247722
rect 252652 247658 252704 247664
rect 250444 246424 250496 246430
rect 250444 246366 250496 246372
rect 252940 246362 252968 303826
rect 253216 252006 253244 308586
rect 253296 308508 253348 308514
rect 253296 308450 253348 308456
rect 253308 254726 253336 308450
rect 253492 308174 253520 310420
rect 253480 308168 253532 308174
rect 253480 308110 253532 308116
rect 253388 307896 253440 307902
rect 253388 307838 253440 307844
rect 253400 278050 253428 307838
rect 253676 306406 253704 310420
rect 253664 306400 253716 306406
rect 253664 306342 253716 306348
rect 253860 303890 253888 310420
rect 254044 306354 254072 310420
rect 254044 306326 254164 306354
rect 254032 306196 254084 306202
rect 254032 306138 254084 306144
rect 253848 303884 253900 303890
rect 253848 303826 253900 303832
rect 253388 278044 253440 278050
rect 253388 277986 253440 277992
rect 254044 269822 254072 306138
rect 254136 286346 254164 306326
rect 254228 289134 254256 310420
rect 254412 308718 254440 310420
rect 254400 308712 254452 308718
rect 254400 308654 254452 308660
rect 254596 306354 254624 310420
rect 254320 306326 254624 306354
rect 254320 290494 254348 306326
rect 254780 306202 254808 310420
rect 254768 306196 254820 306202
rect 254768 306138 254820 306144
rect 254964 302234 254992 310420
rect 255148 305794 255176 310420
rect 255332 306542 255360 310420
rect 255320 306536 255372 306542
rect 255320 306478 255372 306484
rect 255136 305788 255188 305794
rect 255136 305730 255188 305736
rect 254412 302206 254992 302234
rect 254308 290488 254360 290494
rect 254308 290430 254360 290436
rect 254216 289128 254268 289134
rect 254216 289070 254268 289076
rect 254124 286340 254176 286346
rect 254124 286282 254176 286288
rect 254032 269816 254084 269822
rect 254032 269758 254084 269764
rect 254412 261526 254440 302206
rect 254400 261520 254452 261526
rect 254400 261462 254452 261468
rect 255424 257378 255452 310490
rect 255530 310406 255728 310434
rect 255504 306468 255556 306474
rect 255504 306410 255556 306416
rect 255516 279478 255544 306410
rect 255596 306400 255648 306406
rect 255596 306342 255648 306348
rect 255700 306354 255728 310406
rect 255872 306536 255924 306542
rect 255872 306478 255924 306484
rect 255608 283626 255636 306342
rect 255700 306326 255820 306354
rect 255688 306196 255740 306202
rect 255688 306138 255740 306144
rect 255700 291854 255728 306138
rect 255688 291848 255740 291854
rect 255688 291790 255740 291796
rect 255596 283620 255648 283626
rect 255596 283562 255648 283568
rect 255504 279472 255556 279478
rect 255504 279414 255556 279420
rect 255412 257372 255464 257378
rect 255412 257314 255464 257320
rect 255792 256018 255820 306326
rect 255884 296002 255912 306478
rect 255976 306474 256004 310420
rect 255964 306468 256016 306474
rect 255964 306410 256016 306416
rect 256160 306406 256188 310420
rect 256148 306400 256200 306406
rect 256148 306342 256200 306348
rect 256344 306202 256372 310420
rect 256528 307970 256556 310420
rect 256516 307964 256568 307970
rect 256516 307906 256568 307912
rect 256332 306196 256384 306202
rect 256332 306138 256384 306144
rect 256712 305386 256740 310420
rect 256792 306400 256844 306406
rect 256792 306342 256844 306348
rect 256700 305380 256752 305386
rect 256700 305322 256752 305328
rect 255872 295996 255924 296002
rect 255872 295938 255924 295944
rect 255780 256012 255832 256018
rect 255780 255954 255832 255960
rect 253296 254720 253348 254726
rect 253296 254662 253348 254668
rect 253204 252000 253256 252006
rect 253204 251942 253256 251948
rect 256804 247790 256832 306342
rect 256896 306218 256924 310420
rect 257080 306354 257108 310420
rect 257080 306326 257200 306354
rect 256896 306190 257108 306218
rect 256976 305788 257028 305794
rect 256976 305730 257028 305736
rect 256884 305448 256936 305454
rect 256884 305390 256936 305396
rect 256896 260302 256924 305390
rect 256884 260296 256936 260302
rect 256884 260238 256936 260244
rect 256988 260234 257016 305730
rect 257080 280838 257108 306190
rect 257172 287706 257200 306326
rect 257160 287700 257212 287706
rect 257160 287642 257212 287648
rect 257068 280832 257120 280838
rect 257068 280774 257120 280780
rect 256976 260228 257028 260234
rect 256976 260170 257028 260176
rect 256792 247784 256844 247790
rect 256792 247726 256844 247732
rect 252928 246356 252980 246362
rect 252928 246298 252980 246304
rect 257264 244934 257292 310420
rect 257448 305454 257476 310420
rect 257632 305794 257660 310420
rect 257816 307834 257844 310420
rect 257804 307828 257856 307834
rect 257804 307770 257856 307776
rect 258000 306406 258028 310420
rect 258184 306490 258212 310420
rect 258092 306462 258212 306490
rect 258276 310406 258474 310434
rect 257988 306400 258040 306406
rect 257988 306342 258040 306348
rect 258092 306202 258120 306462
rect 258276 306354 258304 310406
rect 258644 306354 258672 310420
rect 258184 306326 258304 306354
rect 258460 306326 258672 306354
rect 258080 306196 258132 306202
rect 258080 306138 258132 306144
rect 257620 305788 257672 305794
rect 257620 305730 257672 305736
rect 257436 305448 257488 305454
rect 257436 305390 257488 305396
rect 257344 305380 257396 305386
rect 257344 305322 257396 305328
rect 257356 301578 257384 305322
rect 257344 301572 257396 301578
rect 257344 301514 257396 301520
rect 258184 276690 258212 306326
rect 258264 305788 258316 305794
rect 258264 305730 258316 305736
rect 258276 282198 258304 305730
rect 258356 304700 258408 304706
rect 258356 304642 258408 304648
rect 258368 285054 258396 304642
rect 258460 294642 258488 306326
rect 258540 306196 258592 306202
rect 258540 306138 258592 306144
rect 258552 300121 258580 306138
rect 258828 305794 258856 310420
rect 259012 308582 259040 310420
rect 259000 308576 259052 308582
rect 259000 308518 259052 308524
rect 258816 305788 258868 305794
rect 258816 305730 258868 305736
rect 259196 304706 259224 310420
rect 259184 304700 259236 304706
rect 259184 304642 259236 304648
rect 258538 300112 258594 300121
rect 258538 300047 258594 300056
rect 259380 296714 259408 310420
rect 259564 307902 259592 310420
rect 259748 308106 259776 310420
rect 259932 309134 259960 310420
rect 259840 309106 259960 309134
rect 259736 308100 259788 308106
rect 259736 308042 259788 308048
rect 259552 307896 259604 307902
rect 259552 307838 259604 307844
rect 259552 306468 259604 306474
rect 259552 306410 259604 306416
rect 258644 296686 259408 296714
rect 258448 294636 258500 294642
rect 258448 294578 258500 294584
rect 258356 285048 258408 285054
rect 258356 284990 258408 284996
rect 258264 282192 258316 282198
rect 258264 282134 258316 282140
rect 258172 276684 258224 276690
rect 258172 276626 258224 276632
rect 258644 247858 258672 296686
rect 259564 251938 259592 306410
rect 259644 306400 259696 306406
rect 259644 306342 259696 306348
rect 259656 267034 259684 306342
rect 259736 306196 259788 306202
rect 259736 306138 259788 306144
rect 259748 286414 259776 306138
rect 259840 290562 259868 309106
rect 260116 308802 260144 310420
rect 260116 308774 260236 308802
rect 260104 308644 260156 308650
rect 260104 308586 260156 308592
rect 260012 308100 260064 308106
rect 260012 308042 260064 308048
rect 259828 290556 259880 290562
rect 259828 290498 259880 290504
rect 259736 286408 259788 286414
rect 259736 286350 259788 286356
rect 259644 267028 259696 267034
rect 259644 266970 259696 266976
rect 259552 251932 259604 251938
rect 259552 251874 259604 251880
rect 260024 251870 260052 308042
rect 260116 257582 260144 308586
rect 260208 302977 260236 308774
rect 260300 306202 260328 310420
rect 260380 308848 260432 308854
rect 260380 308790 260432 308796
rect 260288 306196 260340 306202
rect 260288 306138 260340 306144
rect 260194 302968 260250 302977
rect 260194 302903 260250 302912
rect 260392 296714 260420 308790
rect 260484 306406 260512 310420
rect 260668 306474 260696 310420
rect 260840 306604 260892 306610
rect 260840 306546 260892 306552
rect 260656 306468 260708 306474
rect 260656 306410 260708 306416
rect 260472 306400 260524 306406
rect 260472 306342 260524 306348
rect 260208 296686 260420 296714
rect 260208 271318 260236 296686
rect 260852 293282 260880 306546
rect 260944 306474 260972 310420
rect 260932 306468 260984 306474
rect 260932 306410 260984 306416
rect 261128 306218 261156 310420
rect 261312 306610 261340 310420
rect 261300 306604 261352 306610
rect 261300 306546 261352 306552
rect 261208 306468 261260 306474
rect 261208 306410 261260 306416
rect 260944 306190 261156 306218
rect 260840 293276 260892 293282
rect 260840 293218 260892 293224
rect 260196 271312 260248 271318
rect 260196 271254 260248 271260
rect 260104 257576 260156 257582
rect 260104 257518 260156 257524
rect 260012 251864 260064 251870
rect 260012 251806 260064 251812
rect 260944 250510 260972 306190
rect 261024 305788 261076 305794
rect 261024 305730 261076 305736
rect 261036 271182 261064 305730
rect 261116 305448 261168 305454
rect 261116 305390 261168 305396
rect 261128 272542 261156 305390
rect 261220 279546 261248 306410
rect 261300 306400 261352 306406
rect 261300 306342 261352 306348
rect 261312 283694 261340 306342
rect 261496 305794 261524 310420
rect 261484 305788 261536 305794
rect 261484 305730 261536 305736
rect 261680 305674 261708 310420
rect 261760 307896 261812 307902
rect 261760 307838 261812 307844
rect 261404 305646 261708 305674
rect 261300 283688 261352 283694
rect 261300 283630 261352 283636
rect 261208 279540 261260 279546
rect 261208 279482 261260 279488
rect 261116 272536 261168 272542
rect 261116 272478 261168 272484
rect 261024 271176 261076 271182
rect 261024 271118 261076 271124
rect 260932 250504 260984 250510
rect 260932 250446 260984 250452
rect 261404 249082 261432 305646
rect 261772 302234 261800 307838
rect 261864 306406 261892 310420
rect 261852 306400 261904 306406
rect 261852 306342 261904 306348
rect 262048 305454 262076 310420
rect 262232 306354 262260 310420
rect 262416 308990 262444 310420
rect 262404 308984 262456 308990
rect 262404 308926 262456 308932
rect 262600 307018 262628 310420
rect 262588 307012 262640 307018
rect 262588 306954 262640 306960
rect 262680 306808 262732 306814
rect 262680 306750 262732 306756
rect 262232 306326 262444 306354
rect 262312 305788 262364 305794
rect 262312 305730 262364 305736
rect 262036 305448 262088 305454
rect 262036 305390 262088 305396
rect 261496 302206 261800 302234
rect 261496 257514 261524 302206
rect 261484 257508 261536 257514
rect 261484 257450 261536 257456
rect 261392 249076 261444 249082
rect 261392 249018 261444 249024
rect 258632 247852 258684 247858
rect 258632 247794 258684 247800
rect 262324 246498 262352 305730
rect 262416 249150 262444 306326
rect 262588 306196 262640 306202
rect 262588 306138 262640 306144
rect 262496 304224 262548 304230
rect 262496 304166 262548 304172
rect 262508 250578 262536 304166
rect 262600 250646 262628 306138
rect 262588 250640 262640 250646
rect 262588 250582 262640 250588
rect 262496 250572 262548 250578
rect 262496 250514 262548 250520
rect 262404 249144 262456 249150
rect 262404 249086 262456 249092
rect 262312 246492 262364 246498
rect 262312 246434 262364 246440
rect 262692 245002 262720 306750
rect 262784 304230 262812 310420
rect 262772 304224 262824 304230
rect 262772 304166 262824 304172
rect 262968 296714 262996 310420
rect 263152 305794 263180 310420
rect 263336 306202 263364 310420
rect 263612 306474 263640 310420
rect 263600 306468 263652 306474
rect 263600 306410 263652 306416
rect 263796 306354 263824 310420
rect 263980 306513 264008 310420
rect 263966 306504 264022 306513
rect 263876 306468 263928 306474
rect 264164 306474 264192 310420
rect 263966 306439 264022 306448
rect 264152 306468 264204 306474
rect 263876 306410 263928 306416
rect 264152 306410 264204 306416
rect 263612 306326 263824 306354
rect 263324 306196 263376 306202
rect 263324 306138 263376 306144
rect 263140 305788 263192 305794
rect 263140 305730 263192 305736
rect 262784 296686 262996 296714
rect 262784 296070 262812 296686
rect 262772 296064 262824 296070
rect 262772 296006 262824 296012
rect 263612 293350 263640 306326
rect 263782 306232 263838 306241
rect 263692 306196 263744 306202
rect 263782 306167 263838 306176
rect 263692 306138 263744 306144
rect 263600 293344 263652 293350
rect 263600 293286 263652 293292
rect 263704 253230 263732 306138
rect 263796 261594 263824 306167
rect 263888 267102 263916 306410
rect 264060 306400 264112 306406
rect 264060 306342 264112 306348
rect 263968 305788 264020 305794
rect 263968 305730 264020 305736
rect 263980 268462 264008 305730
rect 264072 269890 264100 306342
rect 264348 306184 264376 310420
rect 264428 306468 264480 306474
rect 264428 306410 264480 306416
rect 264164 306156 264376 306184
rect 264164 278118 264192 306156
rect 264440 299474 264468 306410
rect 264532 306202 264560 310420
rect 264520 306196 264572 306202
rect 264520 306138 264572 306144
rect 264716 305794 264744 310420
rect 264900 306406 264928 310420
rect 265084 306406 265112 310420
rect 265268 306490 265296 310420
rect 265176 306462 265296 306490
rect 264888 306400 264940 306406
rect 264888 306342 264940 306348
rect 265072 306400 265124 306406
rect 265072 306342 265124 306348
rect 265176 306218 265204 306462
rect 265256 306400 265308 306406
rect 265256 306342 265308 306348
rect 265348 306400 265400 306406
rect 265348 306342 265400 306348
rect 265084 306190 265204 306218
rect 264704 305788 264756 305794
rect 264704 305730 264756 305736
rect 264980 304700 265032 304706
rect 264980 304642 265032 304648
rect 264256 299446 264468 299474
rect 264152 278112 264204 278118
rect 264152 278054 264204 278060
rect 264060 269884 264112 269890
rect 264060 269826 264112 269832
rect 263968 268456 264020 268462
rect 263968 268398 264020 268404
rect 263876 267096 263928 267102
rect 263876 267038 263928 267044
rect 263784 261588 263836 261594
rect 263784 261530 263836 261536
rect 263692 253224 263744 253230
rect 263692 253166 263744 253172
rect 264256 250714 264284 299446
rect 264244 250708 264296 250714
rect 264244 250650 264296 250656
rect 264992 249218 265020 304642
rect 265084 256086 265112 306190
rect 265164 303680 265216 303686
rect 265164 303622 265216 303628
rect 265176 264246 265204 303622
rect 265268 271250 265296 306342
rect 265360 272610 265388 306342
rect 265452 276758 265480 310420
rect 265636 306406 265664 310420
rect 265624 306400 265676 306406
rect 265624 306342 265676 306348
rect 265820 296714 265848 310420
rect 265912 310406 266110 310434
rect 265912 304706 265940 310406
rect 265900 304700 265952 304706
rect 265900 304642 265952 304648
rect 266280 303686 266308 310420
rect 266464 306354 266492 310420
rect 266648 306474 266676 310420
rect 266636 306468 266688 306474
rect 266636 306410 266688 306416
rect 266832 306354 266860 310420
rect 267016 308922 267044 310420
rect 267004 308916 267056 308922
rect 267004 308858 267056 308864
rect 267004 308508 267056 308514
rect 267004 308450 267056 308456
rect 266912 306468 266964 306474
rect 266912 306410 266964 306416
rect 266464 306326 266584 306354
rect 266452 305448 266504 305454
rect 266452 305390 266504 305396
rect 266268 303680 266320 303686
rect 266268 303622 266320 303628
rect 265544 296686 265848 296714
rect 265544 285122 265572 296686
rect 265532 285116 265584 285122
rect 265532 285058 265584 285064
rect 265440 276752 265492 276758
rect 265440 276694 265492 276700
rect 265348 272604 265400 272610
rect 265348 272546 265400 272552
rect 265256 271244 265308 271250
rect 265256 271186 265308 271192
rect 265164 264240 265216 264246
rect 265164 264182 265216 264188
rect 265072 256080 265124 256086
rect 265072 256022 265124 256028
rect 264980 249212 265032 249218
rect 264980 249154 265032 249160
rect 266464 247926 266492 305390
rect 266556 249286 266584 306326
rect 266648 306326 266860 306354
rect 266648 254590 266676 306326
rect 266728 306196 266780 306202
rect 266728 306138 266780 306144
rect 266740 254658 266768 306138
rect 266820 305788 266872 305794
rect 266820 305730 266872 305736
rect 266832 269958 266860 305730
rect 266820 269952 266872 269958
rect 266820 269894 266872 269900
rect 266728 254652 266780 254658
rect 266728 254594 266780 254600
rect 266636 254584 266688 254590
rect 266636 254526 266688 254532
rect 266544 249280 266596 249286
rect 266544 249222 266596 249228
rect 266452 247920 266504 247926
rect 266452 247862 266504 247868
rect 266924 246566 266952 306410
rect 267016 258874 267044 308450
rect 267200 305454 267228 310420
rect 267384 306202 267412 310420
rect 267372 306196 267424 306202
rect 267372 306138 267424 306144
rect 267568 305794 267596 310420
rect 267752 306406 267780 310420
rect 267936 307018 267964 310420
rect 267924 307012 267976 307018
rect 267924 306954 267976 306960
rect 268016 306808 268068 306814
rect 268016 306750 268068 306756
rect 267832 306536 267884 306542
rect 267832 306478 267884 306484
rect 267740 306400 267792 306406
rect 267740 306342 267792 306348
rect 267556 305788 267608 305794
rect 267556 305730 267608 305736
rect 267188 305448 267240 305454
rect 267188 305390 267240 305396
rect 267004 258868 267056 258874
rect 267004 258810 267056 258816
rect 267844 253298 267872 306478
rect 267924 306196 267976 306202
rect 267924 306138 267976 306144
rect 267936 264314 267964 306138
rect 268028 273970 268056 306750
rect 268120 306542 268148 310420
rect 268108 306536 268160 306542
rect 268108 306478 268160 306484
rect 268108 306400 268160 306406
rect 268108 306342 268160 306348
rect 268120 275398 268148 306342
rect 268304 306202 268332 310420
rect 268292 306196 268344 306202
rect 268292 306138 268344 306144
rect 268488 302234 268516 310420
rect 268764 308854 268792 310420
rect 268752 308848 268804 308854
rect 268752 308790 268804 308796
rect 268212 302206 268516 302234
rect 268212 278186 268240 302206
rect 268948 296714 268976 310420
rect 269132 306202 269160 310420
rect 269212 306400 269264 306406
rect 269212 306342 269264 306348
rect 269316 306354 269344 310420
rect 269500 308038 269528 310420
rect 269684 309134 269712 310420
rect 269592 309106 269712 309134
rect 269488 308032 269540 308038
rect 269488 307974 269540 307980
rect 269120 306196 269172 306202
rect 269120 306138 269172 306144
rect 268304 296686 268976 296714
rect 268200 278180 268252 278186
rect 268200 278122 268252 278128
rect 268108 275392 268160 275398
rect 268108 275334 268160 275340
rect 268016 273964 268068 273970
rect 268016 273906 268068 273912
rect 267924 264308 267976 264314
rect 267924 264250 267976 264256
rect 267832 253292 267884 253298
rect 267832 253234 267884 253240
rect 266912 246560 266964 246566
rect 266912 246502 266964 246508
rect 268304 245070 268332 296686
rect 269224 246634 269252 306342
rect 269316 306326 269436 306354
rect 269304 303748 269356 303754
rect 269304 303690 269356 303696
rect 269316 254794 269344 303690
rect 269408 272678 269436 306326
rect 269488 306196 269540 306202
rect 269488 306138 269540 306144
rect 269500 276826 269528 306138
rect 269592 304314 269620 309106
rect 269764 308032 269816 308038
rect 269764 307974 269816 307980
rect 269592 304286 269712 304314
rect 269580 302524 269632 302530
rect 269580 302466 269632 302472
rect 269592 282266 269620 302466
rect 269580 282260 269632 282266
rect 269580 282202 269632 282208
rect 269488 276820 269540 276826
rect 269488 276762 269540 276768
rect 269396 272672 269448 272678
rect 269396 272614 269448 272620
rect 269304 254788 269356 254794
rect 269304 254730 269356 254736
rect 269212 246628 269264 246634
rect 269212 246570 269264 246576
rect 269684 245138 269712 304286
rect 269776 289202 269804 307974
rect 269868 307902 269896 310420
rect 269856 307896 269908 307902
rect 269856 307838 269908 307844
rect 270052 302530 270080 310420
rect 270236 306406 270264 310420
rect 270224 306400 270276 306406
rect 270224 306342 270276 306348
rect 270420 303754 270448 310420
rect 270408 303748 270460 303754
rect 270408 303690 270460 303696
rect 270040 302524 270092 302530
rect 270040 302466 270092 302472
rect 269764 289196 269816 289202
rect 269764 289138 269816 289144
rect 270604 253366 270632 310420
rect 270684 306468 270736 306474
rect 270684 306410 270736 306416
rect 270696 264382 270724 306410
rect 270788 306354 270816 310420
rect 270972 306474 271000 310420
rect 271064 310406 271262 310434
rect 270960 306468 271012 306474
rect 270960 306410 271012 306416
rect 270788 306326 271000 306354
rect 270868 306196 270920 306202
rect 270868 306138 270920 306144
rect 270776 305788 270828 305794
rect 270776 305730 270828 305736
rect 270788 265810 270816 305730
rect 270776 265804 270828 265810
rect 270776 265746 270828 265752
rect 270880 265742 270908 306138
rect 270972 275466 271000 306326
rect 271064 306202 271092 310406
rect 271236 308576 271288 308582
rect 271236 308518 271288 308524
rect 271052 306196 271104 306202
rect 271052 306138 271104 306144
rect 271052 305448 271104 305454
rect 271052 305390 271104 305396
rect 270960 275460 271012 275466
rect 270960 275402 271012 275408
rect 270868 265736 270920 265742
rect 270868 265678 270920 265684
rect 270684 264376 270736 264382
rect 270684 264318 270736 264324
rect 271064 253434 271092 305390
rect 271248 302234 271276 308518
rect 271432 305794 271460 310420
rect 271616 308650 271644 310420
rect 271604 308644 271656 308650
rect 271604 308586 271656 308592
rect 271420 305788 271472 305794
rect 271420 305730 271472 305736
rect 271800 305454 271828 310420
rect 271984 306354 272012 310420
rect 271984 306326 272104 306354
rect 271972 306196 272024 306202
rect 271972 306138 272024 306144
rect 271788 305448 271840 305454
rect 271788 305390 271840 305396
rect 271156 302206 271276 302234
rect 271156 291922 271184 302206
rect 271144 291916 271196 291922
rect 271144 291858 271196 291864
rect 271984 256222 272012 306138
rect 271972 256216 272024 256222
rect 271972 256158 272024 256164
rect 272076 256154 272104 306326
rect 272168 274038 272196 310420
rect 272248 306400 272300 306406
rect 272248 306342 272300 306348
rect 272260 280906 272288 306342
rect 272248 280900 272300 280906
rect 272248 280842 272300 280848
rect 272156 274032 272208 274038
rect 272156 273974 272208 273980
rect 272064 256148 272116 256154
rect 272064 256090 272116 256096
rect 271052 253428 271104 253434
rect 271052 253370 271104 253376
rect 270592 253360 270644 253366
rect 270592 253302 270644 253308
rect 272352 246702 272380 310420
rect 272536 306202 272564 310420
rect 272720 308446 272748 310420
rect 272708 308440 272760 308446
rect 272708 308382 272760 308388
rect 272524 306196 272576 306202
rect 272524 306138 272576 306144
rect 272904 296714 272932 310420
rect 273088 306406 273116 310420
rect 273076 306400 273128 306406
rect 273076 306342 273128 306348
rect 273272 306354 273300 310420
rect 273456 308582 273484 310420
rect 273444 308576 273496 308582
rect 273444 308518 273496 308524
rect 273272 306326 273484 306354
rect 273352 306196 273404 306202
rect 273352 306138 273404 306144
rect 272444 296686 272932 296714
rect 272444 296138 272472 296686
rect 272432 296132 272484 296138
rect 272432 296074 272484 296080
rect 273364 265878 273392 306138
rect 273456 275534 273484 306326
rect 273548 282334 273576 310490
rect 273654 310406 273852 310434
rect 273720 306468 273772 306474
rect 273720 306410 273772 306416
rect 273628 306400 273680 306406
rect 273628 306342 273680 306348
rect 273640 289270 273668 306342
rect 273628 289264 273680 289270
rect 273628 289206 273680 289212
rect 273536 282328 273588 282334
rect 273536 282270 273588 282276
rect 273444 275528 273496 275534
rect 273444 275470 273496 275476
rect 273352 265872 273404 265878
rect 273352 265814 273404 265820
rect 273732 250782 273760 306410
rect 273824 296206 273852 310406
rect 274100 306406 274128 310420
rect 274088 306400 274140 306406
rect 274088 306342 274140 306348
rect 274284 306202 274312 310420
rect 274468 306474 274496 310420
rect 274456 306468 274508 306474
rect 274456 306410 274508 306416
rect 274652 306354 274680 310420
rect 274652 306326 274772 306354
rect 274272 306196 274324 306202
rect 274272 306138 274324 306144
rect 274640 304632 274692 304638
rect 274640 304574 274692 304580
rect 273812 296200 273864 296206
rect 273812 296142 273864 296148
rect 274652 290630 274680 304574
rect 274744 294710 274772 306326
rect 274732 294704 274784 294710
rect 274732 294646 274784 294652
rect 274640 290624 274692 290630
rect 274640 290566 274692 290572
rect 274836 276894 274864 310420
rect 274916 306400 274968 306406
rect 274916 306342 274968 306348
rect 274928 280974 274956 306342
rect 275020 283762 275048 310420
rect 275204 306354 275232 310420
rect 275112 306326 275232 306354
rect 275112 287774 275140 306326
rect 275388 302234 275416 310420
rect 275572 306406 275600 310420
rect 275560 306400 275612 306406
rect 275560 306342 275612 306348
rect 275756 304638 275784 310420
rect 275744 304632 275796 304638
rect 275744 304574 275796 304580
rect 275204 302206 275416 302234
rect 275100 287768 275152 287774
rect 275100 287710 275152 287716
rect 275008 283756 275060 283762
rect 275008 283698 275060 283704
rect 274916 280968 274968 280974
rect 274916 280910 274968 280916
rect 274824 276888 274876 276894
rect 274824 276830 274876 276836
rect 273720 250776 273772 250782
rect 273720 250718 273772 250724
rect 275204 247994 275232 302206
rect 275940 296714 275968 310420
rect 276138 310406 276244 310434
rect 276112 306400 276164 306406
rect 276112 306342 276164 306348
rect 276020 305108 276072 305114
rect 276020 305050 276072 305056
rect 275296 296686 275968 296714
rect 275296 264450 275324 296686
rect 276032 290766 276060 305050
rect 276020 290760 276072 290766
rect 276020 290702 276072 290708
rect 275284 264444 275336 264450
rect 275284 264386 275336 264392
rect 276124 262886 276152 306342
rect 276216 268530 276244 310406
rect 276400 307018 276428 310420
rect 276388 307012 276440 307018
rect 276388 306954 276440 306960
rect 276480 306808 276532 306814
rect 276480 306750 276532 306756
rect 276388 305448 276440 305454
rect 276388 305390 276440 305396
rect 276296 300892 276348 300898
rect 276296 300834 276348 300840
rect 276308 278254 276336 300834
rect 276400 285190 276428 305390
rect 276492 286482 276520 306750
rect 276584 300898 276612 310420
rect 276572 300892 276624 300898
rect 276572 300834 276624 300840
rect 276768 296714 276796 310420
rect 276952 305454 276980 310420
rect 276940 305448 276992 305454
rect 276940 305390 276992 305396
rect 277136 305114 277164 310420
rect 277320 306406 277348 310420
rect 277308 306400 277360 306406
rect 277308 306342 277360 306348
rect 277400 306400 277452 306406
rect 277400 306342 277452 306348
rect 277124 305108 277176 305114
rect 277124 305050 277176 305056
rect 276584 296686 276796 296714
rect 276480 286476 276532 286482
rect 276480 286418 276532 286424
rect 276388 285184 276440 285190
rect 276388 285126 276440 285132
rect 276296 278248 276348 278254
rect 276296 278190 276348 278196
rect 276204 268524 276256 268530
rect 276204 268466 276256 268472
rect 276112 262880 276164 262886
rect 276112 262822 276164 262828
rect 276584 261730 276612 296686
rect 276572 261724 276624 261730
rect 276572 261666 276624 261672
rect 277412 252210 277440 306342
rect 277504 306202 277532 310420
rect 277688 306746 277716 310420
rect 277676 306740 277728 306746
rect 277676 306682 277728 306688
rect 277872 306626 277900 310420
rect 277596 306598 277900 306626
rect 277492 306196 277544 306202
rect 277492 306138 277544 306144
rect 277596 306082 277624 306598
rect 277676 306468 277728 306474
rect 277676 306410 277728 306416
rect 277504 306054 277624 306082
rect 277400 252204 277452 252210
rect 277400 252146 277452 252152
rect 277504 252142 277532 306054
rect 277584 305856 277636 305862
rect 277584 305798 277636 305804
rect 277596 261798 277624 305798
rect 277688 262954 277716 306410
rect 278056 306354 278084 310420
rect 277780 306326 278084 306354
rect 277780 282402 277808 306326
rect 277860 306196 277912 306202
rect 277860 306138 277912 306144
rect 277872 283898 277900 306138
rect 278240 305862 278268 310420
rect 278424 306406 278452 310420
rect 278412 306400 278464 306406
rect 278412 306342 278464 306348
rect 278228 305856 278280 305862
rect 278228 305798 278280 305804
rect 278608 300257 278636 310420
rect 278806 310406 278912 310434
rect 278780 306536 278832 306542
rect 278780 306478 278832 306484
rect 278594 300248 278650 300257
rect 278594 300183 278650 300192
rect 278792 294778 278820 306478
rect 278884 306406 278912 310406
rect 278976 310406 279082 310434
rect 278872 306400 278924 306406
rect 278872 306342 278924 306348
rect 278872 305856 278924 305862
rect 278872 305798 278924 305804
rect 278780 294772 278832 294778
rect 278780 294714 278832 294720
rect 277860 283892 277912 283898
rect 277860 283834 277912 283840
rect 277768 282396 277820 282402
rect 277768 282338 277820 282344
rect 278884 270026 278912 305798
rect 278976 274106 279004 310406
rect 279056 306468 279108 306474
rect 279056 306410 279108 306416
rect 279068 279614 279096 306410
rect 279148 306400 279200 306406
rect 279148 306342 279200 306348
rect 279252 306354 279280 310420
rect 279436 306474 279464 310420
rect 279424 306468 279476 306474
rect 279424 306410 279476 306416
rect 279160 291990 279188 306342
rect 279252 306326 279372 306354
rect 279240 306196 279292 306202
rect 279240 306138 279292 306144
rect 279148 291984 279200 291990
rect 279148 291926 279200 291932
rect 279056 279608 279108 279614
rect 279056 279550 279108 279556
rect 278964 274100 279016 274106
rect 278964 274042 279016 274048
rect 278872 270020 278924 270026
rect 278872 269962 278924 269968
rect 277676 262948 277728 262954
rect 277676 262890 277728 262896
rect 277584 261792 277636 261798
rect 277584 261734 277636 261740
rect 277492 252136 277544 252142
rect 277492 252078 277544 252084
rect 275192 247988 275244 247994
rect 275192 247930 275244 247936
rect 272340 246696 272392 246702
rect 272340 246638 272392 246644
rect 279252 245206 279280 306138
rect 279344 300393 279372 306326
rect 279620 305862 279648 310420
rect 279804 306542 279832 310420
rect 279792 306536 279844 306542
rect 279792 306478 279844 306484
rect 279988 306202 280016 310420
rect 279976 306196 280028 306202
rect 279976 306138 280028 306144
rect 280068 306196 280120 306202
rect 280068 306138 280120 306144
rect 279608 305856 279660 305862
rect 279608 305798 279660 305804
rect 280080 305658 280108 306138
rect 280068 305652 280120 305658
rect 280068 305594 280120 305600
rect 280172 305454 280200 310420
rect 280356 306474 280384 310420
rect 280344 306468 280396 306474
rect 280344 306410 280396 306416
rect 280540 306218 280568 310420
rect 280448 306190 280568 306218
rect 280448 305946 280476 306190
rect 280356 305918 280476 305946
rect 280252 305652 280304 305658
rect 280252 305594 280304 305600
rect 280160 305448 280212 305454
rect 280160 305390 280212 305396
rect 279330 300384 279386 300393
rect 279330 300319 279386 300328
rect 280264 248062 280292 305594
rect 280356 252278 280384 305918
rect 280436 305856 280488 305862
rect 280436 305798 280488 305804
rect 280448 253570 280476 305798
rect 280528 305448 280580 305454
rect 280528 305390 280580 305396
rect 280540 254862 280568 305390
rect 280724 302234 280752 310420
rect 280804 306468 280856 306474
rect 280804 306410 280856 306416
rect 280632 302206 280752 302234
rect 280632 258806 280660 302206
rect 280816 296714 280844 306410
rect 280908 305658 280936 310420
rect 281092 305862 281120 310420
rect 281276 308514 281304 310420
rect 281264 308508 281316 308514
rect 281264 308450 281316 308456
rect 281552 306202 281580 310420
rect 281736 306218 281764 310420
rect 281920 306354 281948 310420
rect 282104 306490 282132 310420
rect 282104 306462 282224 306490
rect 281920 306326 282132 306354
rect 281540 306196 281592 306202
rect 281736 306190 281948 306218
rect 281540 306138 281592 306144
rect 281080 305856 281132 305862
rect 281080 305798 281132 305804
rect 281816 305856 281868 305862
rect 281816 305798 281868 305804
rect 280896 305652 280948 305658
rect 280896 305594 280948 305600
rect 281724 305652 281776 305658
rect 281724 305594 281776 305600
rect 280724 296686 280844 296714
rect 280620 258800 280672 258806
rect 280620 258742 280672 258748
rect 280528 254856 280580 254862
rect 280528 254798 280580 254804
rect 280436 253564 280488 253570
rect 280436 253506 280488 253512
rect 280344 252272 280396 252278
rect 280344 252214 280396 252220
rect 280252 248056 280304 248062
rect 280252 247998 280304 248004
rect 280724 245274 280752 296686
rect 281736 276962 281764 305594
rect 281828 278322 281856 305798
rect 281920 287842 281948 306190
rect 281908 287836 281960 287842
rect 281908 287778 281960 287784
rect 281816 278316 281868 278322
rect 281816 278258 281868 278264
rect 281724 276956 281776 276962
rect 281724 276898 281776 276904
rect 282104 271386 282132 306326
rect 282196 302841 282224 306462
rect 282288 305862 282316 310420
rect 282368 305992 282420 305998
rect 282368 305934 282420 305940
rect 282276 305856 282328 305862
rect 282276 305798 282328 305804
rect 282380 305386 282408 305934
rect 282368 305380 282420 305386
rect 282368 305322 282420 305328
rect 282182 302832 282238 302841
rect 282182 302767 282238 302776
rect 282472 296714 282500 310420
rect 282550 306232 282606 306241
rect 282550 306167 282606 306176
rect 282564 306066 282592 306167
rect 282552 306060 282604 306066
rect 282552 306002 282604 306008
rect 282656 302938 282684 310420
rect 282736 306536 282788 306542
rect 282736 306478 282788 306484
rect 282748 306134 282776 306478
rect 282736 306128 282788 306134
rect 282736 306070 282788 306076
rect 282736 305924 282788 305930
rect 282736 305866 282788 305872
rect 282748 305454 282776 305866
rect 282840 305658 282868 310420
rect 282920 306400 282972 306406
rect 282920 306342 282972 306348
rect 282828 305652 282880 305658
rect 282828 305594 282880 305600
rect 282736 305448 282788 305454
rect 282736 305390 282788 305396
rect 282644 302932 282696 302938
rect 282644 302874 282696 302880
rect 282932 301510 282960 306342
rect 283024 302234 283052 310420
rect 283208 306490 283236 310420
rect 283116 306462 283236 306490
rect 283116 304298 283144 306462
rect 283392 306354 283420 310420
rect 283300 306326 283420 306354
rect 283196 305652 283248 305658
rect 283196 305594 283248 305600
rect 283104 304292 283156 304298
rect 283104 304234 283156 304240
rect 283024 302206 283144 302234
rect 282920 301504 282972 301510
rect 282920 301446 282972 301452
rect 282196 296686 282500 296714
rect 282092 271380 282144 271386
rect 282092 271322 282144 271328
rect 282196 249354 282224 296686
rect 283116 272746 283144 302206
rect 283208 275602 283236 305594
rect 283300 286550 283328 306326
rect 283380 306264 283432 306270
rect 283380 306206 283432 306212
rect 283288 286544 283340 286550
rect 283288 286486 283340 286492
rect 283196 275596 283248 275602
rect 283196 275538 283248 275544
rect 283104 272740 283156 272746
rect 283104 272682 283156 272688
rect 282184 249348 282236 249354
rect 282184 249290 282236 249296
rect 283392 245342 283420 306206
rect 283576 296714 283604 310420
rect 283760 306406 283788 310420
rect 283748 306400 283800 306406
rect 283748 306342 283800 306348
rect 283654 306232 283710 306241
rect 283654 306167 283710 306176
rect 283668 306066 283696 306167
rect 283656 306060 283708 306066
rect 283656 306002 283708 306008
rect 283944 305658 283972 310420
rect 284036 310406 284234 310434
rect 284036 306270 284064 310406
rect 284404 306490 284432 310420
rect 284312 306462 284432 306490
rect 284208 306332 284260 306338
rect 284208 306274 284260 306280
rect 284024 306264 284076 306270
rect 284024 306206 284076 306212
rect 284220 305998 284248 306274
rect 284208 305992 284260 305998
rect 284208 305934 284260 305940
rect 284312 305726 284340 306462
rect 284392 306400 284444 306406
rect 284588 306354 284616 310420
rect 284392 306342 284444 306348
rect 284300 305720 284352 305726
rect 284300 305662 284352 305668
rect 283932 305652 283984 305658
rect 283932 305594 283984 305600
rect 283484 296686 283604 296714
rect 283484 265946 283512 296686
rect 284404 272814 284432 306342
rect 284496 306326 284616 306354
rect 284668 306332 284720 306338
rect 284496 274174 284524 306326
rect 284668 306274 284720 306280
rect 284576 306264 284628 306270
rect 284576 306206 284628 306212
rect 284588 289338 284616 306206
rect 284680 293418 284708 306274
rect 284668 293412 284720 293418
rect 284668 293354 284720 293360
rect 284576 289332 284628 289338
rect 284576 289274 284628 289280
rect 284484 274168 284536 274174
rect 284484 274110 284536 274116
rect 284392 272808 284444 272814
rect 284392 272750 284444 272756
rect 283472 265940 283524 265946
rect 283472 265882 283524 265888
rect 284772 248130 284800 310420
rect 284956 307086 284984 310420
rect 284944 307080 284996 307086
rect 284944 307022 284996 307028
rect 285140 306406 285168 310420
rect 285128 306400 285180 306406
rect 285128 306342 285180 306348
rect 285324 306270 285352 310420
rect 285508 306338 285536 310420
rect 285692 308038 285720 310420
rect 285876 309134 285904 310420
rect 285784 309106 285904 309134
rect 285680 308032 285732 308038
rect 285680 307974 285732 307980
rect 285680 306400 285732 306406
rect 285680 306342 285732 306348
rect 285496 306332 285548 306338
rect 285496 306274 285548 306280
rect 285312 306264 285364 306270
rect 285312 306206 285364 306212
rect 284944 305924 284996 305930
rect 284944 305866 284996 305872
rect 284852 305788 284904 305794
rect 284852 305730 284904 305736
rect 284864 305386 284892 305730
rect 284956 305454 284984 305866
rect 284944 305448 284996 305454
rect 284944 305390 284996 305396
rect 284852 305380 284904 305386
rect 284852 305322 284904 305328
rect 285692 304366 285720 306342
rect 285680 304360 285732 304366
rect 285680 304302 285732 304308
rect 285784 300014 285812 309106
rect 285956 308032 286008 308038
rect 285956 307974 286008 307980
rect 285864 306264 285916 306270
rect 285864 306206 285916 306212
rect 285772 300008 285824 300014
rect 285772 299950 285824 299956
rect 285876 271454 285904 306206
rect 285968 284889 285996 307974
rect 286060 306474 286088 310420
rect 286244 306474 286272 310420
rect 286048 306468 286100 306474
rect 286048 306410 286100 306416
rect 286232 306468 286284 306474
rect 286232 306410 286284 306416
rect 286428 306354 286456 310420
rect 286060 306326 286456 306354
rect 286520 310406 286718 310434
rect 285954 284880 286010 284889
rect 285954 284815 286010 284824
rect 285864 271448 285916 271454
rect 285864 271390 285916 271396
rect 286060 250850 286088 306326
rect 286140 306264 286192 306270
rect 286140 306206 286192 306212
rect 286152 269793 286180 306206
rect 286520 296714 286548 310406
rect 286888 306270 286916 310420
rect 287072 306882 287100 310420
rect 287060 306876 287112 306882
rect 287060 306818 287112 306824
rect 287256 306490 287284 310420
rect 287336 306876 287388 306882
rect 287336 306818 287388 306824
rect 287072 306462 287284 306490
rect 286876 306264 286928 306270
rect 286876 306206 286928 306212
rect 287072 303249 287100 306462
rect 287152 306264 287204 306270
rect 287152 306206 287204 306212
rect 287244 306264 287296 306270
rect 287244 306206 287296 306212
rect 287058 303240 287114 303249
rect 287058 303175 287114 303184
rect 286244 296686 286548 296714
rect 286244 296274 286272 296686
rect 286232 296268 286284 296274
rect 286232 296210 286284 296216
rect 286138 269784 286194 269793
rect 286138 269719 286194 269728
rect 287164 254561 287192 306206
rect 287256 256358 287284 306206
rect 287348 261866 287376 306818
rect 287440 306338 287468 310420
rect 287624 306490 287652 310420
rect 287532 306462 287652 306490
rect 287428 306332 287480 306338
rect 287428 306274 287480 306280
rect 287428 305720 287480 305726
rect 287428 305662 287480 305668
rect 287440 301753 287468 305662
rect 287426 301744 287482 301753
rect 287426 301679 287482 301688
rect 287336 261860 287388 261866
rect 287336 261802 287388 261808
rect 287244 256352 287296 256358
rect 287244 256294 287296 256300
rect 287150 254552 287206 254561
rect 287150 254487 287206 254496
rect 286048 250844 286100 250850
rect 286048 250786 286100 250792
rect 287532 250481 287560 306462
rect 287808 305726 287836 310420
rect 287992 306270 288020 310420
rect 287980 306264 288032 306270
rect 287980 306206 288032 306212
rect 287796 305720 287848 305726
rect 287796 305662 287848 305668
rect 288176 302734 288204 310420
rect 288360 306105 288388 310420
rect 288544 306542 288572 310420
rect 288532 306536 288584 306542
rect 288532 306478 288584 306484
rect 288346 306096 288402 306105
rect 288346 306031 288402 306040
rect 288728 303113 288756 310420
rect 288912 305969 288940 310420
rect 289096 306202 289124 310420
rect 289084 306196 289136 306202
rect 289084 306138 289136 306144
rect 288898 305960 288954 305969
rect 288898 305895 288954 305904
rect 289372 303414 289400 310420
rect 289556 305522 289584 310420
rect 289544 305516 289596 305522
rect 289544 305458 289596 305464
rect 289360 303408 289412 303414
rect 289360 303350 289412 303356
rect 288714 303104 288770 303113
rect 288714 303039 288770 303048
rect 289740 302870 289768 310420
rect 289924 303142 289952 310420
rect 290108 305833 290136 310420
rect 290094 305824 290150 305833
rect 290094 305759 290150 305768
rect 290188 304564 290240 304570
rect 290188 304506 290240 304512
rect 289912 303136 289964 303142
rect 289912 303078 289964 303084
rect 289728 302864 289780 302870
rect 289728 302806 289780 302812
rect 288164 302728 288216 302734
rect 288164 302670 288216 302676
rect 290200 297537 290228 304506
rect 290292 302802 290320 310420
rect 290280 302796 290332 302802
rect 290280 302738 290332 302744
rect 290476 302234 290504 310420
rect 290660 305590 290688 310420
rect 290648 305584 290700 305590
rect 290648 305526 290700 305532
rect 290844 303482 290872 310420
rect 291028 304570 291056 310420
rect 291212 305697 291240 310420
rect 291198 305688 291254 305697
rect 291198 305623 291254 305632
rect 291016 304564 291068 304570
rect 291016 304506 291068 304512
rect 291396 303550 291424 310420
rect 291594 310406 291700 310434
rect 291568 306332 291620 306338
rect 291568 306274 291620 306280
rect 291384 303544 291436 303550
rect 291384 303486 291436 303492
rect 290832 303476 290884 303482
rect 290832 303418 290884 303424
rect 290292 302206 290504 302234
rect 290292 299946 290320 302206
rect 290280 299940 290332 299946
rect 290280 299882 290332 299888
rect 290186 297528 290242 297537
rect 290186 297463 290242 297472
rect 291580 297401 291608 306274
rect 291672 297673 291700 310406
rect 291856 305998 291884 310420
rect 291844 305992 291896 305998
rect 291844 305934 291896 305940
rect 292040 303210 292068 310420
rect 292224 306338 292252 310420
rect 292212 306332 292264 306338
rect 292212 306274 292264 306280
rect 292408 305794 292436 310420
rect 292396 305788 292448 305794
rect 292396 305730 292448 305736
rect 292592 303278 292620 310420
rect 292776 307018 292804 310420
rect 292764 307012 292816 307018
rect 292764 306954 292816 306960
rect 292960 306898 292988 310420
rect 292684 306870 292988 306898
rect 292684 305930 292712 306870
rect 293144 306626 293172 310420
rect 292868 306598 293172 306626
rect 292672 305924 292724 305930
rect 292672 305866 292724 305872
rect 292868 303618 292896 306598
rect 293328 306490 293356 310420
rect 293408 307012 293460 307018
rect 293408 306954 293460 306960
rect 293052 306462 293356 306490
rect 293052 305810 293080 306462
rect 293132 306332 293184 306338
rect 293132 306274 293184 306280
rect 292960 305782 293080 305810
rect 292856 303612 292908 303618
rect 292856 303554 292908 303560
rect 292580 303272 292632 303278
rect 292580 303214 292632 303220
rect 292028 303204 292080 303210
rect 292028 303146 292080 303152
rect 292960 301481 292988 305782
rect 293040 305720 293092 305726
rect 293040 305662 293092 305668
rect 292946 301472 293002 301481
rect 292946 301407 293002 301416
rect 291658 297664 291714 297673
rect 291658 297599 291714 297608
rect 293052 297498 293080 305662
rect 293040 297492 293092 297498
rect 293040 297434 293092 297440
rect 291566 297392 291622 297401
rect 293144 297362 293172 306274
rect 293420 302234 293448 306954
rect 293512 306066 293540 310420
rect 293696 306338 293724 310420
rect 293684 306332 293736 306338
rect 293684 306274 293736 306280
rect 293500 306060 293552 306066
rect 293500 306002 293552 306008
rect 293880 305726 293908 310420
rect 293868 305720 293920 305726
rect 293868 305662 293920 305668
rect 294064 303006 294092 310420
rect 294248 306542 294276 310420
rect 294340 310406 294538 310434
rect 294236 306536 294288 306542
rect 294236 306478 294288 306484
rect 294236 306264 294288 306270
rect 294236 306206 294288 306212
rect 294144 304904 294196 304910
rect 294144 304846 294196 304852
rect 294052 303000 294104 303006
rect 294052 302942 294104 302948
rect 293236 302206 293448 302234
rect 291566 297327 291622 297336
rect 293132 297356 293184 297362
rect 293132 297298 293184 297304
rect 293236 297226 293264 302206
rect 294156 297430 294184 304846
rect 294248 297634 294276 306206
rect 294340 304910 294368 310406
rect 294708 305862 294736 310420
rect 294696 305856 294748 305862
rect 294696 305798 294748 305804
rect 294328 304904 294380 304910
rect 294328 304846 294380 304852
rect 294328 304768 294380 304774
rect 294328 304710 294380 304716
rect 294236 297628 294288 297634
rect 294236 297570 294288 297576
rect 294144 297424 294196 297430
rect 294144 297366 294196 297372
rect 293224 297220 293276 297226
rect 293224 297162 293276 297168
rect 294340 294574 294368 304710
rect 294892 302234 294920 310420
rect 295076 304774 295104 310420
rect 295064 304768 295116 304774
rect 295064 304710 295116 304716
rect 294432 302206 294920 302234
rect 294432 297702 294460 302206
rect 294420 297696 294472 297702
rect 294420 297638 294472 297644
rect 295260 297294 295288 310420
rect 295340 304224 295392 304230
rect 295340 304166 295392 304172
rect 295352 301782 295380 304166
rect 295444 303346 295472 310420
rect 295628 307222 295656 310420
rect 295616 307216 295668 307222
rect 295616 307158 295668 307164
rect 295812 306610 295840 310420
rect 295892 307216 295944 307222
rect 295892 307158 295944 307164
rect 295800 306604 295852 306610
rect 295800 306546 295852 306552
rect 295800 306400 295852 306406
rect 295800 306342 295852 306348
rect 295524 306332 295576 306338
rect 295524 306274 295576 306280
rect 295432 303340 295484 303346
rect 295432 303282 295484 303288
rect 295340 301776 295392 301782
rect 295340 301718 295392 301724
rect 295248 297288 295300 297294
rect 295248 297230 295300 297236
rect 295536 294982 295564 306274
rect 295708 306196 295760 306202
rect 295708 306138 295760 306144
rect 295616 306128 295668 306134
rect 295616 306070 295668 306076
rect 295524 294976 295576 294982
rect 295524 294918 295576 294924
rect 295628 294846 295656 306070
rect 295720 295050 295748 306138
rect 295708 295044 295760 295050
rect 295708 294986 295760 294992
rect 295812 294914 295840 306342
rect 295800 294908 295852 294914
rect 295800 294850 295852 294856
rect 295616 294840 295668 294846
rect 295616 294782 295668 294788
rect 294328 294568 294380 294574
rect 294328 294510 294380 294516
rect 295904 294506 295932 307158
rect 295996 306338 296024 310420
rect 295984 306332 296036 306338
rect 295984 306274 296036 306280
rect 296180 304230 296208 310420
rect 296364 306134 296392 310420
rect 296548 306202 296576 310420
rect 296746 310406 296852 310434
rect 296720 306536 296772 306542
rect 296720 306478 296772 306484
rect 296536 306196 296588 306202
rect 296536 306138 296588 306144
rect 296352 306128 296404 306134
rect 296352 306070 296404 306076
rect 296168 304224 296220 304230
rect 296168 304166 296220 304172
rect 296732 295118 296760 306478
rect 296824 301714 296852 310406
rect 296904 306468 296956 306474
rect 296904 306410 296956 306416
rect 296812 301708 296864 301714
rect 296812 301650 296864 301656
rect 296916 295186 296944 306410
rect 297008 295322 297036 310420
rect 297192 306542 297220 310420
rect 297180 306536 297232 306542
rect 297180 306478 297232 306484
rect 297376 306474 297404 310420
rect 297364 306468 297416 306474
rect 297364 306410 297416 306416
rect 297560 306354 297588 310420
rect 297100 306326 297588 306354
rect 296996 295316 297048 295322
rect 296996 295258 297048 295264
rect 297100 295254 297128 306326
rect 297180 306264 297232 306270
rect 297180 306206 297232 306212
rect 297088 295248 297140 295254
rect 297088 295190 297140 295196
rect 296904 295180 296956 295186
rect 296904 295122 296956 295128
rect 296720 295112 296772 295118
rect 296720 295054 296772 295060
rect 295892 294500 295944 294506
rect 295892 294442 295944 294448
rect 287518 250472 287574 250481
rect 287518 250407 287574 250416
rect 284760 248124 284812 248130
rect 284760 248066 284812 248072
rect 283380 245336 283432 245342
rect 283380 245278 283432 245284
rect 280712 245268 280764 245274
rect 280712 245210 280764 245216
rect 279240 245200 279292 245206
rect 279240 245142 279292 245148
rect 269672 245132 269724 245138
rect 269672 245074 269724 245080
rect 268292 245064 268344 245070
rect 268292 245006 268344 245012
rect 262680 244996 262732 245002
rect 262680 244938 262732 244944
rect 257252 244928 257304 244934
rect 257252 244870 257304 244876
rect 297192 243642 297220 306206
rect 297744 296714 297772 310420
rect 297928 306270 297956 310420
rect 298112 306490 298140 310420
rect 298296 306626 298324 310420
rect 298480 308417 298508 310420
rect 298466 308408 298522 308417
rect 298466 308343 298522 308352
rect 298296 306598 298416 306626
rect 298112 306462 298324 306490
rect 298100 306332 298152 306338
rect 298100 306274 298152 306280
rect 297916 306264 297968 306270
rect 297916 306206 297968 306212
rect 297284 296686 297772 296714
rect 219348 243636 219400 243642
rect 219348 243578 219400 243584
rect 297180 243636 297232 243642
rect 297180 243578 297232 243584
rect 219256 155440 219308 155446
rect 219256 155382 219308 155388
rect 218796 155304 218848 155310
rect 218796 155246 218848 155252
rect 217876 155032 217928 155038
rect 217876 154974 217928 154980
rect 218058 3632 218114 3641
rect 216588 3596 216640 3602
rect 218058 3567 218114 3576
rect 216588 3538 216640 3544
rect 216862 3496 216918 3505
rect 216862 3431 216918 3440
rect 216496 3256 216548 3262
rect 216496 3198 216548 3204
rect 216876 480 216904 3431
rect 218072 480 218100 3567
rect 219360 3534 219388 243578
rect 297284 243574 297312 296686
rect 297272 243568 297324 243574
rect 298112 243545 298140 306274
rect 298192 305652 298244 305658
rect 298192 305594 298244 305600
rect 298204 243710 298232 305594
rect 298296 303385 298324 306462
rect 298282 303376 298338 303385
rect 298282 303311 298338 303320
rect 298388 303006 298416 306598
rect 298664 306338 298692 310420
rect 298652 306332 298704 306338
rect 298652 306274 298704 306280
rect 298376 303000 298428 303006
rect 298376 302942 298428 302948
rect 298848 302938 298876 310420
rect 298836 302932 298888 302938
rect 298836 302874 298888 302880
rect 299032 302234 299060 310420
rect 299216 305658 299244 310420
rect 299400 305969 299428 310420
rect 299492 310406 299690 310434
rect 299386 305960 299442 305969
rect 299386 305895 299442 305904
rect 299204 305652 299256 305658
rect 299204 305594 299256 305600
rect 298296 302206 299060 302234
rect 298296 300626 298324 302206
rect 298284 300620 298336 300626
rect 298284 300562 298336 300568
rect 298192 243704 298244 243710
rect 298192 243646 298244 243652
rect 299492 243642 299520 310406
rect 299664 306400 299716 306406
rect 299664 306342 299716 306348
rect 299572 306332 299624 306338
rect 299572 306274 299624 306280
rect 299480 243636 299532 243642
rect 299480 243578 299532 243584
rect 299584 243574 299612 306274
rect 299676 243846 299704 306342
rect 299860 306320 299888 310420
rect 299768 306292 299888 306320
rect 299664 243840 299716 243846
rect 299664 243782 299716 243788
rect 299768 243778 299796 306292
rect 299940 304428 299992 304434
rect 299940 304370 299992 304376
rect 299848 303204 299900 303210
rect 299848 303146 299900 303152
rect 299860 300558 299888 303146
rect 299848 300552 299900 300558
rect 299848 300494 299900 300500
rect 299952 300422 299980 304370
rect 299940 300416 299992 300422
rect 299940 300358 299992 300364
rect 300044 300121 300072 310420
rect 300228 306338 300256 310420
rect 300412 306406 300440 310420
rect 300400 306400 300452 306406
rect 300400 306342 300452 306348
rect 300216 306332 300268 306338
rect 300216 306274 300268 306280
rect 300596 303210 300624 310420
rect 300780 304434 300808 310420
rect 300964 306490 300992 310420
rect 301148 306762 301176 310420
rect 301332 308446 301360 310420
rect 301516 308514 301544 310420
rect 301504 308508 301556 308514
rect 301504 308450 301556 308456
rect 301320 308440 301372 308446
rect 301320 308382 301372 308388
rect 301148 306734 301360 306762
rect 300964 306462 301084 306490
rect 300860 306400 300912 306406
rect 301056 306388 301084 306462
rect 301056 306360 301176 306388
rect 300860 306342 300912 306348
rect 300768 304428 300820 304434
rect 300768 304370 300820 304376
rect 300584 303204 300636 303210
rect 300584 303146 300636 303152
rect 300030 300112 300086 300121
rect 300030 300047 300086 300056
rect 300872 246702 300900 306342
rect 300952 306264 301004 306270
rect 300952 306206 301004 306212
rect 300964 253706 300992 306206
rect 301044 306196 301096 306202
rect 301044 306138 301096 306144
rect 301056 253774 301084 306138
rect 301148 303074 301176 306360
rect 301136 303068 301188 303074
rect 301136 303010 301188 303016
rect 301332 302234 301360 306734
rect 301700 306406 301728 310420
rect 301688 306400 301740 306406
rect 301688 306342 301740 306348
rect 301884 306202 301912 310420
rect 302068 306270 302096 310420
rect 302344 308582 302372 310420
rect 302528 308650 302556 310420
rect 302516 308644 302568 308650
rect 302516 308586 302568 308592
rect 302332 308576 302384 308582
rect 302332 308518 302384 308524
rect 302712 306490 302740 310420
rect 302252 306462 302740 306490
rect 302056 306264 302108 306270
rect 302056 306206 302108 306212
rect 301872 306196 301924 306202
rect 301872 306138 301924 306144
rect 301148 302206 301360 302234
rect 301148 300490 301176 302206
rect 301136 300484 301188 300490
rect 301136 300426 301188 300432
rect 301044 253768 301096 253774
rect 301044 253710 301096 253716
rect 300952 253700 301004 253706
rect 300952 253642 301004 253648
rect 302252 248062 302280 306462
rect 302424 306400 302476 306406
rect 302424 306342 302476 306348
rect 302332 306264 302384 306270
rect 302332 306206 302384 306212
rect 302344 248130 302372 306206
rect 302436 250850 302464 306342
rect 302516 306332 302568 306338
rect 302516 306274 302568 306280
rect 302528 253162 302556 306274
rect 302896 296714 302924 310420
rect 303080 306338 303108 310420
rect 303264 306406 303292 310420
rect 303252 306400 303304 306406
rect 303252 306342 303304 306348
rect 303068 306332 303120 306338
rect 303068 306274 303120 306280
rect 303448 306270 303476 310420
rect 303436 306264 303488 306270
rect 303436 306206 303488 306212
rect 302620 296686 302924 296714
rect 302516 253156 302568 253162
rect 302516 253098 302568 253104
rect 302620 253094 302648 296686
rect 302608 253088 302660 253094
rect 302608 253030 302660 253036
rect 302424 250844 302476 250850
rect 302424 250786 302476 250792
rect 302332 248124 302384 248130
rect 302332 248066 302384 248072
rect 302240 248056 302292 248062
rect 302240 247998 302292 248004
rect 300860 246696 300912 246702
rect 300860 246638 300912 246644
rect 303632 243914 303660 310420
rect 303816 308786 303844 310420
rect 303804 308780 303856 308786
rect 303804 308722 303856 308728
rect 303804 306400 303856 306406
rect 303804 306342 303856 306348
rect 303712 306332 303764 306338
rect 303712 306274 303764 306280
rect 303724 244905 303752 306274
rect 303816 250617 303844 306342
rect 304000 306202 304028 310420
rect 303988 306196 304040 306202
rect 303988 306138 304040 306144
rect 303988 305992 304040 305998
rect 303988 305934 304040 305940
rect 303896 304292 303948 304298
rect 303896 304234 303948 304240
rect 303908 253842 303936 304234
rect 304000 253910 304028 305934
rect 304184 304298 304212 310420
rect 304368 306338 304396 310420
rect 304552 308718 304580 310420
rect 304644 310406 304842 310434
rect 304540 308712 304592 308718
rect 304540 308654 304592 308660
rect 304644 306406 304672 310406
rect 304632 306400 304684 306406
rect 304632 306342 304684 306348
rect 304356 306332 304408 306338
rect 304356 306274 304408 306280
rect 305012 306218 305040 310420
rect 305196 306354 305224 310420
rect 305380 306354 305408 310420
rect 305564 306490 305592 310420
rect 305564 306462 305684 306490
rect 305196 306326 305316 306354
rect 305380 306326 305592 306354
rect 305012 306190 305224 306218
rect 305000 306128 305052 306134
rect 305000 306070 305052 306076
rect 304172 304292 304224 304298
rect 304172 304234 304224 304240
rect 303988 253904 304040 253910
rect 303988 253846 304040 253852
rect 303896 253836 303948 253842
rect 303896 253778 303948 253784
rect 303802 250608 303858 250617
rect 303802 250543 303858 250552
rect 305012 245041 305040 306070
rect 305092 306060 305144 306066
rect 305092 306002 305144 306008
rect 305104 248198 305132 306002
rect 305092 248192 305144 248198
rect 305092 248134 305144 248140
rect 305196 245177 305224 306190
rect 305288 248033 305316 306326
rect 305460 306264 305512 306270
rect 305460 306206 305512 306212
rect 305368 306196 305420 306202
rect 305368 306138 305420 306144
rect 305380 248334 305408 306138
rect 305472 250918 305500 306206
rect 305460 250912 305512 250918
rect 305460 250854 305512 250860
rect 305564 250753 305592 306326
rect 305656 306134 305684 306462
rect 305748 306202 305776 310420
rect 305932 306270 305960 310420
rect 306116 308553 306144 310420
rect 306102 308544 306158 308553
rect 306102 308479 306158 308488
rect 305920 306264 305972 306270
rect 305920 306206 305972 306212
rect 305736 306196 305788 306202
rect 305736 306138 305788 306144
rect 305644 306128 305696 306134
rect 305644 306070 305696 306076
rect 306300 306066 306328 310420
rect 306484 306490 306512 310420
rect 306392 306462 306512 306490
rect 306392 306202 306420 306462
rect 306668 306354 306696 310420
rect 306852 306474 306880 310420
rect 306840 306468 306892 306474
rect 306840 306410 306892 306416
rect 307036 306354 307064 310420
rect 306484 306326 306696 306354
rect 306760 306326 307064 306354
rect 306380 306196 306432 306202
rect 306380 306138 306432 306144
rect 306288 306060 306340 306066
rect 306288 306002 306340 306008
rect 306380 306060 306432 306066
rect 306380 306002 306432 306008
rect 305550 250744 305606 250753
rect 305550 250679 305606 250688
rect 305368 248328 305420 248334
rect 305368 248270 305420 248276
rect 305274 248024 305330 248033
rect 305274 247959 305330 247968
rect 306392 245274 306420 306002
rect 306484 245449 306512 306326
rect 306656 306264 306708 306270
rect 306656 306206 306708 306212
rect 306564 306128 306616 306134
rect 306564 306070 306616 306076
rect 306576 247625 306604 306070
rect 306668 248266 306696 306206
rect 306760 251122 306788 306326
rect 306840 306196 306892 306202
rect 306840 306138 306892 306144
rect 306748 251116 306800 251122
rect 306748 251058 306800 251064
rect 306852 251054 306880 306138
rect 307220 306066 307248 310420
rect 307312 310406 307510 310434
rect 307312 306134 307340 310406
rect 307300 306128 307352 306134
rect 307300 306070 307352 306076
rect 307208 306060 307260 306066
rect 307208 306002 307260 306008
rect 307680 296714 307708 310420
rect 307864 306354 307892 310420
rect 306944 296686 307708 296714
rect 307772 306326 307892 306354
rect 308048 306354 308076 310420
rect 307944 306332 307996 306338
rect 306840 251048 306892 251054
rect 306840 250990 306892 250996
rect 306944 250782 306972 296686
rect 306932 250776 306984 250782
rect 306932 250718 306984 250724
rect 306656 248260 306708 248266
rect 306656 248202 306708 248208
rect 306562 247616 306618 247625
rect 306562 247551 306618 247560
rect 306470 245440 306526 245449
rect 306470 245375 306526 245384
rect 307772 245342 307800 306326
rect 308048 306326 308168 306354
rect 307944 306274 307996 306280
rect 307852 306196 307904 306202
rect 307852 306138 307904 306144
rect 307864 245478 307892 306138
rect 307852 245472 307904 245478
rect 307852 245414 307904 245420
rect 307956 245410 307984 306274
rect 308036 306264 308088 306270
rect 308036 306206 308088 306212
rect 308048 247761 308076 306206
rect 308140 248402 308168 306326
rect 308232 250986 308260 310420
rect 308416 306202 308444 310420
rect 308600 306270 308628 310420
rect 308588 306264 308640 306270
rect 308588 306206 308640 306212
rect 308404 306196 308456 306202
rect 308404 306138 308456 306144
rect 308784 296714 308812 310420
rect 308968 306338 308996 310420
rect 308956 306332 309008 306338
rect 308956 306274 309008 306280
rect 309152 306218 309180 310420
rect 309336 306354 309364 310420
rect 309520 306490 309548 310420
rect 309520 306462 309640 306490
rect 309336 306326 309548 306354
rect 309152 306190 309456 306218
rect 309232 306128 309284 306134
rect 309232 306070 309284 306076
rect 309140 306060 309192 306066
rect 309140 306002 309192 306008
rect 308324 296686 308812 296714
rect 308220 250980 308272 250986
rect 308220 250922 308272 250928
rect 308324 250481 308352 296686
rect 308310 250472 308366 250481
rect 308310 250407 308366 250416
rect 308128 248396 308180 248402
rect 308128 248338 308180 248344
rect 308034 247752 308090 247761
rect 308034 247687 308090 247696
rect 307944 245404 307996 245410
rect 307944 245346 307996 245352
rect 307760 245336 307812 245342
rect 309152 245313 309180 306002
rect 309244 247897 309272 306070
rect 309324 305516 309376 305522
rect 309324 305458 309376 305464
rect 309230 247888 309286 247897
rect 309230 247823 309286 247832
rect 309336 245585 309364 305458
rect 309428 247654 309456 306190
rect 309520 250442 309548 306326
rect 309612 306066 309640 306462
rect 309704 306134 309732 310420
rect 309796 310406 309994 310434
rect 309692 306128 309744 306134
rect 309692 306070 309744 306076
rect 309600 306060 309652 306066
rect 309600 306002 309652 306008
rect 309796 296714 309824 310406
rect 310164 305522 310192 310420
rect 310348 308922 310376 310420
rect 310336 308916 310388 308922
rect 310336 308858 310388 308864
rect 310152 305516 310204 305522
rect 310152 305458 310204 305464
rect 309612 296686 309824 296714
rect 309612 251190 309640 296686
rect 309600 251184 309652 251190
rect 309600 251126 309652 251132
rect 309508 250436 309560 250442
rect 309508 250378 309560 250384
rect 309416 247648 309468 247654
rect 309416 247590 309468 247596
rect 309322 245576 309378 245585
rect 309322 245511 309378 245520
rect 307760 245278 307812 245284
rect 309138 245304 309194 245313
rect 306380 245268 306432 245274
rect 309138 245239 309194 245248
rect 306380 245210 306432 245216
rect 305182 245168 305238 245177
rect 305182 245103 305238 245112
rect 304998 245032 305054 245041
rect 304998 244967 305054 244976
rect 303710 244896 303766 244905
rect 303710 244831 303766 244840
rect 310532 244769 310560 310420
rect 310612 306468 310664 306474
rect 310612 306410 310664 306416
rect 310624 248169 310652 306410
rect 310716 306354 310744 310420
rect 310900 306474 310928 310420
rect 310888 306468 310940 306474
rect 310888 306410 310940 306416
rect 311084 306354 311112 310420
rect 311268 306490 311296 310420
rect 311268 306462 311388 306490
rect 310716 306326 310928 306354
rect 310704 306196 310756 306202
rect 310704 306138 310756 306144
rect 310716 250889 310744 306138
rect 310796 306128 310848 306134
rect 310796 306070 310848 306076
rect 310808 251841 310836 306070
rect 310794 251832 310850 251841
rect 310794 251767 310850 251776
rect 310900 251025 310928 306326
rect 310980 306332 311032 306338
rect 311084 306326 311296 306354
rect 310980 306274 311032 306280
rect 310992 254561 311020 306274
rect 311072 306264 311124 306270
rect 311072 306206 311124 306212
rect 311084 260137 311112 306206
rect 311268 260273 311296 306326
rect 311360 306202 311388 306462
rect 311452 306338 311480 310420
rect 311440 306332 311492 306338
rect 311440 306274 311492 306280
rect 311636 306270 311664 310420
rect 311624 306264 311676 306270
rect 311624 306206 311676 306212
rect 311348 306196 311400 306202
rect 311348 306138 311400 306144
rect 311820 306134 311848 310420
rect 311900 308236 311952 308242
rect 311900 308178 311952 308184
rect 311808 306128 311860 306134
rect 311808 306070 311860 306076
rect 311254 260264 311310 260273
rect 311254 260199 311310 260208
rect 311070 260128 311126 260137
rect 311070 260063 311126 260072
rect 310978 254552 311034 254561
rect 310978 254487 311034 254496
rect 310886 251016 310942 251025
rect 310886 250951 310942 250960
rect 310702 250880 310758 250889
rect 310702 250815 310758 250824
rect 311912 250714 311940 308178
rect 312004 308174 312032 310420
rect 312188 308394 312216 310420
rect 312096 308366 312216 308394
rect 312268 308372 312320 308378
rect 311992 308168 312044 308174
rect 311992 308110 312044 308116
rect 311992 308032 312044 308038
rect 311992 307974 312044 307980
rect 312004 254862 312032 307974
rect 312096 280809 312124 308366
rect 312268 308314 312320 308320
rect 312176 308304 312228 308310
rect 312176 308246 312228 308252
rect 312188 286618 312216 308246
rect 312280 301714 312308 308314
rect 312372 303521 312400 310420
rect 312464 310406 312662 310434
rect 312464 308310 312492 310406
rect 312452 308304 312504 308310
rect 312452 308246 312504 308252
rect 312452 308168 312504 308174
rect 312452 308110 312504 308116
rect 312464 306105 312492 308110
rect 312832 308038 312860 310420
rect 313016 308378 313044 310420
rect 313004 308372 313056 308378
rect 313004 308314 313056 308320
rect 313200 308242 313228 310420
rect 313384 308394 313412 310420
rect 313384 308366 313504 308394
rect 313372 308304 313424 308310
rect 313372 308246 313424 308252
rect 313188 308236 313240 308242
rect 313188 308178 313240 308184
rect 313280 308236 313332 308242
rect 313280 308178 313332 308184
rect 312820 308032 312872 308038
rect 312820 307974 312872 307980
rect 312450 306096 312506 306105
rect 312450 306031 312506 306040
rect 312358 303512 312414 303521
rect 312358 303447 312414 303456
rect 312268 301708 312320 301714
rect 312268 301650 312320 301656
rect 312176 286612 312228 286618
rect 312176 286554 312228 286560
rect 312082 280800 312138 280809
rect 312082 280735 312138 280744
rect 313292 264382 313320 308178
rect 313384 265577 313412 308246
rect 313476 282470 313504 308366
rect 313568 307290 313596 310420
rect 313752 308394 313780 310420
rect 313660 308366 313780 308394
rect 313936 308378 313964 310420
rect 313924 308372 313976 308378
rect 313556 307284 313608 307290
rect 313556 307226 313608 307232
rect 313556 307148 313608 307154
rect 313556 307090 313608 307096
rect 313568 285122 313596 307090
rect 313660 285190 313688 308366
rect 313924 308314 313976 308320
rect 314120 308258 314148 310420
rect 313752 308230 314148 308258
rect 314304 308242 314332 310420
rect 314292 308236 314344 308242
rect 313752 294778 313780 308230
rect 314292 308178 314344 308184
rect 313832 307284 313884 307290
rect 313832 307226 313884 307232
rect 313844 300694 313872 307226
rect 314488 307154 314516 310420
rect 314672 308854 314700 310420
rect 314870 310406 314976 310434
rect 314844 308984 314896 308990
rect 314844 308926 314896 308932
rect 314660 308848 314712 308854
rect 314660 308790 314712 308796
rect 314752 308304 314804 308310
rect 314752 308246 314804 308252
rect 314660 308236 314712 308242
rect 314660 308178 314712 308184
rect 314476 307148 314528 307154
rect 314476 307090 314528 307096
rect 313832 300688 313884 300694
rect 313832 300630 313884 300636
rect 313740 294772 313792 294778
rect 313740 294714 313792 294720
rect 313648 285184 313700 285190
rect 313648 285126 313700 285132
rect 313556 285116 313608 285122
rect 313556 285058 313608 285064
rect 313464 282464 313516 282470
rect 313464 282406 313516 282412
rect 313370 265568 313426 265577
rect 313370 265503 313426 265512
rect 313280 264376 313332 264382
rect 313280 264318 313332 264324
rect 314672 263022 314700 308178
rect 314764 270026 314792 308246
rect 314856 271318 314884 308926
rect 314948 308802 314976 310406
rect 315040 310406 315146 310434
rect 315040 308990 315068 310406
rect 315028 308984 315080 308990
rect 315028 308926 315080 308932
rect 314948 308774 315160 308802
rect 314936 308372 314988 308378
rect 314936 308314 314988 308320
rect 314948 283898 314976 308314
rect 315028 308168 315080 308174
rect 315028 308110 315080 308116
rect 315040 292058 315068 308110
rect 315132 298926 315160 308774
rect 315316 308174 315344 310420
rect 315396 308848 315448 308854
rect 315396 308790 315448 308796
rect 315304 308168 315356 308174
rect 315304 308110 315356 308116
rect 315408 307358 315436 308790
rect 315500 308242 315528 310420
rect 315684 308310 315712 310420
rect 315868 308378 315896 310420
rect 315948 309460 316000 309466
rect 315948 309402 316000 309408
rect 315960 309134 315988 309402
rect 316052 309210 316080 310420
rect 316236 309346 316264 310420
rect 316420 309466 316448 310420
rect 316408 309460 316460 309466
rect 316408 309402 316460 309408
rect 316236 309318 316540 309346
rect 316052 309182 316264 309210
rect 315960 309106 316080 309134
rect 315856 308372 315908 308378
rect 315856 308314 315908 308320
rect 315672 308304 315724 308310
rect 315672 308246 315724 308252
rect 315488 308236 315540 308242
rect 315488 308178 315540 308184
rect 315396 307352 315448 307358
rect 315396 307294 315448 307300
rect 315120 298920 315172 298926
rect 315120 298862 315172 298868
rect 315028 292052 315080 292058
rect 315028 291994 315080 292000
rect 314936 283892 314988 283898
rect 314936 283834 314988 283840
rect 314844 271312 314896 271318
rect 314844 271254 314896 271260
rect 314752 270020 314804 270026
rect 314752 269962 314804 269968
rect 314660 263016 314712 263022
rect 314660 262958 314712 262964
rect 311992 254856 312044 254862
rect 311992 254798 312044 254804
rect 316052 253638 316080 309106
rect 316132 308372 316184 308378
rect 316132 308314 316184 308320
rect 316040 253632 316092 253638
rect 316040 253574 316092 253580
rect 316144 253570 316172 308314
rect 316236 308292 316264 309182
rect 316236 308264 316356 308292
rect 316224 308168 316276 308174
rect 316224 308110 316276 308116
rect 316236 257378 316264 308110
rect 316328 257446 316356 308264
rect 316512 308156 316540 309318
rect 316604 308310 316632 310420
rect 316592 308304 316644 308310
rect 316592 308246 316644 308252
rect 316512 308128 316632 308156
rect 316500 308032 316552 308038
rect 316500 307974 316552 307980
rect 316408 307080 316460 307086
rect 316408 307022 316460 307028
rect 316420 258806 316448 307022
rect 316512 261730 316540 307974
rect 316604 261798 316632 308128
rect 316788 308038 316816 310420
rect 316972 308378 317000 310420
rect 316960 308372 317012 308378
rect 316960 308314 317012 308320
rect 316776 308032 316828 308038
rect 316776 307974 316828 307980
rect 317156 307086 317184 310420
rect 317340 308242 317368 310420
rect 317538 310406 317736 310434
rect 317420 308916 317472 308922
rect 317420 308858 317472 308864
rect 317328 308236 317380 308242
rect 317328 308178 317380 308184
rect 317144 307080 317196 307086
rect 317144 307022 317196 307028
rect 316592 261792 316644 261798
rect 316592 261734 316644 261740
rect 316500 261724 316552 261730
rect 316500 261666 316552 261672
rect 316408 258800 316460 258806
rect 316408 258742 316460 258748
rect 316316 257440 316368 257446
rect 316316 257382 316368 257388
rect 316224 257372 316276 257378
rect 316224 257314 316276 257320
rect 317432 254794 317460 308858
rect 317604 308372 317656 308378
rect 317604 308314 317656 308320
rect 317512 308100 317564 308106
rect 317512 308042 317564 308048
rect 317524 275534 317552 308042
rect 317616 276894 317644 308314
rect 317708 308310 317736 310406
rect 317800 308530 317828 310420
rect 317984 308922 318012 310420
rect 317972 308916 318024 308922
rect 317972 308858 318024 308864
rect 317800 308502 318012 308530
rect 317696 308304 317748 308310
rect 317696 308246 317748 308252
rect 317880 308304 317932 308310
rect 317880 308246 317932 308252
rect 317696 308168 317748 308174
rect 317696 308110 317748 308116
rect 317708 290766 317736 308110
rect 317788 307964 317840 307970
rect 317788 307906 317840 307912
rect 317800 293554 317828 307906
rect 317892 303249 317920 308246
rect 317984 307290 318012 308502
rect 318064 308236 318116 308242
rect 318064 308178 318116 308184
rect 317972 307284 318024 307290
rect 317972 307226 318024 307232
rect 317878 303240 317934 303249
rect 317878 303175 317934 303184
rect 318076 296206 318104 308178
rect 318168 307970 318196 310420
rect 318352 308378 318380 310420
rect 318340 308372 318392 308378
rect 318340 308314 318392 308320
rect 318536 308106 318564 310420
rect 318720 308174 318748 310420
rect 318904 308394 318932 310420
rect 319088 308922 319116 310420
rect 319076 308916 319128 308922
rect 319076 308858 319128 308864
rect 318904 308366 319116 308394
rect 318984 308304 319036 308310
rect 318984 308246 319036 308252
rect 318800 308236 318852 308242
rect 318800 308178 318852 308184
rect 318708 308168 318760 308174
rect 318708 308110 318760 308116
rect 318524 308100 318576 308106
rect 318524 308042 318576 308048
rect 318156 307964 318208 307970
rect 318156 307906 318208 307912
rect 318064 296200 318116 296206
rect 318064 296142 318116 296148
rect 317788 293548 317840 293554
rect 317788 293490 317840 293496
rect 317696 290760 317748 290766
rect 317696 290702 317748 290708
rect 317604 276888 317656 276894
rect 317604 276830 317656 276836
rect 317512 275528 317564 275534
rect 317512 275470 317564 275476
rect 317420 254788 317472 254794
rect 317420 254730 317472 254736
rect 316132 253564 316184 253570
rect 316132 253506 316184 253512
rect 311900 250708 311952 250714
rect 311900 250650 311952 250656
rect 318812 249354 318840 308178
rect 318892 308168 318944 308174
rect 318892 308110 318944 308116
rect 318904 250646 318932 308110
rect 318996 256222 319024 308246
rect 319088 279682 319116 308366
rect 319168 308372 319220 308378
rect 319168 308314 319220 308320
rect 319180 282402 319208 308314
rect 319272 297634 319300 310420
rect 319352 308916 319404 308922
rect 319352 308858 319404 308864
rect 319364 298994 319392 308858
rect 319456 308242 319484 310420
rect 319640 308310 319668 310420
rect 319824 308378 319852 310420
rect 319812 308372 319864 308378
rect 319812 308314 319864 308320
rect 319628 308304 319680 308310
rect 319628 308246 319680 308252
rect 319444 308236 319496 308242
rect 319444 308178 319496 308184
rect 320008 308174 320036 310420
rect 320180 308372 320232 308378
rect 320180 308314 320232 308320
rect 319996 308168 320048 308174
rect 319996 308110 320048 308116
rect 319352 298988 319404 298994
rect 319352 298930 319404 298936
rect 319260 297628 319312 297634
rect 319260 297570 319312 297576
rect 319168 282396 319220 282402
rect 319168 282338 319220 282344
rect 319076 279676 319128 279682
rect 319076 279618 319128 279624
rect 318984 256216 319036 256222
rect 318984 256158 319036 256164
rect 318892 250640 318944 250646
rect 318892 250582 318944 250588
rect 318800 249348 318852 249354
rect 318800 249290 318852 249296
rect 310610 248160 310666 248169
rect 310610 248095 310666 248104
rect 320192 247994 320220 308314
rect 320284 308174 320312 310420
rect 320364 308304 320416 308310
rect 320364 308246 320416 308252
rect 320272 308168 320324 308174
rect 320272 308110 320324 308116
rect 320272 308032 320324 308038
rect 320272 307974 320324 307980
rect 320284 256154 320312 307974
rect 320376 264314 320404 308246
rect 320468 308156 320496 310420
rect 320652 308310 320680 310420
rect 320640 308304 320692 308310
rect 320640 308246 320692 308252
rect 320640 308168 320692 308174
rect 320468 308128 320588 308156
rect 320456 307964 320508 307970
rect 320456 307906 320508 307912
rect 320468 279614 320496 307906
rect 320560 281042 320588 308128
rect 320640 308110 320692 308116
rect 320652 290630 320680 308110
rect 320836 300354 320864 310420
rect 321020 307970 321048 310420
rect 321204 308378 321232 310420
rect 321192 308372 321244 308378
rect 321192 308314 321244 308320
rect 321388 308038 321416 310420
rect 321376 308032 321428 308038
rect 321376 307974 321428 307980
rect 321008 307964 321060 307970
rect 321008 307906 321060 307912
rect 321572 306270 321600 310420
rect 321756 306354 321784 310420
rect 321836 307012 321888 307018
rect 321836 306954 321888 306960
rect 321848 306456 321876 306954
rect 321940 306592 321968 310420
rect 322124 307018 322152 310420
rect 322112 307012 322164 307018
rect 322112 306954 322164 306960
rect 321940 306564 322152 306592
rect 321848 306428 321968 306456
rect 321664 306326 321784 306354
rect 321836 306332 321888 306338
rect 321560 306264 321612 306270
rect 321560 306206 321612 306212
rect 321560 306128 321612 306134
rect 321560 306070 321612 306076
rect 320824 300348 320876 300354
rect 320824 300290 320876 300296
rect 320640 290624 320692 290630
rect 320640 290566 320692 290572
rect 320548 281036 320600 281042
rect 320548 280978 320600 280984
rect 320456 279608 320508 279614
rect 320456 279550 320508 279556
rect 320364 264308 320416 264314
rect 320364 264250 320416 264256
rect 320272 256148 320324 256154
rect 320272 256090 320324 256096
rect 321572 252142 321600 306070
rect 321664 252210 321692 306326
rect 321836 306274 321888 306280
rect 321744 306196 321796 306202
rect 321744 306138 321796 306144
rect 321756 256086 321784 306138
rect 321848 278254 321876 306274
rect 321940 289270 321968 306428
rect 322020 306264 322072 306270
rect 322020 306206 322072 306212
rect 322032 296138 322060 306206
rect 322124 299474 322152 306564
rect 322308 306134 322336 310420
rect 322492 306202 322520 310420
rect 322676 306338 322704 310420
rect 322952 306354 322980 310420
rect 322664 306332 322716 306338
rect 322952 306326 323072 306354
rect 322664 306274 322716 306280
rect 322940 306264 322992 306270
rect 322940 306206 322992 306212
rect 322480 306196 322532 306202
rect 322480 306138 322532 306144
rect 322296 306128 322348 306134
rect 322296 306070 322348 306076
rect 322124 299446 322244 299474
rect 322216 297702 322244 299446
rect 322204 297696 322256 297702
rect 322204 297638 322256 297644
rect 322020 296132 322072 296138
rect 322020 296074 322072 296080
rect 321928 289264 321980 289270
rect 321928 289206 321980 289212
rect 321836 278248 321888 278254
rect 321836 278190 321888 278196
rect 321744 256080 321796 256086
rect 321744 256022 321796 256028
rect 321652 252204 321704 252210
rect 321652 252146 321704 252152
rect 321560 252136 321612 252142
rect 321560 252078 321612 252084
rect 320180 247988 320232 247994
rect 320180 247930 320232 247936
rect 322952 246634 322980 306206
rect 323044 262954 323072 306326
rect 323136 306218 323164 310420
rect 323320 306354 323348 310420
rect 323320 306326 323440 306354
rect 323136 306190 323348 306218
rect 323216 306128 323268 306134
rect 323216 306070 323268 306076
rect 323124 306060 323176 306066
rect 323124 306002 323176 306008
rect 323136 276826 323164 306002
rect 323228 278186 323256 306070
rect 323320 285054 323348 306190
rect 323412 286550 323440 306326
rect 323504 306270 323532 310420
rect 323688 307222 323716 310420
rect 323676 307216 323728 307222
rect 323676 307158 323728 307164
rect 323492 306264 323544 306270
rect 323492 306206 323544 306212
rect 323872 306066 323900 310420
rect 324056 306134 324084 310420
rect 324044 306128 324096 306134
rect 324044 306070 324096 306076
rect 323860 306060 323912 306066
rect 323860 306002 323912 306008
rect 324240 304502 324268 310420
rect 324424 306746 324452 310420
rect 324412 306740 324464 306746
rect 324412 306682 324464 306688
rect 324608 306626 324636 310420
rect 324332 306598 324636 306626
rect 324228 304496 324280 304502
rect 324228 304438 324280 304444
rect 323400 286544 323452 286550
rect 323400 286486 323452 286492
rect 323308 285048 323360 285054
rect 323308 284990 323360 284996
rect 323216 278180 323268 278186
rect 323216 278122 323268 278128
rect 323124 276820 323176 276826
rect 323124 276762 323176 276768
rect 323032 262948 323084 262954
rect 323032 262890 323084 262896
rect 322940 246628 322992 246634
rect 322940 246570 322992 246576
rect 324332 245206 324360 306598
rect 324792 306490 324820 310420
rect 324516 306462 324820 306490
rect 324516 306218 324544 306462
rect 324976 306354 325004 310420
rect 325056 306740 325108 306746
rect 325056 306682 325108 306688
rect 324424 306190 324544 306218
rect 324700 306326 325004 306354
rect 324596 306196 324648 306202
rect 324424 256018 324452 306190
rect 324596 306138 324648 306144
rect 324504 306128 324556 306134
rect 324504 306070 324556 306076
rect 324516 274174 324544 306070
rect 324608 274242 324636 306138
rect 324700 275466 324728 306326
rect 325068 302234 325096 306682
rect 324792 302206 325096 302234
rect 324792 283762 324820 302206
rect 325160 296714 325188 310420
rect 325252 310406 325450 310434
rect 325252 306134 325280 310406
rect 325620 306202 325648 310420
rect 325804 306474 325832 310420
rect 325792 306468 325844 306474
rect 325792 306410 325844 306416
rect 325988 306354 326016 310420
rect 325700 306332 325752 306338
rect 325700 306274 325752 306280
rect 325804 306326 326016 306354
rect 326172 306338 326200 310420
rect 326160 306332 326212 306338
rect 325608 306196 325660 306202
rect 325608 306138 325660 306144
rect 325240 306128 325292 306134
rect 325240 306070 325292 306076
rect 324884 296686 325188 296714
rect 324884 286482 324912 296686
rect 324872 286476 324924 286482
rect 324872 286418 324924 286424
rect 324780 283756 324832 283762
rect 324780 283698 324832 283704
rect 324688 275460 324740 275466
rect 324688 275402 324740 275408
rect 324596 274236 324648 274242
rect 324596 274178 324648 274184
rect 324504 274168 324556 274174
rect 324504 274110 324556 274116
rect 324412 256012 324464 256018
rect 324412 255954 324464 255960
rect 325712 247926 325740 306274
rect 325804 252006 325832 306326
rect 326160 306274 326212 306280
rect 325884 306264 325936 306270
rect 325884 306206 325936 306212
rect 325896 274106 325924 306206
rect 326356 306082 326384 310420
rect 326436 306468 326488 306474
rect 326436 306410 326488 306416
rect 325988 306054 326384 306082
rect 325988 275398 326016 306054
rect 326448 304434 326476 306410
rect 326436 304428 326488 304434
rect 326436 304370 326488 304376
rect 326540 302234 326568 310420
rect 326724 308990 326752 310420
rect 326712 308984 326764 308990
rect 326712 308926 326764 308932
rect 326908 306270 326936 310420
rect 326896 306264 326948 306270
rect 326896 306206 326948 306212
rect 326080 302206 326568 302234
rect 326080 280974 326108 302206
rect 326068 280968 326120 280974
rect 326068 280910 326120 280916
rect 325976 275392 326028 275398
rect 325976 275334 326028 275340
rect 325884 274100 325936 274106
rect 325884 274042 325936 274048
rect 325792 252000 325844 252006
rect 325792 251942 325844 251948
rect 327092 249218 327120 310420
rect 327172 306604 327224 306610
rect 327172 306546 327224 306552
rect 327184 306218 327212 306546
rect 327276 306354 327304 310420
rect 327460 306490 327488 310420
rect 327644 306610 327672 310420
rect 327632 306604 327684 306610
rect 327632 306546 327684 306552
rect 327460 306462 327672 306490
rect 327276 306326 327488 306354
rect 327184 306190 327396 306218
rect 327172 306128 327224 306134
rect 327172 306070 327224 306076
rect 327184 251938 327212 306070
rect 327264 306060 327316 306066
rect 327264 306002 327316 306008
rect 327276 268462 327304 306002
rect 327368 282334 327396 306190
rect 327460 287842 327488 306326
rect 327540 306332 327592 306338
rect 327540 306274 327592 306280
rect 327552 291990 327580 306274
rect 327644 297498 327672 306462
rect 327828 306338 327856 310420
rect 327920 310406 328118 310434
rect 327816 306332 327868 306338
rect 327816 306274 327868 306280
rect 327920 306134 327948 310406
rect 327908 306128 327960 306134
rect 327908 306070 327960 306076
rect 328288 306066 328316 310420
rect 328472 306134 328500 310420
rect 328552 306468 328604 306474
rect 328552 306410 328604 306416
rect 328460 306128 328512 306134
rect 328460 306070 328512 306076
rect 328276 306060 328328 306066
rect 328276 306002 328328 306008
rect 328460 305992 328512 305998
rect 328460 305934 328512 305940
rect 327632 297492 327684 297498
rect 327632 297434 327684 297440
rect 327540 291984 327592 291990
rect 327540 291926 327592 291932
rect 327448 287836 327500 287842
rect 327448 287778 327500 287784
rect 327356 282328 327408 282334
rect 327356 282270 327408 282276
rect 327264 268456 327316 268462
rect 327264 268398 327316 268404
rect 327172 251932 327224 251938
rect 327172 251874 327224 251880
rect 327080 249212 327132 249218
rect 327080 249154 327132 249160
rect 328472 249150 328500 305934
rect 328564 254726 328592 306410
rect 328656 306338 328684 310420
rect 328736 306400 328788 306406
rect 328736 306342 328788 306348
rect 328840 306354 328868 310420
rect 328644 306332 328696 306338
rect 328644 306274 328696 306280
rect 328644 306196 328696 306202
rect 328644 306138 328696 306144
rect 328656 268394 328684 306138
rect 328748 272610 328776 306342
rect 328840 306326 328960 306354
rect 328828 306264 328880 306270
rect 328828 306206 328880 306212
rect 328840 282266 328868 306206
rect 328932 286414 328960 306326
rect 329024 306270 329052 310420
rect 329104 306332 329156 306338
rect 329104 306274 329156 306280
rect 329012 306264 329064 306270
rect 329012 306206 329064 306212
rect 329012 306128 329064 306134
rect 329012 306070 329064 306076
rect 329024 293418 329052 306070
rect 329116 294710 329144 306274
rect 329208 306202 329236 310420
rect 329392 306474 329420 310420
rect 329380 306468 329432 306474
rect 329380 306410 329432 306416
rect 329576 306406 329604 310420
rect 329564 306400 329616 306406
rect 329564 306342 329616 306348
rect 329196 306196 329248 306202
rect 329196 306138 329248 306144
rect 329760 305998 329788 310420
rect 329944 308417 329972 310420
rect 329930 308408 329986 308417
rect 329930 308343 329986 308352
rect 330128 307154 330156 310420
rect 330116 307148 330168 307154
rect 330116 307090 330168 307096
rect 329840 306400 329892 306406
rect 330312 306354 330340 310420
rect 329840 306342 329892 306348
rect 329748 305992 329800 305998
rect 329748 305934 329800 305940
rect 329104 294704 329156 294710
rect 329104 294646 329156 294652
rect 329012 293412 329064 293418
rect 329012 293354 329064 293360
rect 328920 286408 328972 286414
rect 328920 286350 328972 286356
rect 328828 282260 328880 282266
rect 328828 282202 328880 282208
rect 328736 272604 328788 272610
rect 328736 272546 328788 272552
rect 328644 268388 328696 268394
rect 328644 268330 328696 268336
rect 329852 261594 329880 306342
rect 329932 306332 329984 306338
rect 329932 306274 329984 306280
rect 330036 306326 330340 306354
rect 330404 310406 330602 310434
rect 329944 271250 329972 306274
rect 330036 280906 330064 306326
rect 330404 302234 330432 310406
rect 330772 305833 330800 310420
rect 330956 306338 330984 310420
rect 331140 306406 331168 310420
rect 331324 306474 331352 310420
rect 331312 306468 331364 306474
rect 331312 306410 331364 306416
rect 331128 306400 331180 306406
rect 331128 306342 331180 306348
rect 331220 306400 331272 306406
rect 331220 306342 331272 306348
rect 330944 306332 330996 306338
rect 330944 306274 330996 306280
rect 330758 305824 330814 305833
rect 330758 305759 330814 305768
rect 330128 302206 330432 302234
rect 330128 291922 330156 302206
rect 330116 291916 330168 291922
rect 330116 291858 330168 291864
rect 330024 280900 330076 280906
rect 330024 280842 330076 280848
rect 329932 271244 329984 271250
rect 329932 271186 329984 271192
rect 329840 261588 329892 261594
rect 329840 261530 329892 261536
rect 328552 254720 328604 254726
rect 328552 254662 328604 254668
rect 331232 250578 331260 306342
rect 331312 306332 331364 306338
rect 331508 306320 331536 310420
rect 331312 306274 331364 306280
rect 331416 306292 331536 306320
rect 331324 265810 331352 306274
rect 331416 269958 331444 306292
rect 331692 306252 331720 310420
rect 331772 306468 331824 306474
rect 331772 306410 331824 306416
rect 331508 306224 331720 306252
rect 331508 289202 331536 306224
rect 331784 304366 331812 306410
rect 331772 304360 331824 304366
rect 331772 304302 331824 304308
rect 331876 303113 331904 310420
rect 332060 306338 332088 310420
rect 332244 306406 332272 310420
rect 332232 306400 332284 306406
rect 332232 306342 332284 306348
rect 332048 306332 332100 306338
rect 332048 306274 332100 306280
rect 331862 303104 331918 303113
rect 331862 303039 331918 303048
rect 332428 302234 332456 310420
rect 332612 306406 332640 310420
rect 332796 309134 332824 310420
rect 332994 310406 333192 310434
rect 332704 309106 332824 309134
rect 332600 306400 332652 306406
rect 332600 306342 332652 306348
rect 332600 306264 332652 306270
rect 332600 306206 332652 306212
rect 331600 302206 332456 302234
rect 331600 301578 331628 302206
rect 331588 301572 331640 301578
rect 331588 301514 331640 301520
rect 331496 289196 331548 289202
rect 331496 289138 331548 289144
rect 331404 269952 331456 269958
rect 331404 269894 331456 269900
rect 331312 265804 331364 265810
rect 331312 265746 331364 265752
rect 331220 250572 331272 250578
rect 331220 250514 331272 250520
rect 328460 249144 328512 249150
rect 328460 249086 328512 249092
rect 325700 247920 325752 247926
rect 325700 247862 325752 247868
rect 332612 247858 332640 306206
rect 332704 253434 332732 309106
rect 332876 306400 332928 306406
rect 332876 306342 332928 306348
rect 333060 306400 333112 306406
rect 333060 306342 333112 306348
rect 332784 306196 332836 306202
rect 332784 306138 332836 306144
rect 332692 253428 332744 253434
rect 332692 253370 332744 253376
rect 332796 253366 332824 306138
rect 332888 267170 332916 306342
rect 332968 306332 333020 306338
rect 332968 306274 333020 306280
rect 332980 279546 333008 306274
rect 333072 298858 333100 306342
rect 333164 300286 333192 310406
rect 333256 306338 333284 310420
rect 333244 306332 333296 306338
rect 333244 306274 333296 306280
rect 333440 306202 333468 310420
rect 333624 306406 333652 310420
rect 333612 306400 333664 306406
rect 333612 306342 333664 306348
rect 333808 306270 333836 310420
rect 333992 306320 334020 310420
rect 334176 306320 334204 310420
rect 334360 306388 334388 310420
rect 334360 306360 334480 306388
rect 333992 306292 334112 306320
rect 334176 306292 334388 306320
rect 333796 306264 333848 306270
rect 333796 306206 333848 306212
rect 333428 306196 333480 306202
rect 333428 306138 333480 306144
rect 333980 306196 334032 306202
rect 333980 306138 334032 306144
rect 333152 300280 333204 300286
rect 333152 300222 333204 300228
rect 333060 298852 333112 298858
rect 333060 298794 333112 298800
rect 332968 279540 333020 279546
rect 332968 279482 333020 279488
rect 332876 267164 332928 267170
rect 332876 267106 332928 267112
rect 332784 253360 332836 253366
rect 332784 253302 332836 253308
rect 332600 247852 332652 247858
rect 332600 247794 332652 247800
rect 324320 245200 324372 245206
rect 324320 245142 324372 245148
rect 333992 245070 334020 306138
rect 334084 245138 334112 306292
rect 334164 306128 334216 306134
rect 334164 306070 334216 306076
rect 334176 246430 334204 306070
rect 334256 302524 334308 302530
rect 334256 302466 334308 302472
rect 334268 246498 334296 302466
rect 334360 246566 334388 306292
rect 334452 306202 334480 306360
rect 334544 306320 334572 310420
rect 334544 306292 334664 306320
rect 334440 306196 334492 306202
rect 334440 306138 334492 306144
rect 334532 306196 334584 306202
rect 334532 306138 334584 306144
rect 334440 306060 334492 306066
rect 334440 306002 334492 306008
rect 334452 247790 334480 306002
rect 334544 251870 334572 306138
rect 334636 253298 334664 306292
rect 334728 302530 334756 310420
rect 334912 306202 334940 310420
rect 334900 306196 334952 306202
rect 334900 306138 334952 306144
rect 335096 306134 335124 310420
rect 335084 306128 335136 306134
rect 335084 306070 335136 306076
rect 335280 306066 335308 310420
rect 335478 310406 335676 310434
rect 335360 306400 335412 306406
rect 335360 306342 335412 306348
rect 335268 306060 335320 306066
rect 335268 306002 335320 306008
rect 334716 302524 334768 302530
rect 334716 302466 334768 302472
rect 334624 253292 334676 253298
rect 334624 253234 334676 253240
rect 334532 251864 334584 251870
rect 334532 251806 334584 251812
rect 334440 247784 334492 247790
rect 334440 247726 334492 247732
rect 334348 246560 334400 246566
rect 334348 246502 334400 246508
rect 334256 246492 334308 246498
rect 334256 246434 334308 246440
rect 334164 246424 334216 246430
rect 334164 246366 334216 246372
rect 335372 246362 335400 306342
rect 335544 306332 335596 306338
rect 335544 306274 335596 306280
rect 335452 306264 335504 306270
rect 335452 306206 335504 306212
rect 335464 249082 335492 306206
rect 335556 269890 335584 306274
rect 335648 278118 335676 310406
rect 335740 293350 335768 310420
rect 335924 304298 335952 310420
rect 336108 306406 336136 310420
rect 336096 306400 336148 306406
rect 336096 306342 336148 306348
rect 336292 306338 336320 310420
rect 336280 306332 336332 306338
rect 336280 306274 336332 306280
rect 335912 304292 335964 304298
rect 335912 304234 335964 304240
rect 336476 302234 336504 310420
rect 336660 306270 336688 310420
rect 336844 306474 336872 310420
rect 337028 307902 337056 310420
rect 337212 309134 337240 310420
rect 337120 309106 337240 309134
rect 337016 307896 337068 307902
rect 337016 307838 337068 307844
rect 336832 306468 336884 306474
rect 336832 306410 336884 306416
rect 336740 306400 336792 306406
rect 336740 306342 336792 306348
rect 336648 306264 336700 306270
rect 336648 306206 336700 306212
rect 335832 302206 336504 302234
rect 335832 296070 335860 302206
rect 335820 296064 335872 296070
rect 335820 296006 335872 296012
rect 335728 293344 335780 293350
rect 335728 293286 335780 293292
rect 335636 278112 335688 278118
rect 335636 278054 335688 278060
rect 335544 269884 335596 269890
rect 335544 269826 335596 269832
rect 335452 249076 335504 249082
rect 335452 249018 335504 249024
rect 336752 247722 336780 306342
rect 336924 306332 336976 306338
rect 337120 306320 337148 309106
rect 337292 307896 337344 307902
rect 337292 307838 337344 307844
rect 337200 306468 337252 306474
rect 337200 306410 337252 306416
rect 336924 306274 336976 306280
rect 337028 306292 337148 306320
rect 336832 306264 336884 306270
rect 336832 306206 336884 306212
rect 336844 253230 336872 306206
rect 336936 275330 336964 306274
rect 337028 276758 337056 306292
rect 337212 306252 337240 306410
rect 337120 306224 337240 306252
rect 337120 283694 337148 306224
rect 337304 302977 337332 307838
rect 337396 306406 337424 310420
rect 337384 306400 337436 306406
rect 337384 306342 337436 306348
rect 337290 302968 337346 302977
rect 337290 302903 337346 302912
rect 337580 302234 337608 310420
rect 337764 306338 337792 310420
rect 337752 306332 337804 306338
rect 337752 306274 337804 306280
rect 337948 306270 337976 310420
rect 338146 310406 338252 310434
rect 338120 306332 338172 306338
rect 338120 306274 338172 306280
rect 337936 306264 337988 306270
rect 337936 306206 337988 306212
rect 337212 302206 337608 302234
rect 337212 294642 337240 302206
rect 337200 294636 337252 294642
rect 337200 294578 337252 294584
rect 337108 283688 337160 283694
rect 337108 283630 337160 283636
rect 337016 276752 337068 276758
rect 337016 276694 337068 276700
rect 336924 275324 336976 275330
rect 336924 275266 336976 275272
rect 336832 253224 336884 253230
rect 336832 253166 336884 253172
rect 336740 247716 336792 247722
rect 336740 247658 336792 247664
rect 335360 246356 335412 246362
rect 335360 246298 335412 246304
rect 334072 245132 334124 245138
rect 334072 245074 334124 245080
rect 333980 245064 334032 245070
rect 333980 245006 334032 245012
rect 338132 245002 338160 306274
rect 338224 306202 338252 310406
rect 338316 310406 338422 310434
rect 338212 306196 338264 306202
rect 338212 306138 338264 306144
rect 338212 306060 338264 306066
rect 338212 306002 338264 306008
rect 338224 265742 338252 306002
rect 338316 274038 338344 310406
rect 338592 306388 338620 310420
rect 338408 306360 338620 306388
rect 338408 279478 338436 306360
rect 338776 306320 338804 310420
rect 338856 308984 338908 308990
rect 338856 308926 338908 308932
rect 338592 306292 338804 306320
rect 338488 306264 338540 306270
rect 338488 306206 338540 306212
rect 338500 291854 338528 306206
rect 338592 293282 338620 306292
rect 338672 306196 338724 306202
rect 338672 306138 338724 306144
rect 338684 301510 338712 306138
rect 338672 301504 338724 301510
rect 338672 301446 338724 301452
rect 338868 296714 338896 308926
rect 338960 306338 338988 310420
rect 338948 306332 339000 306338
rect 338948 306274 339000 306280
rect 339144 306066 339172 310420
rect 339328 306270 339356 310420
rect 339512 306354 339540 310420
rect 339696 306474 339724 310420
rect 339684 306468 339736 306474
rect 339684 306410 339736 306416
rect 339512 306326 339816 306354
rect 339316 306264 339368 306270
rect 339316 306206 339368 306212
rect 339684 306264 339736 306270
rect 339684 306206 339736 306212
rect 339500 306196 339552 306202
rect 339500 306138 339552 306144
rect 339132 306060 339184 306066
rect 339132 306002 339184 306008
rect 338776 296686 338896 296714
rect 338580 293276 338632 293282
rect 338580 293218 338632 293224
rect 338488 291848 338540 291854
rect 338488 291790 338540 291796
rect 338396 279472 338448 279478
rect 338396 279414 338448 279420
rect 338304 274032 338356 274038
rect 338304 273974 338356 273980
rect 338212 265736 338264 265742
rect 338212 265678 338264 265684
rect 338776 249286 338804 296686
rect 339512 260234 339540 306138
rect 339592 306128 339644 306134
rect 339592 306070 339644 306076
rect 339604 271182 339632 306070
rect 339696 272542 339724 306206
rect 339788 283626 339816 306326
rect 339880 300218 339908 310420
rect 339960 306468 340012 306474
rect 339960 306410 340012 306416
rect 339972 302841 340000 306410
rect 340064 306270 340092 310420
rect 340052 306264 340104 306270
rect 340052 306206 340104 306212
rect 340248 306202 340276 310420
rect 340432 307086 340460 310420
rect 340420 307080 340472 307086
rect 340420 307022 340472 307028
rect 340236 306196 340288 306202
rect 340236 306138 340288 306144
rect 340616 306134 340644 310420
rect 340892 306626 340920 310420
rect 340892 306598 341012 306626
rect 340880 306468 340932 306474
rect 340880 306410 340932 306416
rect 340604 306128 340656 306134
rect 340604 306070 340656 306076
rect 339958 302832 340014 302841
rect 339958 302767 340014 302776
rect 339868 300212 339920 300218
rect 339868 300154 339920 300160
rect 339776 283620 339828 283626
rect 339776 283562 339828 283568
rect 339684 272536 339736 272542
rect 339684 272478 339736 272484
rect 339592 271176 339644 271182
rect 339592 271118 339644 271124
rect 340892 264246 340920 306410
rect 340984 306202 341012 306598
rect 341076 306270 341104 310420
rect 341064 306264 341116 306270
rect 341064 306206 341116 306212
rect 340972 306196 341024 306202
rect 340972 306138 341024 306144
rect 341064 306128 341116 306134
rect 341064 306070 341116 306076
rect 340972 306060 341024 306066
rect 340972 306002 341024 306008
rect 340984 267102 341012 306002
rect 341076 269822 341104 306070
rect 341156 302796 341208 302802
rect 341156 302738 341208 302744
rect 341168 289134 341196 302738
rect 341260 290562 341288 310420
rect 341444 306474 341472 310420
rect 341432 306468 341484 306474
rect 341432 306410 341484 306416
rect 341628 306354 341656 310420
rect 341352 306326 341656 306354
rect 341248 290556 341300 290562
rect 341248 290498 341300 290504
rect 341352 290494 341380 306326
rect 341432 306264 341484 306270
rect 341432 306206 341484 306212
rect 341444 298790 341472 306206
rect 341524 306196 341576 306202
rect 341524 306138 341576 306144
rect 341536 300150 341564 306138
rect 341812 306134 341840 310420
rect 341800 306128 341852 306134
rect 341800 306070 341852 306076
rect 341996 306066 342024 310420
rect 341984 306060 342036 306066
rect 341984 306002 342036 306008
rect 342180 302802 342208 310420
rect 342260 306332 342312 306338
rect 342260 306274 342312 306280
rect 342168 302796 342220 302802
rect 342168 302738 342220 302744
rect 341524 300144 341576 300150
rect 341524 300086 341576 300092
rect 341432 298784 341484 298790
rect 341432 298726 341484 298732
rect 341340 290488 341392 290494
rect 341340 290430 341392 290436
rect 341156 289128 341208 289134
rect 341156 289070 341208 289076
rect 341064 269816 341116 269822
rect 341064 269758 341116 269764
rect 340972 267096 341024 267102
rect 340972 267038 341024 267044
rect 340880 264240 340932 264246
rect 340880 264182 340932 264188
rect 339500 260228 339552 260234
rect 339500 260170 339552 260176
rect 342272 260166 342300 306274
rect 342364 306218 342392 310420
rect 342548 306354 342576 310420
rect 342732 306354 342760 310420
rect 342548 306326 342668 306354
rect 342732 306326 342852 306354
rect 342916 306338 342944 310420
rect 342364 306190 342576 306218
rect 342444 306128 342496 306134
rect 342444 306070 342496 306076
rect 342352 306060 342404 306066
rect 342352 306002 342404 306008
rect 342364 265674 342392 306002
rect 342456 276690 342484 306070
rect 342548 282198 342576 306190
rect 342640 287774 342668 306326
rect 342720 306264 342772 306270
rect 342720 306206 342772 306212
rect 342628 287768 342680 287774
rect 342628 287710 342680 287716
rect 342732 287706 342760 306206
rect 342824 297430 342852 306326
rect 342904 306332 342956 306338
rect 342904 306274 342956 306280
rect 343100 306134 343128 310420
rect 343284 306270 343312 310420
rect 343376 310406 343574 310434
rect 343272 306264 343324 306270
rect 343272 306206 343324 306212
rect 343088 306128 343140 306134
rect 343088 306070 343140 306076
rect 343376 306066 343404 310406
rect 343364 306060 343416 306066
rect 343364 306002 343416 306008
rect 343640 305244 343692 305250
rect 343640 305186 343692 305192
rect 342812 297424 342864 297430
rect 342812 297366 342864 297372
rect 342720 287700 342772 287706
rect 342720 287642 342772 287648
rect 342536 282192 342588 282198
rect 342536 282134 342588 282140
rect 342444 276684 342496 276690
rect 342444 276626 342496 276632
rect 342352 265668 342404 265674
rect 342352 265610 342404 265616
rect 342260 260160 342312 260166
rect 342260 260102 342312 260108
rect 338764 249280 338816 249286
rect 338764 249222 338816 249228
rect 338120 244996 338172 245002
rect 338120 244938 338172 244944
rect 343652 244934 343680 305186
rect 343744 254658 343772 310420
rect 343824 306332 343876 306338
rect 343824 306274 343876 306280
rect 343732 254652 343784 254658
rect 343732 254594 343784 254600
rect 343836 254590 343864 306274
rect 343928 305998 343956 310420
rect 344112 306354 344140 310420
rect 344020 306326 344140 306354
rect 344296 306338 344324 310420
rect 344284 306332 344336 306338
rect 343916 305992 343968 305998
rect 343916 305934 343968 305940
rect 343916 305856 343968 305862
rect 343916 305798 343968 305804
rect 343928 261526 343956 305798
rect 344020 267034 344048 306326
rect 344284 306274 344336 306280
rect 344480 306082 344508 310420
rect 344112 306054 344508 306082
rect 344112 286346 344140 306054
rect 344192 305992 344244 305998
rect 344192 305934 344244 305940
rect 344204 296002 344232 305934
rect 344664 305862 344692 310420
rect 344652 305856 344704 305862
rect 344652 305798 344704 305804
rect 344848 305250 344876 310420
rect 345032 306474 345060 310420
rect 345020 306468 345072 306474
rect 345020 306410 345072 306416
rect 345112 306400 345164 306406
rect 345112 306342 345164 306348
rect 345020 306332 345072 306338
rect 345020 306274 345072 306280
rect 344836 305244 344888 305250
rect 344836 305186 344888 305192
rect 344192 295996 344244 296002
rect 344192 295938 344244 295944
rect 344100 286340 344152 286346
rect 344100 286282 344152 286288
rect 344008 267028 344060 267034
rect 344008 266970 344060 266976
rect 343916 261520 343968 261526
rect 343916 261462 343968 261468
rect 343824 254584 343876 254590
rect 343824 254526 343876 254532
rect 345032 250510 345060 306274
rect 345124 261662 345152 306342
rect 345216 306082 345244 310420
rect 345400 306490 345428 310420
rect 345308 306462 345428 306490
rect 345480 306468 345532 306474
rect 345308 306270 345336 306462
rect 345480 306410 345532 306416
rect 345296 306264 345348 306270
rect 345296 306206 345348 306212
rect 345216 306054 345428 306082
rect 345204 305992 345256 305998
rect 345204 305934 345256 305940
rect 345296 305992 345348 305998
rect 345296 305934 345348 305940
rect 345216 262886 345244 305934
rect 345308 278050 345336 305934
rect 345400 280838 345428 306054
rect 345492 305697 345520 306410
rect 345478 305688 345534 305697
rect 345478 305623 345534 305632
rect 345584 302234 345612 310420
rect 345768 306338 345796 310420
rect 345860 310406 346058 310434
rect 345756 306332 345808 306338
rect 345756 306274 345808 306280
rect 345860 305998 345888 310406
rect 346228 306406 346256 310420
rect 346216 306400 346268 306406
rect 346216 306342 346268 306348
rect 345848 305992 345900 305998
rect 345848 305934 345900 305940
rect 345492 302206 345612 302234
rect 345492 284986 345520 302206
rect 345480 284980 345532 284986
rect 345480 284922 345532 284928
rect 345388 280832 345440 280838
rect 345388 280774 345440 280780
rect 345296 278044 345348 278050
rect 345296 277986 345348 277992
rect 345204 262880 345256 262886
rect 345204 262822 345256 262828
rect 345112 261656 345164 261662
rect 345112 261598 345164 261604
rect 345020 250504 345072 250510
rect 345020 250446 345072 250452
rect 346412 246770 346440 310420
rect 346596 306354 346624 310420
rect 346780 309097 346808 310420
rect 346766 309088 346822 309097
rect 346766 309023 346822 309032
rect 346964 308961 346992 310420
rect 346950 308952 347006 308961
rect 346950 308887 347006 308896
rect 346504 306326 346624 306354
rect 346504 258738 346532 306326
rect 347148 305658 347176 310420
rect 347136 305652 347188 305658
rect 347136 305594 347188 305600
rect 347332 302234 347360 310420
rect 347516 308825 347544 310420
rect 347700 309126 347728 310420
rect 347688 309120 347740 309126
rect 347688 309062 347740 309068
rect 347502 308816 347558 308825
rect 347502 308751 347558 308760
rect 347884 306490 347912 310420
rect 347884 306462 348004 306490
rect 347780 306400 347832 306406
rect 347780 306342 347832 306348
rect 346596 302206 347360 302234
rect 346596 297566 346624 302206
rect 346584 297560 346636 297566
rect 346584 297502 346636 297508
rect 346492 258732 346544 258738
rect 346492 258674 346544 258680
rect 347792 252074 347820 306342
rect 347872 306332 347924 306338
rect 347872 306274 347924 306280
rect 347884 267238 347912 306274
rect 347976 303550 348004 306462
rect 347964 303544 348016 303550
rect 347964 303486 348016 303492
rect 348068 302234 348096 310420
rect 348252 306338 348280 310420
rect 348436 308689 348464 310420
rect 348712 309058 348740 310420
rect 348700 309052 348752 309058
rect 348700 308994 348752 309000
rect 348516 308984 348568 308990
rect 348516 308926 348568 308932
rect 348422 308680 348478 308689
rect 348422 308615 348478 308624
rect 348424 307828 348476 307834
rect 348424 307770 348476 307776
rect 348240 306332 348292 306338
rect 348240 306274 348292 306280
rect 347976 302206 348096 302234
rect 347976 301646 348004 302206
rect 347964 301640 348016 301646
rect 347964 301582 348016 301588
rect 347872 267232 347924 267238
rect 347872 267174 347924 267180
rect 348436 253502 348464 307770
rect 348528 290698 348556 308926
rect 348896 303210 348924 310420
rect 349080 306406 349108 310420
rect 349068 306400 349120 306406
rect 349264 306377 349292 310420
rect 349068 306342 349120 306348
rect 349250 306368 349306 306377
rect 349250 306303 349306 306312
rect 349448 305454 349476 310420
rect 349436 305448 349488 305454
rect 349436 305390 349488 305396
rect 348884 303204 348936 303210
rect 348884 303146 348936 303152
rect 349632 303142 349660 310420
rect 349620 303136 349672 303142
rect 349620 303078 349672 303084
rect 349816 302234 349844 310420
rect 350000 306241 350028 310420
rect 349986 306232 350042 306241
rect 349986 306167 350042 306176
rect 350184 303414 350212 310420
rect 350368 307834 350396 310420
rect 350356 307828 350408 307834
rect 350356 307770 350408 307776
rect 350552 306490 350580 310420
rect 350552 306462 350672 306490
rect 350540 306332 350592 306338
rect 350540 306274 350592 306280
rect 350172 303408 350224 303414
rect 350172 303350 350224 303356
rect 349724 302206 349844 302234
rect 349724 293486 349752 302206
rect 349712 293480 349764 293486
rect 349712 293422 349764 293428
rect 348516 290692 348568 290698
rect 348516 290634 348568 290640
rect 350552 256290 350580 306274
rect 350644 305561 350672 306462
rect 350630 305552 350686 305561
rect 350630 305487 350686 305496
rect 350736 302870 350764 310420
rect 350724 302864 350776 302870
rect 350724 302806 350776 302812
rect 350920 302234 350948 310420
rect 351196 305726 351224 310420
rect 351184 305720 351236 305726
rect 351184 305662 351236 305668
rect 351380 302734 351408 310420
rect 351564 306338 351592 310420
rect 351552 306332 351604 306338
rect 351552 306274 351604 306280
rect 351748 305250 351776 310420
rect 351736 305244 351788 305250
rect 351736 305186 351788 305192
rect 351932 303278 351960 310420
rect 352116 308990 352144 310420
rect 352104 308984 352156 308990
rect 352104 308926 352156 308932
rect 352300 305590 352328 310420
rect 352288 305584 352340 305590
rect 352288 305526 352340 305532
rect 352484 303482 352512 310420
rect 352668 305318 352696 310420
rect 352656 305312 352708 305318
rect 352656 305254 352708 305260
rect 352472 303476 352524 303482
rect 352472 303418 352524 303424
rect 352852 303346 352880 310420
rect 353036 307834 353064 310420
rect 353024 307828 353076 307834
rect 353024 307770 353076 307776
rect 353220 306338 353248 310420
rect 353404 307902 353432 310420
rect 353392 307896 353444 307902
rect 353392 307838 353444 307844
rect 353208 306332 353260 306338
rect 353208 306274 353260 306280
rect 353588 305862 353616 310420
rect 353864 308310 353892 310420
rect 353852 308304 353904 308310
rect 353852 308246 353904 308252
rect 354048 306066 354076 310420
rect 354232 309194 354260 310420
rect 354220 309188 354272 309194
rect 354220 309130 354272 309136
rect 354036 306060 354088 306066
rect 354036 306002 354088 306008
rect 353576 305856 353628 305862
rect 353576 305798 353628 305804
rect 354416 305794 354444 310420
rect 354600 308174 354628 310420
rect 354588 308168 354640 308174
rect 354588 308110 354640 308116
rect 354784 305998 354812 310420
rect 354968 308242 354996 310420
rect 354956 308236 355008 308242
rect 354956 308178 355008 308184
rect 354772 305992 354824 305998
rect 354772 305934 354824 305940
rect 355152 305930 355180 310420
rect 355232 308780 355284 308786
rect 355232 308722 355284 308728
rect 355140 305924 355192 305930
rect 355140 305866 355192 305872
rect 354404 305788 354456 305794
rect 354404 305730 354456 305736
rect 352840 303340 352892 303346
rect 352840 303282 352892 303288
rect 351920 303272 351972 303278
rect 351920 303214 351972 303220
rect 351368 302728 351420 302734
rect 351368 302670 351420 302676
rect 350644 302206 350948 302234
rect 355244 302234 355272 308722
rect 355336 308378 355364 310420
rect 355520 308802 355548 310420
rect 355704 309126 355732 310420
rect 355692 309120 355744 309126
rect 355692 309062 355744 309068
rect 355520 308774 355824 308802
rect 355508 308712 355560 308718
rect 355508 308654 355560 308660
rect 355416 308508 355468 308514
rect 355416 308450 355468 308456
rect 355324 308372 355376 308378
rect 355324 308314 355376 308320
rect 355244 302206 355364 302234
rect 350644 283830 350672 302206
rect 350632 283824 350684 283830
rect 350632 283766 350684 283772
rect 350540 256284 350592 256290
rect 350540 256226 350592 256232
rect 348424 253496 348476 253502
rect 348424 253438 348476 253444
rect 347780 252068 347832 252074
rect 347780 252010 347832 252016
rect 346400 246764 346452 246770
rect 346400 246706 346452 246712
rect 343640 244928 343692 244934
rect 343640 244870 343692 244876
rect 310518 244760 310574 244769
rect 310518 244695 310574 244704
rect 355336 244526 355364 302206
rect 355324 244520 355376 244526
rect 355324 244462 355376 244468
rect 355428 244322 355456 308450
rect 355520 245546 355548 308654
rect 355692 308644 355744 308650
rect 355692 308586 355744 308592
rect 355600 308576 355652 308582
rect 355600 308518 355652 308524
rect 355612 245614 355640 308518
rect 355704 247586 355732 308586
rect 355796 305522 355824 308774
rect 355784 305516 355836 305522
rect 355784 305458 355836 305464
rect 355888 303618 355916 310420
rect 356072 308650 356100 310420
rect 356060 308644 356112 308650
rect 356060 308586 356112 308592
rect 356348 306202 356376 310420
rect 356532 308854 356560 310420
rect 356520 308848 356572 308854
rect 356520 308790 356572 308796
rect 356520 308440 356572 308446
rect 356520 308382 356572 308388
rect 356532 306270 356560 308382
rect 356716 306626 356744 310420
rect 356900 308446 356928 310420
rect 356888 308440 356940 308446
rect 356888 308382 356940 308388
rect 356624 306598 356744 306626
rect 356520 306264 356572 306270
rect 356520 306206 356572 306212
rect 356336 306196 356388 306202
rect 356336 306138 356388 306144
rect 355876 303612 355928 303618
rect 355876 303554 355928 303560
rect 356624 302802 356652 306598
rect 357084 306490 357112 310420
rect 357164 308780 357216 308786
rect 357164 308722 357216 308728
rect 356716 306462 357112 306490
rect 356612 302796 356664 302802
rect 356612 302738 356664 302744
rect 355692 247580 355744 247586
rect 355692 247522 355744 247528
rect 355600 245608 355652 245614
rect 355600 245550 355652 245556
rect 355508 245540 355560 245546
rect 355508 245482 355560 245488
rect 355416 244316 355468 244322
rect 355416 244258 355468 244264
rect 303620 243908 303672 243914
rect 303620 243850 303672 243856
rect 299756 243772 299808 243778
rect 299756 243714 299808 243720
rect 299572 243568 299624 243574
rect 297272 243510 297324 243516
rect 298098 243536 298154 243545
rect 299572 243510 299624 243516
rect 298098 243471 298154 243480
rect 278134 159896 278190 159905
rect 278134 159831 278190 159840
rect 271050 159624 271106 159633
rect 271050 159559 271106 159568
rect 275834 159624 275890 159633
rect 275834 159559 275890 159568
rect 256700 159520 256752 159526
rect 256700 159462 256752 159468
rect 239588 158772 239640 158778
rect 239588 158714 239640 158720
rect 238116 158704 238168 158710
rect 220818 158672 220874 158681
rect 238114 158672 238116 158681
rect 239600 158681 239628 158714
rect 238168 158672 238170 158681
rect 220818 158607 220874 158616
rect 230480 158636 230532 158642
rect 219438 157856 219494 157865
rect 219438 157791 219494 157800
rect 219452 16574 219480 157791
rect 220832 16574 220860 158607
rect 238114 158607 238170 158616
rect 239586 158672 239642 158681
rect 239586 158607 239642 158616
rect 240690 158672 240746 158681
rect 240690 158607 240746 158616
rect 248326 158672 248382 158681
rect 248326 158607 248382 158616
rect 250442 158672 250498 158681
rect 250442 158607 250498 158616
rect 252374 158672 252430 158681
rect 252374 158607 252430 158616
rect 254950 158672 255006 158681
rect 254950 158607 255006 158616
rect 255870 158672 255926 158681
rect 255870 158607 255926 158616
rect 230480 158578 230532 158584
rect 224958 158536 225014 158545
rect 224958 158471 225014 158480
rect 223578 158400 223634 158409
rect 223578 158335 223634 158344
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219348 3528 219400 3534
rect 219254 3496 219310 3505
rect 219348 3470 219400 3476
rect 219254 3431 219310 3440
rect 219268 480 219296 3431
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222752 3324 222804 3330
rect 222752 3266 222804 3272
rect 222764 480 222792 3266
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 158335
rect 224972 16574 225000 158471
rect 227718 158264 227774 158273
rect 227718 158199 227774 158208
rect 227732 16574 227760 158199
rect 229100 157820 229152 157826
rect 229100 157762 229152 157768
rect 229112 16574 229140 157762
rect 230492 16574 230520 158578
rect 236000 158568 236052 158574
rect 236000 158510 236052 158516
rect 234712 158500 234764 158506
rect 234712 158442 234764 158448
rect 231858 158128 231914 158137
rect 231858 158063 231914 158072
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 225156 480 225184 16546
rect 227536 3392 227588 3398
rect 227536 3334 227588 3340
rect 226340 3256 226392 3262
rect 226340 3198 226392 3204
rect 226352 480 226380 3198
rect 227548 480 227576 3334
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 158063
rect 233240 157956 233292 157962
rect 233240 157898 233292 157904
rect 233252 16574 233280 157898
rect 234620 157888 234672 157894
rect 234620 157830 234672 157836
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11762 234660 157830
rect 234620 11756 234672 11762
rect 234620 11698 234672 11704
rect 234724 6914 234752 158442
rect 236012 16574 236040 158510
rect 238758 157992 238814 158001
rect 238758 157927 238814 157936
rect 237380 155848 237432 155854
rect 237380 155790 237432 155796
rect 237392 16574 237420 155790
rect 238772 16574 238800 157927
rect 240704 157758 240732 158607
rect 242992 158432 243044 158438
rect 242992 158374 243044 158380
rect 242900 158364 242952 158370
rect 242900 158306 242952 158312
rect 240692 157752 240744 157758
rect 240692 157694 240744 157700
rect 241520 155780 241572 155786
rect 241520 155722 241572 155728
rect 241532 16574 241560 155722
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 235816 11756 235868 11762
rect 235816 11698 235868 11704
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11698
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240508 4140 240560 4146
rect 240508 4082 240560 4088
rect 240520 480 240548 4082
rect 241716 480 241744 16546
rect 242912 11762 242940 158306
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 243004 6914 243032 158374
rect 245660 158296 245712 158302
rect 245660 158238 245712 158244
rect 245672 16574 245700 158238
rect 247040 158228 247092 158234
rect 247040 158170 247092 158176
rect 246854 158128 246910 158137
rect 246854 158063 246910 158072
rect 246868 155961 246896 158063
rect 246854 155952 246910 155961
rect 246854 155887 246910 155896
rect 247052 16574 247080 158170
rect 248340 157350 248368 158607
rect 249800 158024 249852 158030
rect 248694 157992 248750 158001
rect 249800 157966 249852 157972
rect 248694 157927 248750 157936
rect 248328 157344 248380 157350
rect 248328 157286 248380 157292
rect 248708 155922 248736 157927
rect 248696 155916 248748 155922
rect 248696 155858 248748 155864
rect 248420 155712 248472 155718
rect 248420 155654 248472 155660
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11698
rect 245200 4072 245252 4078
rect 245200 4014 245252 4020
rect 245212 480 245240 4014
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 155654
rect 249812 16574 249840 157966
rect 250456 157214 250484 158607
rect 251180 158160 251232 158166
rect 251180 158102 251232 158108
rect 250444 157208 250496 157214
rect 250444 157150 250496 157156
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 158102
rect 252282 157992 252338 158001
rect 252282 157927 252338 157936
rect 252296 155854 252324 157927
rect 252388 157282 252416 158607
rect 252560 158092 252612 158098
rect 252560 158034 252612 158040
rect 252376 157276 252428 157282
rect 252376 157218 252428 157224
rect 252284 155848 252336 155854
rect 252284 155790 252336 155796
rect 251270 155544 251326 155553
rect 251270 155479 251326 155488
rect 251284 16574 251312 155479
rect 252572 16574 252600 158034
rect 253570 157992 253626 158001
rect 253570 157927 253626 157936
rect 253584 155786 253612 157927
rect 253662 157448 253718 157457
rect 253662 157383 253718 157392
rect 253572 155780 253624 155786
rect 253572 155722 253624 155728
rect 253676 154562 253704 157383
rect 254964 157146 254992 158607
rect 254952 157140 255004 157146
rect 254952 157082 255004 157088
rect 255884 156942 255912 158607
rect 256238 157448 256294 157457
rect 256238 157383 256294 157392
rect 255872 156936 255924 156942
rect 255872 156878 255924 156884
rect 253940 155644 253992 155650
rect 253940 155586 253992 155592
rect 253664 154556 253716 154562
rect 253664 154498 253716 154504
rect 253952 16574 253980 155586
rect 255320 155508 255372 155514
rect 255320 155450 255372 155456
rect 255332 16574 255360 155450
rect 256252 154494 256280 157383
rect 256240 154488 256292 154494
rect 256240 154430 256292 154436
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 159462
rect 259460 159452 259512 159458
rect 259460 159394 259512 159400
rect 257250 158672 257306 158681
rect 257250 158607 257306 158616
rect 259090 158672 259146 158681
rect 259090 158607 259146 158616
rect 257264 157078 257292 158607
rect 257252 157072 257304 157078
rect 257252 157014 257304 157020
rect 259104 157010 259132 158607
rect 259092 157004 259144 157010
rect 259092 156946 259144 156952
rect 259472 151814 259500 159394
rect 263692 159384 263744 159390
rect 263692 159326 263744 159332
rect 259550 158672 259606 158681
rect 259550 158607 259606 158616
rect 261482 158672 261538 158681
rect 261482 158607 261538 158616
rect 262862 158672 262918 158681
rect 262862 158607 262918 158616
rect 263598 158672 263654 158681
rect 263598 158607 263654 158616
rect 259564 158506 259592 158607
rect 259552 158500 259604 158506
rect 259552 158442 259604 158448
rect 260654 157992 260710 158001
rect 260654 157927 260710 157936
rect 260668 155718 260696 157927
rect 261496 157690 261524 158607
rect 262876 158574 262904 158607
rect 262864 158568 262916 158574
rect 262864 158510 262916 158516
rect 263612 158438 263640 158607
rect 263600 158432 263652 158438
rect 263600 158374 263652 158380
rect 261758 157856 261814 157865
rect 261758 157791 261814 157800
rect 261484 157684 261536 157690
rect 261484 157626 261536 157632
rect 260656 155712 260708 155718
rect 260656 155654 260708 155660
rect 261772 155650 261800 157791
rect 261760 155644 261812 155650
rect 261760 155586 261812 155592
rect 260840 155372 260892 155378
rect 260840 155314 260892 155320
rect 259472 151786 259592 151814
rect 259564 6914 259592 151786
rect 260852 16574 260880 155314
rect 263704 142154 263732 159326
rect 268750 158672 268806 158681
rect 268750 158607 268806 158616
rect 269854 158672 269910 158681
rect 269854 158607 269910 158616
rect 268764 158370 268792 158607
rect 268752 158364 268804 158370
rect 268752 158306 268804 158312
rect 269868 158302 269896 158607
rect 269856 158296 269908 158302
rect 267646 158264 267702 158273
rect 269856 158238 269908 158244
rect 267646 158199 267702 158208
rect 264518 157856 264574 157865
rect 264518 157791 264574 157800
rect 266910 157856 266966 157865
rect 266910 157791 266966 157800
rect 264532 155514 264560 157791
rect 265990 157720 266046 157729
rect 265990 157655 266046 157664
rect 264520 155508 264572 155514
rect 264520 155450 264572 155456
rect 264980 155440 265032 155446
rect 264980 155382 265032 155388
rect 263612 142126 263732 142154
rect 263612 16574 263640 142126
rect 260852 16546 261800 16574
rect 263612 16546 264192 16574
rect 259472 6886 259592 6914
rect 258264 4004 258316 4010
rect 258264 3946 258316 3952
rect 258276 480 258304 3946
rect 259472 480 259500 6886
rect 260656 3936 260708 3942
rect 260656 3878 260708 3884
rect 260668 480 260696 3878
rect 261772 480 261800 16546
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 262968 480 262996 3810
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 155382
rect 266004 155378 266032 157655
rect 266924 155446 266952 157791
rect 266912 155440 266964 155446
rect 266912 155382 266964 155388
rect 265992 155372 266044 155378
rect 265992 155314 266044 155320
rect 267660 155310 267688 158199
rect 268934 157856 268990 157865
rect 268934 157791 268990 157800
rect 268948 155582 268976 157791
rect 271064 156874 271092 159559
rect 275848 158846 275876 159559
rect 278148 158982 278176 159831
rect 300950 159760 301006 159769
rect 300950 159695 301006 159704
rect 279238 159624 279294 159633
rect 279238 159559 279294 159568
rect 288346 159624 288402 159633
rect 288346 159559 288402 159568
rect 295890 159624 295946 159633
rect 295890 159559 295946 159568
rect 279252 159050 279280 159559
rect 288360 159118 288388 159559
rect 295904 159186 295932 159559
rect 300964 159254 300992 159695
rect 322940 159656 322992 159662
rect 322940 159598 322992 159604
rect 318708 159588 318760 159594
rect 318708 159530 318760 159536
rect 314660 159520 314712 159526
rect 314660 159462 314712 159468
rect 310428 159452 310480 159458
rect 310428 159394 310480 159400
rect 305000 159384 305052 159390
rect 305000 159326 305052 159332
rect 300952 159248 301004 159254
rect 300952 159190 301004 159196
rect 295892 159180 295944 159186
rect 295892 159122 295944 159128
rect 288348 159112 288400 159118
rect 288348 159054 288400 159060
rect 279240 159044 279292 159050
rect 279240 158986 279292 158992
rect 278136 158976 278188 158982
rect 278136 158918 278188 158924
rect 277032 158908 277084 158914
rect 277032 158850 277084 158856
rect 275836 158840 275888 158846
rect 275836 158782 275888 158788
rect 274456 158772 274508 158778
rect 274456 158714 274508 158720
rect 274468 158681 274496 158714
rect 277044 158681 277072 158850
rect 305012 158710 305040 159326
rect 298560 158704 298612 158710
rect 271142 158672 271198 158681
rect 271142 158607 271198 158616
rect 272246 158672 272302 158681
rect 272246 158607 272302 158616
rect 274454 158672 274510 158681
rect 274454 158607 274510 158616
rect 277030 158672 277086 158681
rect 277030 158607 277086 158616
rect 298558 158672 298560 158681
rect 305000 158704 305052 158710
rect 298612 158672 298614 158681
rect 298558 158607 298614 158616
rect 303526 158672 303582 158681
rect 306104 158704 306156 158710
rect 305000 158646 305052 158652
rect 306102 158672 306104 158681
rect 306156 158672 306158 158681
rect 303526 158607 303582 158616
rect 306102 158607 306158 158616
rect 308770 158672 308826 158681
rect 308770 158607 308772 158616
rect 271156 158234 271184 158607
rect 271144 158228 271196 158234
rect 271144 158170 271196 158176
rect 272260 157894 272288 158607
rect 274454 158400 274510 158409
rect 274454 158335 274510 158344
rect 276110 158400 276166 158409
rect 276110 158335 276166 158344
rect 281354 158400 281410 158409
rect 281354 158335 281410 158344
rect 286322 158400 286378 158409
rect 286322 158335 286378 158344
rect 293682 158400 293738 158409
rect 293682 158335 293738 158344
rect 272248 157888 272300 157894
rect 272248 157830 272300 157836
rect 271052 156868 271104 156874
rect 271052 156810 271104 156816
rect 274468 156602 274496 158335
rect 274546 157720 274602 157729
rect 274546 157655 274602 157664
rect 274456 156596 274508 156602
rect 274456 156538 274508 156544
rect 267832 155576 267884 155582
rect 267832 155518 267884 155524
rect 268936 155576 268988 155582
rect 268936 155518 268988 155524
rect 266360 155304 266412 155310
rect 266360 155246 266412 155252
rect 267648 155304 267700 155310
rect 267648 155246 267700 155252
rect 266372 16574 266400 155246
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267844 6914 267872 155518
rect 269118 155408 269174 155417
rect 269118 155343 269174 155352
rect 269132 16574 269160 155343
rect 270498 155272 270554 155281
rect 274560 155242 274588 157655
rect 276124 156806 276152 158335
rect 278686 157720 278742 157729
rect 278686 157655 278742 157664
rect 276112 156800 276164 156806
rect 276112 156742 276164 156748
rect 270498 155207 270554 155216
rect 273260 155236 273312 155242
rect 270512 16574 270540 155207
rect 273260 155178 273312 155184
rect 274548 155236 274600 155242
rect 274548 155178 274600 155184
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 267752 6886 267872 6914
rect 267752 480 267780 6886
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 268856 480 268884 3742
rect 270052 480 270080 16546
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 3732 272484 3738
rect 272432 3674 272484 3680
rect 272444 480 272472 3674
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 155178
rect 278700 155174 278728 157655
rect 281368 156738 281396 158335
rect 283930 157584 283986 157593
rect 283930 157519 283986 157528
rect 281356 156732 281408 156738
rect 281356 156674 281408 156680
rect 277400 155168 277452 155174
rect 277400 155110 277452 155116
rect 278688 155168 278740 155174
rect 278688 155110 278740 155116
rect 274640 155032 274692 155038
rect 274640 154974 274692 154980
rect 274652 16574 274680 154974
rect 277412 16574 277440 155110
rect 283944 155106 283972 157519
rect 286336 156670 286364 158335
rect 291014 157584 291070 157593
rect 291014 157519 291070 157528
rect 286324 156664 286376 156670
rect 286324 156606 286376 156612
rect 278780 155100 278832 155106
rect 278780 155042 278832 155048
rect 283932 155100 283984 155106
rect 283932 155042 283984 155048
rect 278792 16574 278820 155042
rect 291028 155038 291056 157519
rect 293696 156534 293724 158335
rect 303540 158166 303568 158607
rect 308824 158607 308826 158616
rect 308772 158578 308824 158584
rect 310440 158166 310468 159394
rect 314672 158710 314700 159462
rect 314660 158704 314712 158710
rect 313462 158672 313518 158681
rect 314660 158646 314712 158652
rect 315854 158672 315910 158681
rect 313462 158607 313518 158616
rect 315854 158607 315910 158616
rect 318614 158672 318670 158681
rect 318720 158642 318748 159530
rect 321006 158672 321062 158681
rect 318614 158607 318670 158616
rect 318708 158636 318760 158642
rect 311070 158264 311126 158273
rect 311070 158199 311126 158208
rect 303528 158160 303580 158166
rect 303528 158102 303580 158108
rect 310428 158160 310480 158166
rect 310428 158102 310480 158108
rect 299478 157992 299534 158001
rect 299478 157927 299534 157936
rect 293684 156528 293736 156534
rect 293684 156470 293736 156476
rect 291016 155032 291068 155038
rect 291016 154974 291068 154980
rect 295340 154216 295392 154222
rect 295340 154158 295392 154164
rect 288440 154080 288492 154086
rect 288440 154022 288492 154028
rect 285680 153876 285732 153882
rect 285680 153818 285732 153824
rect 285692 16574 285720 153818
rect 288452 16574 288480 154022
rect 293960 153944 294012 153950
rect 293960 153886 294012 153892
rect 292578 153776 292634 153785
rect 292578 153711 292634 153720
rect 292592 16574 292620 153711
rect 293972 16574 294000 153886
rect 295352 16574 295380 154158
rect 298100 154012 298152 154018
rect 298100 153954 298152 153960
rect 274652 16546 274864 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 285692 16546 286640 16574
rect 288452 16546 289032 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 274836 480 274864 16546
rect 276020 3664 276072 3670
rect 276020 3606 276072 3612
rect 276032 480 276060 3606
rect 277124 3460 277176 3466
rect 277124 3402 277176 3408
rect 277136 480 277164 3402
rect 278332 480 278360 16546
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 285404 3664 285456 3670
rect 285404 3606 285456 3612
rect 284300 3596 284352 3602
rect 284300 3538 284352 3544
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 280724 480 280752 3470
rect 281920 480 281948 3470
rect 283104 3460 283156 3466
rect 283104 3402 283156 3408
rect 283116 480 283144 3402
rect 284312 480 284340 3538
rect 285416 480 285444 3606
rect 286612 480 286640 16546
rect 287796 3596 287848 3602
rect 287796 3538 287848 3544
rect 287808 480 287836 3538
rect 289004 480 289032 16546
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 290186 3360 290242 3369
rect 290186 3295 290242 3304
rect 290200 480 290228 3295
rect 291396 480 291424 3810
rect 292580 3800 292632 3806
rect 292580 3742 292632 3748
rect 292592 480 292620 3742
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297272 3392 297324 3398
rect 297272 3334 297324 3340
rect 297284 480 297312 3334
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 153954
rect 299492 3482 299520 157927
rect 311084 156466 311112 158199
rect 313476 158098 313504 158607
rect 313464 158092 313516 158098
rect 313464 158034 313516 158040
rect 315868 158030 315896 158607
rect 315856 158024 315908 158030
rect 315856 157966 315908 157972
rect 318628 157962 318656 158607
rect 321006 158607 321062 158616
rect 318708 158578 318760 158584
rect 321020 158166 321048 158607
rect 321008 158160 321060 158166
rect 321008 158102 321060 158108
rect 318616 157956 318668 157962
rect 318616 157898 318668 157904
rect 322952 157894 322980 159598
rect 356716 159390 356744 306462
rect 356796 306264 356848 306270
rect 356796 306206 356848 306212
rect 356704 159384 356756 159390
rect 356704 159326 356756 159332
rect 323398 158672 323454 158681
rect 323398 158607 323454 158616
rect 325974 158672 326030 158681
rect 325974 158607 326030 158616
rect 323412 157894 323440 158607
rect 322940 157888 322992 157894
rect 322940 157830 322992 157836
rect 323400 157888 323452 157894
rect 323400 157830 323452 157836
rect 325988 157826 326016 158607
rect 354126 158264 354182 158273
rect 354126 158199 354182 158208
rect 353942 158128 353998 158137
rect 353942 158063 353998 158072
rect 325976 157820 326028 157826
rect 325976 157762 326028 157768
rect 352562 156904 352618 156913
rect 352562 156839 352618 156848
rect 348422 156768 348478 156777
rect 348422 156703 348478 156712
rect 345662 156632 345718 156641
rect 345662 156567 345718 156576
rect 311072 156460 311124 156466
rect 311072 156402 311124 156408
rect 299572 154148 299624 154154
rect 299572 154090 299624 154096
rect 299584 3738 299612 154090
rect 319720 9444 319772 9450
rect 319720 9386 319772 9392
rect 316224 9376 316276 9382
rect 316224 9318 316276 9324
rect 303160 9240 303212 9246
rect 303160 9182 303212 9188
rect 301964 3936 302016 3942
rect 301964 3878 302016 3884
rect 299572 3732 299624 3738
rect 299572 3674 299624 3680
rect 300768 3732 300820 3738
rect 300768 3674 300820 3680
rect 301780 3732 301832 3738
rect 301780 3674 301832 3680
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3674
rect 301792 3398 301820 3674
rect 301780 3392 301832 3398
rect 301780 3334 301832 3340
rect 301976 480 302004 3878
rect 303172 480 303200 9182
rect 306748 9172 306800 9178
rect 306748 9114 306800 9120
rect 305552 9036 305604 9042
rect 305552 8978 305604 8984
rect 304356 8968 304408 8974
rect 304356 8910 304408 8916
rect 304368 480 304396 8910
rect 305564 480 305592 8978
rect 306760 480 306788 9114
rect 309048 9104 309100 9110
rect 309048 9046 309100 9052
rect 307944 6248 307996 6254
rect 307944 6190 307996 6196
rect 307956 480 307984 6190
rect 309060 480 309088 9046
rect 313832 6588 313884 6594
rect 313832 6530 313884 6536
rect 312636 6384 312688 6390
rect 312636 6326 312688 6332
rect 311440 6316 311492 6322
rect 311440 6258 311492 6264
rect 310244 6180 310296 6186
rect 310244 6122 310296 6128
rect 310256 480 310284 6122
rect 311452 480 311480 6258
rect 312648 480 312676 6326
rect 313844 480 313872 6530
rect 315028 6452 315080 6458
rect 315028 6394 315080 6400
rect 315040 480 315068 6394
rect 316236 480 316264 9318
rect 318524 6656 318576 6662
rect 318524 6598 318576 6604
rect 317328 6520 317380 6526
rect 317328 6462 317380 6468
rect 317340 480 317368 6462
rect 318536 480 318564 6598
rect 319732 480 319760 9386
rect 322112 9308 322164 9314
rect 322112 9250 322164 9256
rect 320914 6216 320970 6225
rect 320914 6151 320970 6160
rect 320928 480 320956 6151
rect 322124 480 322152 9250
rect 337476 6860 337528 6866
rect 337476 6802 337528 6808
rect 333888 6792 333940 6798
rect 333888 6734 333940 6740
rect 330392 6724 330444 6730
rect 330392 6666 330444 6672
rect 326802 6488 326858 6497
rect 326802 6423 326858 6432
rect 323306 6352 323362 6361
rect 323306 6287 323362 6296
rect 323320 480 323348 6287
rect 325606 3632 325662 3641
rect 325606 3567 325662 3576
rect 324410 3496 324466 3505
rect 324410 3431 324466 3440
rect 324424 480 324452 3431
rect 325620 480 325648 3567
rect 326816 480 326844 6423
rect 329196 4004 329248 4010
rect 329196 3946 329248 3952
rect 327998 3768 328054 3777
rect 327998 3703 328054 3712
rect 328012 480 328040 3703
rect 329208 480 329236 3946
rect 330404 480 330432 6666
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 331586 3904 331642 3913
rect 331586 3839 331642 3848
rect 331600 480 331628 3839
rect 332704 480 332732 4014
rect 333900 480 333928 6734
rect 336280 4140 336332 4146
rect 336280 4082 336332 4088
rect 335082 4040 335138 4049
rect 335082 3975 335138 3984
rect 335096 480 335124 3975
rect 336292 480 336320 4082
rect 337488 480 337516 6802
rect 340972 6112 341024 6118
rect 340972 6054 341024 6060
rect 338672 3392 338724 3398
rect 338672 3334 338724 3340
rect 338684 480 338712 3334
rect 339866 3224 339922 3233
rect 339866 3159 339922 3168
rect 339880 480 339908 3159
rect 340984 480 341012 6054
rect 344560 6044 344612 6050
rect 344560 5986 344612 5992
rect 343364 3324 343416 3330
rect 343364 3266 343416 3272
rect 342168 3256 342220 3262
rect 342168 3198 342220 3204
rect 342180 480 342208 3198
rect 343376 480 343404 3266
rect 344572 480 344600 5986
rect 345676 3670 345704 156567
rect 345756 154284 345808 154290
rect 345756 154226 345808 154232
rect 345768 3874 345796 154226
rect 348054 6624 348110 6633
rect 348054 6559 348110 6568
rect 345756 3868 345808 3874
rect 345756 3810 345808 3816
rect 345664 3664 345716 3670
rect 345664 3606 345716 3612
rect 346952 3664 347004 3670
rect 346952 3606 347004 3612
rect 345756 3188 345808 3194
rect 345756 3130 345808 3136
rect 345768 480 345796 3130
rect 346964 480 346992 3606
rect 348068 480 348096 6559
rect 348436 3806 348464 156703
rect 351642 6760 351698 6769
rect 351642 6695 351698 6704
rect 350448 5976 350500 5982
rect 350448 5918 350500 5924
rect 348424 3800 348476 3806
rect 348424 3742 348476 3748
rect 349252 3800 349304 3806
rect 349252 3742 349304 3748
rect 349264 480 349292 3742
rect 350460 480 350488 5918
rect 351656 480 351684 6695
rect 352576 3942 352604 156839
rect 352564 3936 352616 3942
rect 352564 3878 352616 3884
rect 353956 3738 353984 158063
rect 354036 3868 354088 3874
rect 354036 3810 354088 3816
rect 353944 3732 353996 3738
rect 353944 3674 353996 3680
rect 352840 3120 352892 3126
rect 352840 3062 352892 3068
rect 352852 480 352880 3062
rect 354048 480 354076 3810
rect 354140 3602 354168 158199
rect 356808 156913 356836 306206
rect 357176 302234 357204 308722
rect 357268 308582 357296 310420
rect 357256 308576 357308 308582
rect 357256 308518 357308 308524
rect 357452 306134 357480 310420
rect 357532 306604 357584 306610
rect 357532 306546 357584 306552
rect 357440 306128 357492 306134
rect 357440 306070 357492 306076
rect 357438 303376 357494 303385
rect 357438 303311 357494 303320
rect 356900 302206 357204 302234
rect 356900 243545 356928 302206
rect 356886 243536 356942 243545
rect 356886 243471 356942 243480
rect 357346 159624 357402 159633
rect 357346 159559 357402 159568
rect 357360 158953 357388 159559
rect 357346 158944 357402 158953
rect 357346 158879 357402 158888
rect 356794 156904 356850 156913
rect 356794 156839 356850 156848
rect 355966 3768 356022 3777
rect 355966 3703 356022 3712
rect 354128 3596 354180 3602
rect 354128 3538 354180 3544
rect 355232 3596 355284 3602
rect 355232 3538 355284 3544
rect 355244 480 355272 3538
rect 355980 3233 356008 3703
rect 356334 3632 356390 3641
rect 356334 3567 356390 3576
rect 355966 3224 356022 3233
rect 355966 3159 356022 3168
rect 356348 480 356376 3567
rect 357452 3534 357480 303311
rect 357544 158302 357572 306546
rect 357636 306474 357664 310420
rect 357624 306468 357676 306474
rect 357624 306410 357676 306416
rect 357820 306406 357848 310420
rect 358004 306610 358032 310420
rect 357992 306604 358044 306610
rect 357992 306546 358044 306552
rect 358188 306490 358216 310420
rect 358372 306513 358400 310420
rect 357912 306462 358216 306490
rect 358358 306504 358414 306513
rect 357808 306400 357860 306406
rect 357808 306342 357860 306348
rect 357716 306264 357768 306270
rect 357912 306218 357940 306462
rect 358358 306439 358414 306448
rect 357992 306400 358044 306406
rect 358556 306354 358584 310420
rect 357992 306342 358044 306348
rect 357716 306206 357768 306212
rect 357622 304328 357678 304337
rect 357622 304263 357678 304272
rect 357532 158296 357584 158302
rect 357532 158238 357584 158244
rect 357636 158234 357664 304263
rect 357728 158370 357756 306206
rect 357820 306190 357940 306218
rect 357820 159526 357848 306190
rect 357900 306128 357952 306134
rect 357900 306070 357952 306076
rect 357808 159520 357860 159526
rect 357808 159462 357860 159468
rect 357912 159254 357940 306070
rect 358004 159458 358032 306342
rect 358096 306326 358584 306354
rect 358096 159594 358124 306326
rect 358740 306218 358768 310420
rect 358188 306190 358768 306218
rect 358832 310406 359030 310434
rect 358188 159662 358216 306190
rect 358266 305960 358322 305969
rect 358266 305895 358322 305904
rect 358280 160177 358308 305895
rect 358832 301646 358860 310406
rect 359200 306354 359228 310420
rect 358924 306326 359228 306354
rect 358820 301640 358872 301646
rect 358820 301582 358872 301588
rect 358820 253088 358872 253094
rect 358820 253030 358872 253036
rect 358266 160168 358322 160177
rect 358266 160103 358322 160112
rect 358360 160132 358412 160138
rect 358360 160074 358412 160080
rect 358176 159656 358228 159662
rect 358176 159598 358228 159604
rect 358084 159588 358136 159594
rect 358084 159530 358136 159536
rect 357992 159452 358044 159458
rect 357992 159394 358044 159400
rect 357900 159248 357952 159254
rect 357900 159190 357952 159196
rect 358372 159066 358400 160074
rect 358280 159038 358400 159066
rect 357716 158364 357768 158370
rect 357716 158306 357768 158312
rect 357624 158228 357676 158234
rect 357624 158170 357676 158176
rect 358280 9246 358308 159038
rect 358358 158944 358414 158953
rect 358358 158879 358414 158888
rect 358268 9240 358320 9246
rect 358268 9182 358320 9188
rect 358372 6914 358400 158879
rect 357544 6886 358400 6914
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 357544 480 357572 6886
rect 358832 6322 358860 253030
rect 358924 156602 358952 306326
rect 359384 306218 359412 310420
rect 359568 306354 359596 310420
rect 359108 306190 359412 306218
rect 359476 306326 359596 306354
rect 359648 306400 359700 306406
rect 359648 306342 359700 306348
rect 359004 301640 359056 301646
rect 359004 301582 359056 301588
rect 358912 156596 358964 156602
rect 358912 156538 358964 156544
rect 359016 156466 359044 301582
rect 359108 158098 359136 306190
rect 359280 306128 359332 306134
rect 359280 306070 359332 306076
rect 359188 305448 359240 305454
rect 359188 305390 359240 305396
rect 359096 158092 359148 158098
rect 359096 158034 359148 158040
rect 359200 157962 359228 305390
rect 359292 158030 359320 306070
rect 359372 306060 359424 306066
rect 359372 306002 359424 306008
rect 359384 158846 359412 306002
rect 359372 158840 359424 158846
rect 359372 158782 359424 158788
rect 359476 158778 359504 306326
rect 359660 305726 359688 306342
rect 359752 306134 359780 310420
rect 359740 306128 359792 306134
rect 359740 306070 359792 306076
rect 359832 306128 359884 306134
rect 359832 306070 359884 306076
rect 359844 305862 359872 306070
rect 359936 306066 359964 310420
rect 359924 306060 359976 306066
rect 359924 306002 359976 306008
rect 359832 305856 359884 305862
rect 359832 305798 359884 305804
rect 359924 305856 359976 305862
rect 359924 305798 359976 305804
rect 359648 305720 359700 305726
rect 359648 305662 359700 305668
rect 359740 305720 359792 305726
rect 359740 305662 359792 305668
rect 359556 305380 359608 305386
rect 359556 305322 359608 305328
rect 359464 158772 359516 158778
rect 359464 158714 359516 158720
rect 359280 158024 359332 158030
rect 359280 157966 359332 157972
rect 359188 157956 359240 157962
rect 359188 157898 359240 157904
rect 359004 156460 359056 156466
rect 359004 156402 359056 156408
rect 359568 154494 359596 305322
rect 359752 305250 359780 305662
rect 359936 305590 359964 305798
rect 359924 305584 359976 305590
rect 359924 305526 359976 305532
rect 360016 305584 360068 305590
rect 360016 305526 360068 305532
rect 360028 305318 360056 305526
rect 360120 305454 360148 310420
rect 360200 308508 360252 308514
rect 360200 308450 360252 308456
rect 360212 306374 360240 308450
rect 360304 308038 360332 310420
rect 360488 308156 360516 310420
rect 360672 308394 360700 310420
rect 360856 308514 360884 310420
rect 360844 308508 360896 308514
rect 360844 308450 360896 308456
rect 361040 308394 361068 310420
rect 360672 308366 360792 308394
rect 360488 308128 360608 308156
rect 360292 308032 360344 308038
rect 360292 307974 360344 307980
rect 360476 307964 360528 307970
rect 360476 307906 360528 307912
rect 360212 306346 360424 306374
rect 360108 305448 360160 305454
rect 360108 305390 360160 305396
rect 360016 305312 360068 305318
rect 360016 305254 360068 305260
rect 359740 305244 359792 305250
rect 359740 305186 359792 305192
rect 360200 253156 360252 253162
rect 360200 253098 360252 253104
rect 359646 243672 359702 243681
rect 359646 243607 359702 243616
rect 359660 156641 359688 243607
rect 359646 156632 359702 156641
rect 359646 156567 359702 156576
rect 359556 154488 359608 154494
rect 359556 154430 359608 154436
rect 360212 6390 360240 253098
rect 360292 250844 360344 250850
rect 360292 250786 360344 250792
rect 360304 6594 360332 250786
rect 360396 157894 360424 306346
rect 360384 157888 360436 157894
rect 360384 157830 360436 157836
rect 360488 157826 360516 307906
rect 360580 158166 360608 308128
rect 360660 308032 360712 308038
rect 360660 307974 360712 307980
rect 360672 158914 360700 307974
rect 360764 158982 360792 308366
rect 360856 308366 361068 308394
rect 360856 159050 360884 308366
rect 361224 307970 361252 310420
rect 362130 309088 362186 309097
rect 362130 309023 362186 309032
rect 361212 307964 361264 307970
rect 361212 307906 361264 307912
rect 360936 307896 360988 307902
rect 360936 307838 360988 307844
rect 360844 159044 360896 159050
rect 360844 158986 360896 158992
rect 360752 158976 360804 158982
rect 360752 158918 360804 158924
rect 360660 158908 360712 158914
rect 360660 158850 360712 158856
rect 360568 158160 360620 158166
rect 360568 158102 360620 158108
rect 360476 157820 360528 157826
rect 360476 157762 360528 157768
rect 360948 156942 360976 307838
rect 361580 250436 361632 250442
rect 361580 250378 361632 250384
rect 361028 243704 361080 243710
rect 361028 243646 361080 243652
rect 360936 156936 360988 156942
rect 360936 156878 360988 156884
rect 361040 154086 361068 243646
rect 361028 154080 361080 154086
rect 361028 154022 361080 154028
rect 361592 6769 361620 250378
rect 362040 248124 362092 248130
rect 362040 248066 362092 248072
rect 361764 245472 361816 245478
rect 361764 245414 361816 245420
rect 361672 245336 361724 245342
rect 361672 245278 361724 245284
rect 361578 6760 361634 6769
rect 361578 6695 361634 6704
rect 360292 6588 360344 6594
rect 360292 6530 360344 6536
rect 360200 6384 360252 6390
rect 360200 6326 360252 6332
rect 358820 6316 358872 6322
rect 358820 6258 358872 6264
rect 358726 3496 358782 3505
rect 358726 3431 358782 3440
rect 359922 3496 359978 3505
rect 359922 3431 359978 3440
rect 361118 3496 361174 3505
rect 361118 3431 361174 3440
rect 358740 480 358768 3431
rect 359936 480 359964 3431
rect 361132 480 361160 3431
rect 361684 3262 361712 245278
rect 361672 3256 361724 3262
rect 361672 3198 361724 3204
rect 361776 3194 361804 245414
rect 361856 245404 361908 245410
rect 361856 245346 361908 245352
rect 361868 3806 361896 245346
rect 361948 245268 362000 245274
rect 361948 245210 362000 245216
rect 361856 3800 361908 3806
rect 361856 3742 361908 3748
rect 361960 3398 361988 245210
rect 362052 6458 362080 248066
rect 362144 159633 362172 309023
rect 362236 273970 362264 444042
rect 362316 441788 362368 441794
rect 362316 441730 362368 441736
rect 362328 325650 362356 441730
rect 362420 353258 362448 444110
rect 362500 443216 362552 443222
rect 362500 443158 362552 443164
rect 362512 405686 362540 443158
rect 362604 431934 362632 445946
rect 363604 445936 363656 445942
rect 363604 445878 363656 445884
rect 362592 431928 362644 431934
rect 362592 431870 362644 431876
rect 362500 405680 362552 405686
rect 362500 405622 362552 405628
rect 363616 365702 363644 445878
rect 378784 445868 378836 445874
rect 378784 445810 378836 445816
rect 374644 444780 374696 444786
rect 374644 444722 374696 444728
rect 371976 444712 372028 444718
rect 371976 444654 372028 444660
rect 363696 441924 363748 441930
rect 363696 441866 363748 441872
rect 363708 379506 363736 441866
rect 364984 440632 365036 440638
rect 364984 440574 365036 440580
rect 364996 419490 365024 440574
rect 364984 419484 365036 419490
rect 364984 419426 365036 419432
rect 363696 379500 363748 379506
rect 363696 379442 363748 379448
rect 363604 365696 363656 365702
rect 363604 365638 363656 365644
rect 362408 353252 362460 353258
rect 362408 353194 362460 353200
rect 362316 325644 362368 325650
rect 362316 325586 362368 325592
rect 367744 309120 367796 309126
rect 367744 309062 367796 309068
rect 366272 309052 366324 309058
rect 366272 308994 366324 309000
rect 364982 308952 365038 308961
rect 364982 308887 365038 308896
rect 364890 308816 364946 308825
rect 364890 308751 364946 308760
rect 364800 308168 364852 308174
rect 364800 308110 364852 308116
rect 363512 307828 363564 307834
rect 363512 307770 363564 307776
rect 362316 306536 362368 306542
rect 362316 306478 362368 306484
rect 362328 306066 362356 306478
rect 362316 306060 362368 306066
rect 362316 306002 362368 306008
rect 362316 302728 362368 302734
rect 362316 302670 362368 302676
rect 362224 273964 362276 273970
rect 362224 273906 362276 273912
rect 362224 243840 362276 243846
rect 362224 243782 362276 243788
rect 362130 159624 362186 159633
rect 362130 159559 362186 159568
rect 362236 154222 362264 243782
rect 362328 158438 362356 302670
rect 363144 251116 363196 251122
rect 363144 251058 363196 251064
rect 362960 248328 363012 248334
rect 362960 248270 363012 248276
rect 362408 243772 362460 243778
rect 362408 243714 362460 243720
rect 362316 158432 362368 158438
rect 362316 158374 362368 158380
rect 362420 156777 362448 243714
rect 362498 158944 362554 158953
rect 362498 158879 362554 158888
rect 362406 156768 362462 156777
rect 362406 156703 362462 156712
rect 362224 154216 362276 154222
rect 362224 154158 362276 154164
rect 362040 6452 362092 6458
rect 362040 6394 362092 6400
rect 362314 3496 362370 3505
rect 362314 3431 362370 3440
rect 361948 3392 362000 3398
rect 361948 3334 362000 3340
rect 361764 3188 361816 3194
rect 361764 3130 361816 3136
rect 362328 480 362356 3431
rect 362512 3126 362540 158879
rect 362972 4010 363000 248270
rect 363052 248192 363104 248198
rect 363052 248134 363104 248140
rect 363064 4078 363092 248134
rect 363156 6866 363184 251058
rect 363236 251048 363288 251054
rect 363236 250990 363288 250996
rect 363144 6860 363196 6866
rect 363144 6802 363196 6808
rect 363248 6798 363276 250990
rect 363328 250912 363380 250918
rect 363328 250854 363380 250860
rect 363236 6792 363288 6798
rect 363236 6734 363288 6740
rect 363340 6730 363368 250854
rect 363420 244520 363472 244526
rect 363420 244462 363472 244468
rect 363328 6724 363380 6730
rect 363328 6666 363380 6672
rect 363432 6526 363460 244462
rect 363524 157146 363552 307770
rect 363604 305584 363656 305590
rect 363604 305526 363656 305532
rect 363512 157140 363564 157146
rect 363512 157082 363564 157088
rect 363616 155786 363644 305526
rect 363696 303068 363748 303074
rect 363696 303010 363748 303016
rect 363708 158001 363736 303010
rect 364340 253904 364392 253910
rect 364340 253846 364392 253852
rect 363788 244316 363840 244322
rect 363788 244258 363840 244264
rect 363800 160138 363828 244258
rect 363878 160168 363934 160177
rect 363788 160132 363840 160138
rect 363878 160103 363934 160112
rect 363788 160074 363840 160080
rect 363694 157992 363750 158001
rect 363694 157927 363750 157936
rect 363786 157448 363842 157457
rect 363786 157383 363842 157392
rect 363604 155780 363656 155786
rect 363604 155722 363656 155728
rect 363420 6520 363472 6526
rect 363420 6462 363472 6468
rect 363052 4072 363104 4078
rect 363052 4014 363104 4020
rect 362960 4004 363012 4010
rect 362960 3946 363012 3952
rect 363800 3874 363828 157383
rect 363788 3868 363840 3874
rect 363788 3810 363840 3816
rect 363892 3670 363920 160103
rect 364352 6662 364380 253846
rect 364524 248396 364576 248402
rect 364524 248338 364576 248344
rect 364432 248260 364484 248266
rect 364432 248202 364484 248208
rect 364340 6656 364392 6662
rect 364340 6598 364392 6604
rect 364444 4146 364472 248202
rect 364432 4140 364484 4146
rect 364432 4082 364484 4088
rect 363880 3664 363932 3670
rect 363880 3606 363932 3612
rect 363510 3496 363566 3505
rect 363510 3431 363566 3440
rect 362500 3120 362552 3126
rect 362500 3062 362552 3068
rect 363524 480 363552 3431
rect 364536 3330 364564 248338
rect 364616 247648 364668 247654
rect 364616 247590 364668 247596
rect 364628 5982 364656 247590
rect 364708 243908 364760 243914
rect 364708 243850 364760 243856
rect 364720 9382 364748 243850
rect 364812 158506 364840 308110
rect 364904 158817 364932 308751
rect 364996 158953 365024 308887
rect 366180 308304 366232 308310
rect 366180 308246 366232 308252
rect 365076 305516 365128 305522
rect 365076 305458 365128 305464
rect 365088 159118 365116 305458
rect 365168 300620 365220 300626
rect 365168 300562 365220 300568
rect 365076 159112 365128 159118
rect 365076 159054 365128 159060
rect 364982 158944 365038 158953
rect 364982 158879 365038 158888
rect 364890 158808 364946 158817
rect 364890 158743 364946 158752
rect 364800 158500 364852 158506
rect 364800 158442 364852 158448
rect 365180 158273 365208 300562
rect 365812 253836 365864 253842
rect 365812 253778 365864 253784
rect 365720 251184 365772 251190
rect 365720 251126 365772 251132
rect 365166 158264 365222 158273
rect 365166 158199 365222 158208
rect 364708 9376 364760 9382
rect 364708 9318 364760 9324
rect 364616 5976 364668 5982
rect 364616 5918 364668 5924
rect 365732 3602 365760 251126
rect 365824 9450 365852 253778
rect 365996 250980 366048 250986
rect 365996 250922 366048 250928
rect 365904 250776 365956 250782
rect 365904 250718 365956 250724
rect 365812 9444 365864 9450
rect 365812 9386 365864 9392
rect 365916 6118 365944 250718
rect 365904 6112 365956 6118
rect 365904 6054 365956 6060
rect 366008 6050 366036 250922
rect 366088 246696 366140 246702
rect 366088 246638 366140 246644
rect 366100 8974 366128 246638
rect 366192 157078 366220 308246
rect 366180 157072 366232 157078
rect 366180 157014 366232 157020
rect 366284 157010 366312 308994
rect 367652 308984 367704 308990
rect 367652 308926 367704 308932
rect 367376 308712 367428 308718
rect 367376 308654 367428 308660
rect 367284 308236 367336 308242
rect 367284 308178 367336 308184
rect 366364 306332 366416 306338
rect 366364 306274 366416 306280
rect 366376 157214 366404 306274
rect 367100 303000 367152 303006
rect 367100 302942 367152 302948
rect 366456 302864 366508 302870
rect 366456 302806 366508 302812
rect 366468 157690 366496 302806
rect 366548 243636 366600 243642
rect 366548 243578 366600 243584
rect 366456 157684 366508 157690
rect 366456 157626 366508 157632
rect 366364 157208 366416 157214
rect 366364 157150 366416 157156
rect 366272 157004 366324 157010
rect 366272 156946 366324 156952
rect 366560 154290 366588 243578
rect 366548 154284 366600 154290
rect 366548 154226 366600 154232
rect 366088 8968 366140 8974
rect 366088 8910 366140 8916
rect 365996 6044 366048 6050
rect 365996 5986 366048 5992
rect 367006 3632 367062 3641
rect 365720 3596 365772 3602
rect 367006 3567 367062 3576
rect 365720 3538 365772 3544
rect 364614 3496 364670 3505
rect 364614 3431 364670 3440
rect 365810 3496 365866 3505
rect 365810 3431 365866 3440
rect 364524 3324 364576 3330
rect 364524 3266 364576 3272
rect 364628 480 364656 3431
rect 365824 480 365852 3431
rect 367020 480 367048 3567
rect 367112 3466 367140 302942
rect 367192 253768 367244 253774
rect 367192 253710 367244 253716
rect 367204 9042 367232 253710
rect 367296 155718 367324 308178
rect 367284 155712 367336 155718
rect 367284 155654 367336 155660
rect 367388 155378 367416 308654
rect 367560 308644 367612 308650
rect 367560 308586 367612 308592
rect 367468 308372 367520 308378
rect 367468 308314 367520 308320
rect 367480 155650 367508 308314
rect 367468 155644 367520 155650
rect 367468 155586 367520 155592
rect 367572 155514 367600 308586
rect 367664 157185 367692 308926
rect 367756 158574 367784 309062
rect 371424 308916 371476 308922
rect 371424 308858 371476 308864
rect 370134 308680 370190 308689
rect 370134 308615 370190 308624
rect 368572 308576 368624 308582
rect 368572 308518 368624 308524
rect 367928 303544 367980 303550
rect 367928 303486 367980 303492
rect 367836 302932 367888 302938
rect 367836 302874 367888 302880
rect 367744 158568 367796 158574
rect 367744 158510 367796 158516
rect 367650 157176 367706 157185
rect 367650 157111 367706 157120
rect 367560 155508 367612 155514
rect 367560 155450 367612 155456
rect 367376 155372 367428 155378
rect 367376 155314 367428 155320
rect 367848 153882 367876 302874
rect 367940 159225 367968 303486
rect 368480 253700 368532 253706
rect 368480 253642 368532 253648
rect 367926 159216 367982 159225
rect 367926 159151 367982 159160
rect 367836 153876 367888 153882
rect 367836 153818 367888 153824
rect 368492 9178 368520 253642
rect 368584 155310 368612 308518
rect 370044 308508 370096 308514
rect 370044 308450 370096 308456
rect 368662 306368 368718 306377
rect 368662 306303 368718 306312
rect 368676 155961 368704 306303
rect 368940 306196 368992 306202
rect 368940 306138 368992 306144
rect 368756 306060 368808 306066
rect 368756 306002 368808 306008
rect 368662 155952 368718 155961
rect 368662 155887 368718 155896
rect 368572 155304 368624 155310
rect 368572 155246 368624 155252
rect 368768 155242 368796 306002
rect 368846 305552 368902 305561
rect 368846 305487 368902 305496
rect 368860 155922 368888 305487
rect 368848 155916 368900 155922
rect 368848 155858 368900 155864
rect 368756 155236 368808 155242
rect 368756 155178 368808 155184
rect 368952 155174 368980 306138
rect 369032 306128 369084 306134
rect 369032 306070 369084 306076
rect 369044 156806 369072 306070
rect 369124 305856 369176 305862
rect 369124 305798 369176 305804
rect 369136 157282 369164 305798
rect 369216 300552 369268 300558
rect 369216 300494 369268 300500
rect 369228 158137 369256 300494
rect 369952 247580 370004 247586
rect 369952 247522 370004 247528
rect 369860 245608 369912 245614
rect 369860 245550 369912 245556
rect 369308 243568 369360 243574
rect 369308 243510 369360 243516
rect 369214 158128 369270 158137
rect 369214 158063 369270 158072
rect 369124 157276 369176 157282
rect 369124 157218 369176 157224
rect 369032 156800 369084 156806
rect 369032 156742 369084 156748
rect 368940 155168 368992 155174
rect 368940 155110 368992 155116
rect 369320 153950 369348 243510
rect 369308 153944 369360 153950
rect 369308 153886 369360 153892
rect 368480 9172 368532 9178
rect 368480 9114 368532 9120
rect 367192 9036 367244 9042
rect 367192 8978 367244 8984
rect 369872 6254 369900 245550
rect 369964 9110 369992 247522
rect 370056 155446 370084 308450
rect 370148 157321 370176 308615
rect 370318 306232 370374 306241
rect 370318 306167 370374 306176
rect 370228 305720 370280 305726
rect 370228 305662 370280 305668
rect 370134 157312 370190 157321
rect 370134 157247 370190 157256
rect 370240 155854 370268 305662
rect 370332 157049 370360 306167
rect 370412 305652 370464 305658
rect 370412 305594 370464 305600
rect 370424 157350 370452 305594
rect 370596 303408 370648 303414
rect 370596 303350 370648 303356
rect 370504 300484 370556 300490
rect 370504 300426 370556 300432
rect 370412 157344 370464 157350
rect 370412 157286 370464 157292
rect 370318 157040 370374 157049
rect 370318 156975 370374 156984
rect 370228 155848 370280 155854
rect 370228 155790 370280 155796
rect 370044 155440 370096 155446
rect 370044 155382 370096 155388
rect 370516 154154 370544 300426
rect 370608 159361 370636 303350
rect 370688 302796 370740 302802
rect 370688 302738 370740 302744
rect 370594 159352 370650 159361
rect 370594 159287 370650 159296
rect 370700 159186 370728 302738
rect 371240 286612 371292 286618
rect 371240 286554 371292 286560
rect 370688 159180 370740 159186
rect 370688 159122 370740 159128
rect 370504 154148 370556 154154
rect 370504 154090 370556 154096
rect 369952 9104 370004 9110
rect 369952 9046 370004 9052
rect 369860 6248 369912 6254
rect 369860 6190 369912 6196
rect 368202 3496 368258 3505
rect 367100 3460 367152 3466
rect 368202 3431 368258 3440
rect 369398 3496 369454 3505
rect 369398 3431 369454 3440
rect 370594 3496 370650 3505
rect 370594 3431 370650 3440
rect 367100 3402 367152 3408
rect 368216 480 368244 3431
rect 369412 480 369440 3431
rect 370608 480 370636 3431
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 286554
rect 371332 248056 371384 248062
rect 371332 247998 371384 248004
rect 371344 6186 371372 247998
rect 371436 154562 371464 308858
rect 371608 306264 371660 306270
rect 371608 306206 371660 306212
rect 371516 305992 371568 305998
rect 371516 305934 371568 305940
rect 371528 155106 371556 305934
rect 371620 156534 371648 306206
rect 371792 305924 371844 305930
rect 371792 305866 371844 305872
rect 371700 305788 371752 305794
rect 371700 305730 371752 305736
rect 371712 156738 371740 305730
rect 371700 156732 371752 156738
rect 371700 156674 371752 156680
rect 371804 156670 371832 305866
rect 371884 282464 371936 282470
rect 371884 282406 371936 282412
rect 371792 156664 371844 156670
rect 371792 156606 371844 156612
rect 371608 156528 371660 156534
rect 371608 156470 371660 156476
rect 371516 155100 371568 155106
rect 371516 155042 371568 155048
rect 371424 154556 371476 154562
rect 371424 154498 371476 154504
rect 371332 6180 371384 6186
rect 371332 6122 371384 6128
rect 371896 3194 371924 282406
rect 371988 167006 372016 444654
rect 373356 440496 373408 440502
rect 373356 440438 373408 440444
rect 373264 307352 373316 307358
rect 373264 307294 373316 307300
rect 372068 303612 372120 303618
rect 372068 303554 372120 303560
rect 371976 167000 372028 167006
rect 371976 166942 372028 166948
rect 372080 155038 372108 303554
rect 372804 303476 372856 303482
rect 372804 303418 372856 303424
rect 372620 254856 372672 254862
rect 372620 254798 372672 254804
rect 372068 155032 372120 155038
rect 372068 154974 372120 154980
rect 372632 6914 372660 254798
rect 372712 245540 372764 245546
rect 372712 245482 372764 245488
rect 372724 9314 372752 245482
rect 372816 155582 372844 303418
rect 372988 303204 373040 303210
rect 372988 303146 373040 303152
rect 372896 300416 372948 300422
rect 372896 300358 372948 300364
rect 372804 155576 372856 155582
rect 372804 155518 372856 155524
rect 372908 154018 372936 300358
rect 373000 157758 373028 303146
rect 372988 157752 373040 157758
rect 372988 157694 373040 157700
rect 372896 154012 372948 154018
rect 372896 153954 372948 153960
rect 372712 9308 372764 9314
rect 372712 9250 372764 9256
rect 372632 6886 372936 6914
rect 371884 3188 371936 3194
rect 371884 3130 371936 3136
rect 372908 480 372936 6886
rect 373276 3466 373304 307294
rect 373368 206990 373396 440438
rect 374184 303340 374236 303346
rect 374184 303282 374236 303288
rect 374000 301708 374052 301714
rect 374000 301650 374052 301656
rect 373356 206984 373408 206990
rect 373356 206926 373408 206932
rect 373264 3460 373316 3466
rect 373264 3402 373316 3408
rect 374012 3346 374040 301650
rect 374092 250708 374144 250714
rect 374092 250650 374144 250656
rect 374104 3534 374132 250650
rect 374196 156874 374224 303282
rect 374368 303272 374420 303278
rect 374368 303214 374420 303220
rect 374276 303136 374328 303142
rect 374276 303078 374328 303084
rect 374288 158545 374316 303078
rect 374380 159497 374408 303214
rect 374656 259418 374684 444722
rect 377404 440564 377456 440570
rect 377404 440506 377456 440512
rect 377416 313274 377444 440506
rect 377404 313268 377456 313274
rect 377404 313210 377456 313216
rect 376760 300688 376812 300694
rect 376760 300630 376812 300636
rect 374644 259412 374696 259418
rect 374644 259354 374696 259360
rect 374366 159488 374422 159497
rect 374366 159423 374422 159432
rect 374274 158536 374330 158545
rect 374274 158471 374330 158480
rect 374184 156868 374236 156874
rect 374184 156810 374236 156816
rect 376772 16574 376800 300630
rect 377404 298988 377456 298994
rect 377404 298930 377456 298936
rect 376772 16546 377352 16574
rect 374092 3528 374144 3534
rect 374092 3470 374144 3476
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 377324 3482 377352 16546
rect 377416 3602 377444 298930
rect 378140 285184 378192 285190
rect 378140 285126 378192 285132
rect 378152 16574 378180 285126
rect 378796 60722 378824 445810
rect 578884 444440 578936 444446
rect 578884 444382 578936 444388
rect 577502 443184 577558 443193
rect 388444 443148 388496 443154
rect 577502 443119 577558 443128
rect 388444 443090 388496 443096
rect 385040 298920 385092 298926
rect 385040 298862 385092 298868
rect 381544 297696 381596 297702
rect 381544 297638 381596 297644
rect 380900 294772 380952 294778
rect 380900 294714 380952 294720
rect 378784 60716 378836 60722
rect 378784 60658 378836 60664
rect 380912 16574 380940 294714
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 377404 3596 377456 3602
rect 377404 3538 377456 3544
rect 374012 3318 374132 3346
rect 374104 480 374132 3318
rect 375300 480 375328 3470
rect 377324 3454 377720 3482
rect 376484 3188 376536 3194
rect 376484 3130 376536 3136
rect 376496 480 376524 3130
rect 377692 480 377720 3454
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379978 3360 380034 3369
rect 379978 3295 380034 3304
rect 379992 480 380020 3295
rect 381188 480 381216 16546
rect 381556 3534 381584 297638
rect 382280 285116 382332 285122
rect 382280 285058 382332 285064
rect 381544 3528 381596 3534
rect 381544 3470 381596 3476
rect 382292 3398 382320 285058
rect 382372 264376 382424 264382
rect 382372 264318 382424 264324
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 264318
rect 385052 16574 385080 298862
rect 387064 292052 387116 292058
rect 387064 291994 387116 292000
rect 386420 271312 386472 271318
rect 386420 271254 386472 271260
rect 386432 16574 386460 271254
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 384764 3460 384816 3466
rect 384764 3402 384816 3408
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 384776 480 384804 3402
rect 385972 480 386000 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387076 3466 387104 291994
rect 387064 3460 387116 3466
rect 387064 3402 387116 3408
rect 388260 3460 388312 3466
rect 388260 3402 388312 3408
rect 388272 480 388300 3402
rect 388456 3398 388484 443090
rect 462962 308408 463018 308417
rect 462962 308343 463018 308352
rect 402980 307284 403032 307290
rect 402980 307226 403032 307232
rect 396722 303240 396778 303249
rect 396722 303175 396778 303184
rect 390560 283892 390612 283898
rect 390560 283834 390612 283840
rect 389180 263016 389232 263022
rect 389180 262958 389232 262964
rect 389192 16574 389220 262958
rect 389192 16546 389496 16574
rect 388444 3392 388496 3398
rect 388444 3334 388496 3340
rect 389468 480 389496 16546
rect 390572 3466 390600 283834
rect 390652 270020 390704 270026
rect 390652 269962 390704 269968
rect 390560 3460 390612 3466
rect 390560 3402 390612 3408
rect 390664 480 390692 269962
rect 393320 261792 393372 261798
rect 393320 261734 393372 261740
rect 391940 257440 391992 257446
rect 391940 257382 391992 257388
rect 391952 16574 391980 257382
rect 393332 16574 393360 261734
rect 396080 257372 396132 257378
rect 396080 257314 396132 257320
rect 394700 253632 394752 253638
rect 394700 253574 394752 253580
rect 394712 16574 394740 253574
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 391860 480 391888 3402
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 257314
rect 396736 2990 396764 303175
rect 400220 296200 400272 296206
rect 400220 296142 400272 296148
rect 397460 261724 397512 261730
rect 397460 261666 397512 261672
rect 397472 16574 397500 261666
rect 398840 258800 398892 258806
rect 398840 258742 398892 258748
rect 397472 16546 397776 16574
rect 396724 2984 396776 2990
rect 396724 2926 396776 2932
rect 397748 480 397776 16546
rect 398852 3398 398880 258742
rect 398932 253564 398984 253570
rect 398932 253506 398984 253512
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 253506
rect 400232 16574 400260 296142
rect 402992 16574 403020 307226
rect 427084 307216 427136 307222
rect 427084 307158 427136 307164
rect 422300 300348 422352 300354
rect 422300 300290 422352 300296
rect 412640 297628 412692 297634
rect 412640 297570 412692 297576
rect 405740 293548 405792 293554
rect 405740 293490 405792 293496
rect 405004 275528 405056 275534
rect 405004 275470 405056 275476
rect 404360 254788 404412 254794
rect 404360 254730 404412 254736
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 2984 402572 2990
rect 402520 2926 402572 2932
rect 402532 480 402560 2926
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 254730
rect 405016 3262 405044 275470
rect 405752 16574 405780 293490
rect 408500 290760 408552 290766
rect 408500 290702 408552 290708
rect 407212 276888 407264 276894
rect 407212 276830 407264 276836
rect 405752 16546 406056 16574
rect 405004 3256 405056 3262
rect 405004 3198 405056 3204
rect 406028 480 406056 16546
rect 407224 480 407252 276830
rect 408512 16574 408540 290702
rect 409880 279676 409932 279682
rect 409880 279618 409932 279624
rect 409892 16574 409920 279618
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 3256 408460 3262
rect 408408 3198 408460 3204
rect 408420 480 408448 3198
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 411916 480 411944 3538
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 297570
rect 421564 296132 421616 296138
rect 421564 296074 421616 296080
rect 418160 290624 418212 290630
rect 418160 290566 418212 290572
rect 414664 282396 414716 282402
rect 414664 282338 414716 282344
rect 413284 256216 413336 256222
rect 413284 256158 413336 256164
rect 413296 3058 413324 256158
rect 414020 249348 414072 249354
rect 414020 249290 414072 249296
rect 414032 16574 414060 249290
rect 414032 16546 414336 16574
rect 413284 3052 413336 3058
rect 413284 2994 413336 3000
rect 414308 480 414336 16546
rect 414676 3466 414704 282338
rect 417424 281036 417476 281042
rect 417424 280978 417476 280984
rect 416780 250640 416832 250646
rect 416780 250582 416832 250588
rect 416792 6914 416820 250582
rect 417436 16574 417464 280978
rect 418172 16574 418200 290566
rect 420920 264308 420972 264314
rect 420920 264250 420972 264256
rect 417436 16546 417556 16574
rect 418172 16546 418568 16574
rect 416792 6886 417464 6914
rect 414664 3460 414716 3466
rect 414664 3402 414716 3408
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 415492 3052 415544 3058
rect 415492 2994 415544 3000
rect 415504 480 415532 2994
rect 416700 480 416728 3402
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 6886
rect 417528 3058 417556 16546
rect 417516 3052 417568 3058
rect 417516 2994 417568 3000
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420184 3052 420236 3058
rect 420184 2994 420236 3000
rect 420196 480 420224 2994
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 264250
rect 421576 3602 421604 296074
rect 422312 16574 422340 300290
rect 423680 279608 423732 279614
rect 423680 279550 423732 279556
rect 422312 16546 422616 16574
rect 421564 3596 421616 3602
rect 421564 3538 421616 3544
rect 422588 480 422616 16546
rect 423692 3346 423720 279550
rect 425060 256148 425112 256154
rect 425060 256090 425112 256096
rect 423772 247988 423824 247994
rect 423772 247930 423824 247936
rect 423784 3534 423812 247930
rect 425072 16574 425100 256090
rect 425072 16546 425744 16574
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 423692 3318 423812 3346
rect 423784 480 423812 3318
rect 424980 480 425008 3470
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 427096 3670 427124 307158
rect 440884 304496 440936 304502
rect 440884 304438 440936 304444
rect 430580 289264 430632 289270
rect 430580 289206 430632 289212
rect 428464 278248 428516 278254
rect 428464 278190 428516 278196
rect 427820 252204 427872 252210
rect 427820 252146 427872 252152
rect 427832 6914 427860 252146
rect 428476 16574 428504 278190
rect 430592 16574 430620 289206
rect 435364 286544 435416 286550
rect 435364 286486 435416 286492
rect 434720 262948 434772 262954
rect 434720 262890 434772 262896
rect 431960 256080 432012 256086
rect 431960 256022 432012 256028
rect 428476 16546 428596 16574
rect 430592 16546 430896 16574
rect 427832 6886 428504 6914
rect 427084 3664 427136 3670
rect 427084 3606 427136 3612
rect 427268 3596 427320 3602
rect 427268 3538 427320 3544
rect 427280 480 427308 3538
rect 428476 480 428504 6886
rect 428568 4146 428596 16546
rect 428556 4140 428608 4146
rect 428556 4082 428608 4088
rect 429660 3392 429712 3398
rect 429660 3334 429712 3340
rect 429672 480 429700 3334
rect 430868 480 430896 16546
rect 431972 3534 432000 256022
rect 432052 252136 432104 252142
rect 432052 252078 432104 252084
rect 431960 3528 432012 3534
rect 431960 3470 432012 3476
rect 432064 480 432092 252078
rect 434732 16574 434760 262890
rect 434732 16546 435128 16574
rect 434444 4140 434496 4146
rect 434444 4082 434496 4088
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 433260 480 433288 3470
rect 434456 480 434484 4082
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426134 -960 426246 326
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 435376 3194 435404 286486
rect 436100 285048 436152 285054
rect 436100 284990 436152 284996
rect 436112 16574 436140 284990
rect 439504 276820 439556 276826
rect 439504 276762 439556 276768
rect 438860 246628 438912 246634
rect 438860 246570 438912 246576
rect 438872 16574 438900 246570
rect 436112 16546 436784 16574
rect 438872 16546 439176 16574
rect 435364 3188 435416 3194
rect 435364 3130 435416 3136
rect 436756 480 436784 16546
rect 437940 3188 437992 3194
rect 437940 3130 437992 3136
rect 437952 480 437980 3130
rect 439148 480 439176 16546
rect 439516 3534 439544 276762
rect 440896 3874 440924 304438
rect 452660 304428 452712 304434
rect 452660 304370 452712 304376
rect 448520 286476 448572 286482
rect 448520 286418 448572 286424
rect 442264 283756 442316 283762
rect 442264 283698 442316 283704
rect 441620 278180 441672 278186
rect 441620 278122 441672 278128
rect 441632 16574 441660 278122
rect 441632 16546 442212 16574
rect 440884 3868 440936 3874
rect 440884 3810 440936 3816
rect 440332 3664 440384 3670
rect 440332 3606 440384 3612
rect 439504 3528 439556 3534
rect 439504 3470 439556 3476
rect 440344 480 440372 3606
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442184 3482 442212 16546
rect 442276 3602 442304 283698
rect 445024 280968 445076 280974
rect 445024 280910 445076 280916
rect 443828 3868 443880 3874
rect 443828 3810 443880 3816
rect 442264 3596 442316 3602
rect 442264 3538 442316 3544
rect 441540 480 441568 3470
rect 442184 3454 442672 3482
rect 442644 480 442672 3454
rect 443840 480 443868 3810
rect 445036 3738 445064 280910
rect 446404 274236 446456 274242
rect 446404 274178 446456 274184
rect 445116 256012 445168 256018
rect 445116 255954 445168 255960
rect 445024 3732 445076 3738
rect 445024 3674 445076 3680
rect 445024 3596 445076 3602
rect 445024 3538 445076 3544
rect 445036 480 445064 3538
rect 445128 3126 445156 255954
rect 445760 245200 445812 245206
rect 445760 245142 445812 245148
rect 445116 3120 445168 3126
rect 445116 3062 445168 3068
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 245142
rect 446416 3330 446444 274178
rect 448532 3534 448560 286418
rect 448612 275460 448664 275466
rect 448612 275402 448664 275408
rect 448520 3528 448572 3534
rect 448520 3470 448572 3476
rect 446404 3324 446456 3330
rect 446404 3266 446456 3272
rect 447416 3120 447468 3126
rect 447416 3062 447468 3068
rect 447428 480 447456 3062
rect 448624 480 448652 275402
rect 449900 274168 449952 274174
rect 449900 274110 449952 274116
rect 449912 16574 449940 274110
rect 452672 16574 452700 304370
rect 460204 287836 460256 287842
rect 460204 287778 460256 287784
rect 458824 282328 458876 282334
rect 458824 282270 458876 282276
rect 454684 275392 454736 275398
rect 454684 275334 454736 275340
rect 454040 252000 454092 252006
rect 454040 251942 454092 251948
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449820 480 449848 3470
rect 450924 480 450952 16546
rect 452108 3324 452160 3330
rect 452108 3266 452160 3272
rect 452120 480 452148 3266
rect 453316 480 453344 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 251942
rect 454696 3534 454724 275334
rect 458180 249280 458232 249286
rect 458180 249222 458232 249228
rect 455420 247920 455472 247926
rect 455420 247862 455472 247868
rect 455432 16574 455460 247862
rect 458192 16574 458220 249222
rect 455432 16546 455736 16574
rect 458192 16546 458772 16574
rect 454684 3528 454736 3534
rect 454684 3470 454736 3476
rect 455708 480 455736 16546
rect 458088 3732 458140 3738
rect 458088 3674 458140 3680
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 456904 480 456932 3470
rect 458100 480 458128 3674
rect 458744 3482 458772 16546
rect 458836 3602 458864 282270
rect 459560 274100 459612 274106
rect 459560 274042 459612 274048
rect 459572 16574 459600 274042
rect 459572 16546 459968 16574
rect 458824 3596 458876 3602
rect 458824 3538 458876 3544
rect 458744 3454 459232 3482
rect 459204 480 459232 3454
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 460216 4146 460244 287778
rect 460940 249212 460992 249218
rect 460940 249154 460992 249160
rect 460952 16574 460980 249154
rect 460952 16546 461624 16574
rect 460204 4140 460256 4146
rect 460204 4082 460256 4088
rect 461596 480 461624 16546
rect 462780 4140 462832 4146
rect 462780 4082 462832 4088
rect 462792 480 462820 4082
rect 462976 3534 463004 308343
rect 480260 307148 480312 307154
rect 480260 307090 480312 307096
rect 476762 305824 476818 305833
rect 476762 305759 476818 305768
rect 463700 297492 463752 297498
rect 463700 297434 463752 297440
rect 463712 16574 463740 297434
rect 468484 294704 468536 294710
rect 468484 294646 468536 294652
rect 467104 293412 467156 293418
rect 467104 293354 467156 293360
rect 464344 291984 464396 291990
rect 464344 291926 464396 291932
rect 463712 16546 464016 16574
rect 462964 3528 463016 3534
rect 462964 3470 463016 3476
rect 463988 480 464016 16546
rect 464356 3058 464384 291926
rect 466460 251932 466512 251938
rect 466460 251874 466512 251880
rect 466472 16574 466500 251874
rect 466472 16546 467052 16574
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 3538
rect 467024 3482 467052 16546
rect 467116 3602 467144 293354
rect 467840 268456 467892 268462
rect 467840 268398 467892 268404
rect 467852 16574 467880 268398
rect 467852 16546 468248 16574
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 467024 3454 467512 3482
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 3454
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 4146 468524 294646
rect 471980 286408 472032 286414
rect 471980 286350 472032 286356
rect 471244 282260 471296 282266
rect 471244 282202 471296 282208
rect 468484 4140 468536 4146
rect 468484 4082 468536 4088
rect 471060 4140 471112 4146
rect 471060 4082 471112 4088
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 471072 480 471100 4082
rect 471256 3534 471284 282202
rect 471992 16574 472020 286350
rect 475384 272604 475436 272610
rect 475384 272546 475436 272552
rect 473452 268388 473504 268394
rect 473452 268330 473504 268336
rect 473464 16574 473492 268330
rect 474740 254720 474792 254726
rect 474740 254662 474792 254668
rect 474752 16574 474780 254662
rect 471992 16546 472296 16574
rect 473464 16546 474136 16574
rect 474752 16546 475332 16574
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 472268 480 472296 16546
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475304 3482 475332 16546
rect 475396 3602 475424 272546
rect 476776 3670 476804 305759
rect 478144 291916 478196 291922
rect 478144 291858 478196 291864
rect 477500 249144 477552 249150
rect 477500 249086 477552 249092
rect 477512 6914 477540 249086
rect 478156 16574 478184 291858
rect 480272 16574 480300 307090
rect 543740 307080 543792 307086
rect 543740 307022 543792 307028
rect 485044 304360 485096 304366
rect 485044 304302 485096 304308
rect 481732 280900 481784 280906
rect 481732 280842 481784 280848
rect 478156 16546 478276 16574
rect 480272 16546 480576 16574
rect 477512 6886 478184 6914
rect 476764 3664 476816 3670
rect 476764 3606 476816 3612
rect 475384 3596 475436 3602
rect 475384 3538 475436 3544
rect 476948 3596 477000 3602
rect 476948 3538 477000 3544
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 476960 480 476988 3538
rect 478156 480 478184 6886
rect 478248 4146 478276 16546
rect 478236 4140 478288 4146
rect 478236 4082 478288 4088
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481744 480 481772 280842
rect 484400 271244 484452 271250
rect 484400 271186 484452 271192
rect 484412 16574 484440 271186
rect 484412 16546 484808 16574
rect 482836 4140 482888 4146
rect 482836 4082 482888 4088
rect 482848 480 482876 4082
rect 484032 3596 484084 3602
rect 484032 3538 484084 3544
rect 484044 480 484072 3538
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485056 3194 485084 304302
rect 514024 304292 514076 304298
rect 514024 304234 514076 304240
rect 489182 303104 489238 303113
rect 489182 303039 489238 303048
rect 486424 269952 486476 269958
rect 486424 269894 486476 269900
rect 485780 261588 485832 261594
rect 485780 261530 485832 261536
rect 485792 6914 485820 261530
rect 486436 16574 486464 269894
rect 486436 16546 486556 16574
rect 485792 6886 486464 6914
rect 485044 3188 485096 3194
rect 485044 3130 485096 3136
rect 486436 480 486464 6886
rect 486528 3058 486556 16546
rect 489196 3738 489224 303039
rect 494060 301572 494112 301578
rect 494060 301514 494112 301520
rect 490012 289196 490064 289202
rect 490012 289138 490064 289144
rect 490024 6914 490052 289138
rect 493324 279540 493376 279546
rect 493324 279482 493376 279488
rect 491300 265804 491352 265810
rect 491300 265746 491352 265752
rect 491312 16574 491340 265746
rect 492680 250572 492732 250578
rect 492680 250514 492732 250520
rect 492692 16574 492720 250514
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 489932 6886 490052 6914
rect 489184 3732 489236 3738
rect 489184 3674 489236 3680
rect 487620 3188 487672 3194
rect 487620 3130 487672 3136
rect 486516 3052 486568 3058
rect 486516 2994 486568 3000
rect 487632 480 487660 3130
rect 488816 3052 488868 3058
rect 488816 2994 488868 3000
rect 488828 480 488856 2994
rect 489932 480 489960 6886
rect 491116 3732 491168 3738
rect 491116 3674 491168 3680
rect 491128 480 491156 3674
rect 492324 480 492352 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 493336 3398 493364 279482
rect 494072 16574 494100 301514
rect 498292 300280 498344 300286
rect 498292 300222 498344 300228
rect 495440 267164 495492 267170
rect 495440 267106 495492 267112
rect 494072 16546 494744 16574
rect 493324 3392 493376 3398
rect 493324 3334 493376 3340
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 267106
rect 496084 253428 496136 253434
rect 496084 253370 496136 253376
rect 496096 3534 496124 253370
rect 498304 6914 498332 300222
rect 500224 298852 500276 298858
rect 500224 298794 500276 298800
rect 499580 253360 499632 253366
rect 499580 253302 499632 253308
rect 499592 16574 499620 253302
rect 499592 16546 500172 16574
rect 498212 6886 498332 6914
rect 496084 3528 496136 3534
rect 496084 3470 496136 3476
rect 497096 3528 497148 3534
rect 497096 3470 497148 3476
rect 497108 480 497136 3470
rect 498212 480 498240 6886
rect 500144 3482 500172 16546
rect 500236 3602 500264 298794
rect 509884 293344 509936 293350
rect 509884 293286 509936 293292
rect 506480 253292 506532 253298
rect 506480 253234 506532 253240
rect 502340 247852 502392 247858
rect 502340 247794 502392 247800
rect 502352 16574 502380 247794
rect 505100 246560 505152 246566
rect 505100 246502 505152 246508
rect 503720 245132 503772 245138
rect 503720 245074 503772 245080
rect 502352 16546 503024 16574
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 500144 3454 500632 3482
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500604 480 500632 3454
rect 501800 480 501828 3538
rect 502996 480 503024 16546
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 245074
rect 505112 16574 505140 246502
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 3534 506520 253234
rect 509240 251864 509292 251870
rect 509240 251806 509292 251812
rect 507860 246492 507912 246498
rect 507860 246434 507912 246440
rect 506572 245064 506624 245070
rect 506572 245006 506624 245012
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3380 506612 245006
rect 507872 16574 507900 246434
rect 509252 16574 509280 251806
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3352 506612 3380
rect 506492 480 506520 3352
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 509896 3330 509924 293286
rect 511264 278112 511316 278118
rect 511264 278054 511316 278060
rect 510620 246424 510672 246430
rect 510620 246366 510672 246372
rect 510632 16574 510660 246366
rect 510632 16546 511212 16574
rect 511184 3482 511212 16546
rect 511276 3602 511304 278054
rect 512000 247784 512052 247790
rect 512000 247726 512052 247732
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511184 3454 511304 3482
rect 509884 3324 509936 3330
rect 509884 3266 509936 3272
rect 511276 480 511304 3454
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 247726
rect 513564 3596 513616 3602
rect 513564 3538 513616 3544
rect 513576 480 513604 3538
rect 514036 3058 514064 304234
rect 520922 302968 520978 302977
rect 520922 302903 520978 302912
rect 516784 296064 516836 296070
rect 516784 296006 516836 296012
rect 516140 246356 516192 246362
rect 516140 246298 516192 246304
rect 516152 16574 516180 246298
rect 516152 16546 516732 16574
rect 516704 3482 516732 16546
rect 516796 3874 516824 296006
rect 517520 269884 517572 269890
rect 517520 269826 517572 269832
rect 517532 16574 517560 269826
rect 520280 249076 520332 249082
rect 520280 249018 520332 249024
rect 517532 16546 517928 16574
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 516704 3454 517192 3482
rect 514760 3324 514812 3330
rect 514760 3266 514812 3272
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 3266
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 3454
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3868 519596 3874
rect 519544 3810 519596 3816
rect 519556 480 519584 3810
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 249018
rect 520936 3534 520964 302903
rect 539690 302832 539746 302841
rect 539690 302767 539746 302776
rect 529940 301504 529992 301510
rect 529940 301446 529992 301452
rect 525800 294636 525852 294642
rect 525800 294578 525852 294584
rect 521660 283688 521712 283694
rect 521660 283630 521712 283636
rect 520924 3528 520976 3534
rect 520924 3470 520976 3476
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 283630
rect 522304 276752 522356 276758
rect 522304 276694 522356 276700
rect 522316 3058 522344 276694
rect 525064 275324 525116 275330
rect 525064 275266 525116 275272
rect 524420 247716 524472 247722
rect 524420 247658 524472 247664
rect 524432 16574 524460 247658
rect 524432 16546 525012 16574
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 524984 3482 525012 16546
rect 525076 3602 525104 275266
rect 525812 16574 525840 294578
rect 527824 293276 527876 293282
rect 527824 293218 527876 293224
rect 525812 16546 526208 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 522304 3052 522356 3058
rect 522304 2994 522356 3000
rect 523052 480 523080 3470
rect 524984 3454 525472 3482
rect 524236 3052 524288 3058
rect 524236 2994 524288 3000
rect 524248 480 524276 2994
rect 525444 480 525472 3454
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527732 3596 527784 3602
rect 527732 3538 527784 3544
rect 527744 3346 527772 3538
rect 527836 3534 527864 293218
rect 528560 253224 528612 253230
rect 528560 253166 528612 253172
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 527744 3318 527864 3346
rect 527836 480 527864 3318
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 253166
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 301446
rect 538864 300212 538916 300218
rect 538864 300154 538916 300160
rect 534724 291848 534776 291854
rect 534724 291790 534776 291796
rect 531320 279472 531372 279478
rect 531320 279414 531372 279420
rect 531332 3534 531360 279414
rect 531412 274032 531464 274038
rect 531412 273974 531464 273980
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 273974
rect 534080 244996 534132 245002
rect 534080 244938 534132 244944
rect 534092 16574 534120 244938
rect 534092 16546 534488 16574
rect 533712 3596 533764 3602
rect 533712 3538 533764 3544
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 3538
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3194 534764 291790
rect 536104 283620 536156 283626
rect 536104 283562 536156 283568
rect 535460 265736 535512 265742
rect 535460 265678 535512 265684
rect 535472 6914 535500 265678
rect 536116 16574 536144 283562
rect 536116 16546 536236 16574
rect 535472 6886 536144 6914
rect 534724 3188 534776 3194
rect 534724 3130 534776 3136
rect 536116 480 536144 6886
rect 536208 4146 536236 16546
rect 536196 4140 536248 4146
rect 536196 4082 536248 4088
rect 538404 4140 538456 4146
rect 538404 4082 538456 4088
rect 537208 3188 537260 3194
rect 537208 3130 537260 3136
rect 537220 480 537248 3130
rect 538416 480 538444 4082
rect 538876 3058 538904 300154
rect 539704 6914 539732 302767
rect 543004 290556 543056 290562
rect 543004 290498 543056 290504
rect 540244 272536 540296 272542
rect 540244 272478 540296 272484
rect 539612 6886 539732 6914
rect 538864 3052 538916 3058
rect 538864 2994 538916 3000
rect 539612 480 539640 6886
rect 540256 2990 540284 272478
rect 542360 260228 542412 260234
rect 542360 260170 542412 260176
rect 542372 16574 542400 260170
rect 542372 16546 542768 16574
rect 540796 3052 540848 3058
rect 540796 2994 540848 3000
rect 540244 2984 540296 2990
rect 540244 2926 540296 2932
rect 540808 480 540836 2994
rect 541992 2984 542044 2990
rect 541992 2926 542044 2932
rect 542004 480 542032 2926
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3398 543044 290498
rect 543752 16574 543780 307022
rect 570602 305688 570658 305697
rect 570602 305623 570658 305632
rect 545764 300144 545816 300150
rect 545764 300086 545816 300092
rect 545120 271176 545172 271182
rect 545120 271118 545172 271124
rect 545132 16574 545160 271118
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 543004 3392 543056 3398
rect 543004 3334 543056 3340
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 545776 3534 545804 300086
rect 547972 298784 548024 298790
rect 547972 298726 548024 298732
rect 547984 6914 548012 298726
rect 557540 297424 557592 297430
rect 557540 297366 557592 297372
rect 549904 290488 549956 290494
rect 549904 290430 549956 290436
rect 549260 264240 549312 264246
rect 549260 264182 549312 264188
rect 549272 16574 549300 264182
rect 549272 16546 549852 16574
rect 547892 6886 548012 6914
rect 545764 3528 545816 3534
rect 545764 3470 545816 3476
rect 546684 3528 546736 3534
rect 546684 3470 546736 3476
rect 546696 480 546724 3470
rect 547892 480 547920 6886
rect 549824 3482 549852 16546
rect 549916 3602 549944 290430
rect 552664 289128 552716 289134
rect 552664 289070 552716 289076
rect 552020 269816 552072 269822
rect 552020 269758 552072 269764
rect 552032 6914 552060 269758
rect 552676 16574 552704 289070
rect 554044 287768 554096 287774
rect 554044 287710 554096 287716
rect 553400 267096 553452 267102
rect 553400 267038 553452 267044
rect 553412 16574 553440 267038
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 549904 3596 549956 3602
rect 549904 3538 549956 3544
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 549824 3454 550312 3482
rect 549076 3392 549128 3398
rect 549076 3334 549128 3340
rect 549088 480 549116 3334
rect 550284 480 550312 3454
rect 551480 480 551508 3538
rect 552676 480 552704 6886
rect 552768 2990 552796 16546
rect 552756 2984 552808 2990
rect 552756 2926 552808 2932
rect 553780 480 553808 16546
rect 554056 3262 554084 287710
rect 556252 282192 556304 282198
rect 556252 282134 556304 282140
rect 556264 6914 556292 282134
rect 557552 16574 557580 297366
rect 563704 295996 563756 296002
rect 563704 295938 563756 295944
rect 561680 287700 561732 287706
rect 561680 287642 561732 287648
rect 560300 276684 560352 276690
rect 560300 276626 560352 276632
rect 558920 260160 558972 260166
rect 558920 260102 558972 260108
rect 558932 16574 558960 260102
rect 560312 16574 560340 276626
rect 560944 265668 560996 265674
rect 560944 265610 560996 265616
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 556172 6886 556292 6914
rect 554044 3256 554096 3262
rect 554044 3198 554096 3204
rect 554964 2984 555016 2990
rect 554964 2926 555016 2932
rect 554976 480 555004 2926
rect 556172 480 556200 6886
rect 557356 3256 557408 3262
rect 557356 3198 557408 3204
rect 557368 480 557396 3198
rect 558564 480 558592 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 560956 3194 560984 265610
rect 561692 16574 561720 287642
rect 561692 16546 562088 16574
rect 560944 3188 560996 3194
rect 560944 3130 560996 3136
rect 562060 480 562088 16546
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 563716 3058 563744 295938
rect 566464 286340 566516 286346
rect 566464 286282 566516 286288
rect 565820 267028 565872 267034
rect 565820 266970 565872 266976
rect 564532 254652 564584 254658
rect 564532 254594 564584 254600
rect 564544 6914 564572 254594
rect 565832 16574 565860 266970
rect 565832 16546 566412 16574
rect 564452 6886 564572 6914
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 564452 480 564480 6886
rect 566384 3482 566412 16546
rect 566476 3874 566504 286282
rect 569960 261520 570012 261526
rect 569960 261462 570012 261468
rect 567200 254584 567252 254590
rect 567200 254526 567252 254532
rect 567212 16574 567240 254526
rect 569972 16574 570000 261462
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 566464 3868 566516 3874
rect 566464 3810 566516 3816
rect 566384 3454 566872 3482
rect 565636 3052 565688 3058
rect 565636 2994 565688 3000
rect 565648 480 565676 2994
rect 566844 480 566872 3454
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 3868 569184 3874
rect 569132 3810 569184 3816
rect 569144 480 569172 3810
rect 570340 480 570368 16546
rect 570616 3534 570644 305623
rect 575480 284980 575532 284986
rect 575480 284922 575532 284928
rect 571984 280832 572036 280838
rect 571984 280774 572036 280780
rect 571340 244928 571392 244934
rect 571340 244870 571392 244876
rect 570604 3528 570656 3534
rect 570604 3470 570656 3476
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 244870
rect 571996 3058 572024 280774
rect 574100 262880 574152 262886
rect 574100 262822 574152 262828
rect 574112 16574 574140 262822
rect 575492 16574 575520 284922
rect 576860 250504 576912 250510
rect 576860 250446 576912 250452
rect 576872 16574 576900 250446
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 3470
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 577516 6798 577544 443119
rect 577596 441652 577648 441658
rect 577596 441594 577648 441600
rect 577608 193186 577636 441594
rect 578240 278044 578292 278050
rect 578240 277986 578292 277992
rect 577596 193180 577648 193186
rect 577596 193122 577648 193128
rect 578252 16574 578280 277986
rect 578896 245585 578924 444382
rect 581092 443080 581144 443086
rect 580354 443048 580410 443057
rect 581092 443022 581144 443028
rect 580354 442983 580410 442992
rect 580264 442536 580316 442542
rect 580264 442478 580316 442484
rect 580172 440904 580224 440910
rect 580172 440846 580224 440852
rect 579804 431928 579856 431934
rect 579804 431870 579856 431876
rect 579816 431633 579844 431870
rect 579802 431624 579858 431633
rect 579802 431559 579858 431568
rect 579988 419484 580040 419490
rect 579988 419426 580040 419432
rect 580000 418305 580028 419426
rect 579986 418296 580042 418305
rect 579986 418231 580042 418240
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404977 579844 405622
rect 579802 404968 579858 404977
rect 579802 404903 579858 404912
rect 580080 379500 580132 379506
rect 580080 379442 580132 379448
rect 580092 378457 580120 379442
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580080 365696 580132 365702
rect 580080 365638 580132 365644
rect 580092 365129 580120 365638
rect 580078 365120 580134 365129
rect 580078 365055 580134 365064
rect 579988 353252 580040 353258
rect 579988 353194 580040 353200
rect 580000 351937 580028 353194
rect 579986 351928 580042 351937
rect 579986 351863 580042 351872
rect 580080 325644 580132 325650
rect 580080 325586 580132 325592
rect 580092 325281 580120 325586
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 579988 313268 580040 313274
rect 579988 313210 580040 313216
rect 580000 312089 580028 313210
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580184 298761 580212 440846
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273964 580224 273970
rect 580172 273906 580224 273912
rect 580184 272241 580212 273906
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 578882 245576 578938 245585
rect 578882 245511 578938 245520
rect 579620 206984 579672 206990
rect 579620 206926 579672 206932
rect 579632 205737 579660 206926
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580276 19825 580304 442478
rect 580368 33153 580396 442983
rect 580724 442672 580776 442678
rect 580724 442614 580776 442620
rect 580632 442604 580684 442610
rect 580632 442546 580684 442552
rect 580540 442332 580592 442338
rect 580540 442274 580592 442280
rect 580448 442264 580500 442270
rect 580448 442206 580500 442212
rect 580460 73001 580488 442206
rect 580552 112849 580580 442274
rect 580644 139369 580672 442546
rect 580736 152697 580764 442614
rect 580816 442468 580868 442474
rect 580816 442410 580868 442416
rect 580828 219065 580856 442410
rect 580908 442400 580960 442406
rect 580908 442342 580960 442348
rect 580920 232393 580948 442342
rect 580906 232384 580962 232393
rect 580906 232319 580962 232328
rect 580814 219056 580870 219065
rect 580814 218991 580870 219000
rect 580816 193180 580868 193186
rect 580816 193122 580868 193128
rect 580828 192545 580856 193122
rect 580814 192536 580870 192545
rect 580814 192471 580870 192480
rect 580722 152688 580778 152697
rect 580722 152623 580778 152632
rect 580630 139360 580686 139369
rect 580630 139295 580686 139304
rect 580538 112840 580594 112849
rect 580538 112775 580594 112784
rect 580446 72992 580502 73001
rect 580446 72927 580502 72936
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 581104 16574 581132 443022
rect 582380 443012 582432 443018
rect 582380 442954 582432 442960
rect 582392 16574 582420 442954
rect 578252 16546 578648 16574
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 577504 6792 577556 6798
rect 577504 6734 577556 6740
rect 578620 480 578648 16546
rect 580264 6792 580316 6798
rect 580264 6734 580316 6740
rect 580276 6633 580304 6734
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3146 619112 3202 619168
rect 3422 606076 3478 606112
rect 3422 606056 3424 606076
rect 3424 606056 3476 606076
rect 3476 606056 3478 606076
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 217598 516840 217654 516896
rect 217506 513712 217562 513768
rect 217414 489912 217470 489968
rect 217322 488008 217378 488064
rect 4066 449520 4122 449576
rect 217690 515888 217746 515944
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3330 254088 3386 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3698 358400 3754 358456
rect 3606 345344 3662 345400
rect 3514 241032 3570 241088
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 34518 300056 34574 300112
rect 134154 372680 134210 372736
rect 159914 374040 159970 374096
rect 133878 371612 133934 371648
rect 133878 371592 133886 371612
rect 133886 371592 133934 371612
rect 135166 371628 135168 371648
rect 135168 371628 135220 371648
rect 135220 371628 135222 371648
rect 135166 371592 135222 371628
rect 143262 371612 143318 371648
rect 143262 371592 143264 371612
rect 143264 371592 143316 371612
rect 143316 371592 143318 371612
rect 153014 371628 153016 371648
rect 153016 371628 153068 371648
rect 153068 371628 153070 371648
rect 153014 371592 153070 371628
rect 99838 370640 99894 370696
rect 97906 367376 97962 367432
rect 97814 364656 97870 364712
rect 97722 361936 97778 361992
rect 99286 359216 99342 359272
rect 99194 356496 99250 356552
rect 97906 353776 97962 353832
rect 97630 351056 97686 351112
rect 97814 345616 97870 345672
rect 97722 340176 97778 340232
rect 97630 334736 97686 334792
rect 97538 332016 97594 332072
rect 97446 326576 97502 326632
rect 97354 323856 97410 323912
rect 97262 310256 97318 310312
rect 97262 299104 97318 299160
rect 99102 348336 99158 348392
rect 99010 342896 99066 342952
rect 98918 337456 98974 337512
rect 98826 329296 98882 329352
rect 98734 321136 98790 321192
rect 98642 315696 98698 315752
rect 98550 307536 98606 307592
rect 97906 304816 97962 304872
rect 97538 299376 97594 299432
rect 97354 298016 97410 298072
rect 99378 318416 99434 318472
rect 99286 300736 99342 300792
rect 99470 312976 99526 313032
rect 170770 309440 170826 309496
rect 171690 358536 171746 358592
rect 172334 369416 172390 369472
rect 172426 366696 172482 366752
rect 171874 363976 171930 364032
rect 170954 309304 171010 309360
rect 99838 302096 99894 302152
rect 164238 300328 164294 300384
rect 160098 300192 160154 300248
rect 99194 299240 99250 299296
rect 109682 297880 109738 297936
rect 150898 297744 150954 297800
rect 170494 302912 170550 302968
rect 171966 361256 172022 361312
rect 171874 350376 171930 350432
rect 171414 325896 171470 325952
rect 172426 355816 172482 355872
rect 172426 353096 172482 353152
rect 172426 347656 172482 347712
rect 172058 344936 172114 344992
rect 172426 342252 172428 342272
rect 172428 342252 172480 342272
rect 172480 342252 172482 342272
rect 172426 342216 172482 342252
rect 172150 339496 172206 339552
rect 172426 336796 172482 336832
rect 172426 336776 172428 336796
rect 172428 336776 172480 336796
rect 172480 336776 172482 336796
rect 172426 334056 172482 334112
rect 172426 331336 172482 331392
rect 172426 328616 172482 328672
rect 172242 323176 172298 323232
rect 172058 310800 172114 310856
rect 172426 320456 172482 320512
rect 172426 317736 172482 317792
rect 172426 315016 172482 315072
rect 172426 312296 172482 312352
rect 172426 309576 172482 309632
rect 174726 309168 174782 309224
rect 174634 308896 174690 308952
rect 173254 308216 173310 308272
rect 172426 306856 172482 306912
rect 172334 304136 172390 304192
rect 172426 301416 172482 301472
rect 182178 302776 182234 302832
rect 205086 3304 205142 3360
rect 210974 155352 211030 155408
rect 210790 155216 210846 155272
rect 211986 297472 212042 297528
rect 212354 297336 212410 297392
rect 212170 3576 212226 3632
rect 213550 297608 213606 297664
rect 214746 157800 214802 157856
rect 214470 3440 214526 3496
rect 219162 512760 219218 512816
rect 219070 509904 219126 509960
rect 218978 508136 219034 508192
rect 218886 488280 218942 488336
rect 219254 510992 219310 511048
rect 238482 477264 238538 477320
rect 242806 477128 242862 477184
rect 240046 476856 240102 476912
rect 241426 476876 241482 476912
rect 241426 476856 241428 476876
rect 241428 476856 241480 476876
rect 241480 476856 241482 476876
rect 237286 476740 237342 476776
rect 237286 476720 237288 476740
rect 237288 476720 237340 476740
rect 237340 476720 237342 476740
rect 237194 476176 237250 476232
rect 256606 476992 256662 477048
rect 253754 476448 253810 476504
rect 245474 476312 245530 476368
rect 248326 476312 248382 476368
rect 251086 476312 251142 476368
rect 252374 476312 252430 476368
rect 244186 476176 244242 476232
rect 245566 476176 245622 476232
rect 246946 476176 247002 476232
rect 248234 476176 248290 476232
rect 249706 476176 249762 476232
rect 250994 476176 251050 476232
rect 252466 476176 252522 476232
rect 241794 445848 241850 445904
rect 216586 308352 216642 308408
rect 215666 3440 215722 3496
rect 217230 195880 217286 195936
rect 217138 192752 217194 192808
rect 217322 168000 217378 168056
rect 217690 196832 217746 196888
rect 217598 193704 217654 193760
rect 217506 169904 217562 169960
rect 217782 168272 217838 168328
rect 218426 243480 218482 243536
rect 218518 189896 218574 189952
rect 218702 190984 218758 191040
rect 218610 188128 218666 188184
rect 218886 158208 218942 158264
rect 225694 310528 225750 310584
rect 227074 309576 227130 309632
rect 234618 444624 234674 444680
rect 233974 443400 234030 443456
rect 232686 443128 232742 443184
rect 233330 442992 233386 443048
rect 237838 445712 237894 445768
rect 236550 444352 236606 444408
rect 238574 444488 238630 444544
rect 239862 443264 239918 443320
rect 253846 476176 253902 476232
rect 255226 476176 255282 476232
rect 256514 476176 256570 476232
rect 259366 476720 259422 476776
rect 264794 476720 264850 476776
rect 257986 476176 258042 476232
rect 259274 476176 259330 476232
rect 262126 476448 262182 476504
rect 260746 476312 260802 476368
rect 260654 476176 260710 476232
rect 262034 476176 262090 476232
rect 263506 476176 263562 476232
rect 266266 476584 266322 476640
rect 267646 476312 267702 476368
rect 264886 476176 264942 476232
rect 266174 476176 266230 476232
rect 267554 476176 267610 476232
rect 268934 476312 268990 476368
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476604 271842 476640
rect 271786 476584 271788 476604
rect 271788 476584 271840 476604
rect 271840 476584 271842 476604
rect 274454 476448 274510 476504
rect 271694 476176 271750 476232
rect 273166 476176 273222 476232
rect 274362 476176 274418 476232
rect 274546 476312 274602 476368
rect 277306 476312 277362 476368
rect 278594 476312 278650 476368
rect 275926 476176 275982 476232
rect 277214 476176 277270 476232
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 281446 476176 281502 476232
rect 279974 443400 280030 443456
rect 284206 476176 284262 476232
rect 286506 476176 286562 476232
rect 288346 476176 288402 476232
rect 291106 476176 291162 476232
rect 293866 476176 293922 476232
rect 296626 476176 296682 476232
rect 299386 476176 299442 476232
rect 302146 476176 302202 476232
rect 303526 476176 303582 476232
rect 306286 476176 306342 476232
rect 299386 444760 299442 444816
rect 298098 441632 298154 441688
rect 300858 443264 300914 443320
rect 309046 476720 309102 476776
rect 311806 476312 311862 476368
rect 314566 476720 314622 476776
rect 315946 476196 316002 476232
rect 315946 476176 315948 476196
rect 315948 476176 316000 476196
rect 316000 476176 316002 476196
rect 318706 476468 318762 476504
rect 318706 476448 318708 476468
rect 318708 476448 318760 476468
rect 318760 476448 318762 476468
rect 321466 476176 321522 476232
rect 324226 476176 324282 476232
rect 326986 476448 327042 476504
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580262 630808 580318 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 283562 441088 283618 441144
rect 283102 440988 283104 441008
rect 283104 440988 283156 441008
rect 283156 440988 283158 441008
rect 283102 440952 283158 440988
rect 304998 441088 305054 441144
rect 298650 440952 298706 441008
rect 228638 308760 228694 308816
rect 231122 309848 231178 309904
rect 231306 309032 231362 309088
rect 232318 310664 232374 310720
rect 232962 310392 233018 310448
rect 234434 310528 234490 310584
rect 235814 310528 235870 310584
rect 234342 299240 234398 299296
rect 238022 308488 238078 308544
rect 237654 298016 237710 298072
rect 239034 301552 239090 301608
rect 241242 309440 241298 309496
rect 243358 308624 243414 308680
rect 244646 309848 244702 309904
rect 244278 308896 244334 308952
rect 245842 300736 245898 300792
rect 246394 309304 246450 309360
rect 246578 308760 246634 308816
rect 247314 309712 247370 309768
rect 248326 309032 248382 309088
rect 249062 309576 249118 309632
rect 248510 301144 248566 301200
rect 250626 309168 250682 309224
rect 249890 299376 249946 299432
rect 252650 308216 252706 308272
rect 258538 300056 258594 300112
rect 260194 302912 260250 302968
rect 263966 306448 264022 306504
rect 263782 306176 263838 306232
rect 278594 300192 278650 300248
rect 279330 300328 279386 300384
rect 282182 302776 282238 302832
rect 282550 306176 282606 306232
rect 283654 306176 283710 306232
rect 285954 284824 286010 284880
rect 287058 303184 287114 303240
rect 286138 269728 286194 269784
rect 287426 301688 287482 301744
rect 287150 254496 287206 254552
rect 288346 306040 288402 306096
rect 288898 305904 288954 305960
rect 288714 303048 288770 303104
rect 290094 305768 290150 305824
rect 291198 305632 291254 305688
rect 290186 297472 290242 297528
rect 292946 301416 293002 301472
rect 291658 297608 291714 297664
rect 291566 297336 291622 297392
rect 287518 250416 287574 250472
rect 298466 308352 298522 308408
rect 218058 3576 218114 3632
rect 216862 3440 216918 3496
rect 298282 303320 298338 303376
rect 299386 305904 299442 305960
rect 300030 300056 300086 300112
rect 303802 250552 303858 250608
rect 306102 308488 306158 308544
rect 305550 250688 305606 250744
rect 305274 247968 305330 248024
rect 306562 247560 306618 247616
rect 306470 245384 306526 245440
rect 308310 250416 308366 250472
rect 308034 247696 308090 247752
rect 309230 247832 309286 247888
rect 309322 245520 309378 245576
rect 309138 245248 309194 245304
rect 305182 245112 305238 245168
rect 304998 244976 305054 245032
rect 303710 244840 303766 244896
rect 310794 251776 310850 251832
rect 311254 260208 311310 260264
rect 311070 260072 311126 260128
rect 310978 254496 311034 254552
rect 310886 250960 310942 251016
rect 310702 250824 310758 250880
rect 312450 306040 312506 306096
rect 312358 303456 312414 303512
rect 312082 280744 312138 280800
rect 313370 265512 313426 265568
rect 317878 303184 317934 303240
rect 310610 248104 310666 248160
rect 329930 308352 329986 308408
rect 330758 305768 330814 305824
rect 331862 303048 331918 303104
rect 337290 302912 337346 302968
rect 339958 302776 340014 302832
rect 345478 305632 345534 305688
rect 346766 309032 346822 309088
rect 346950 308896 347006 308952
rect 347502 308760 347558 308816
rect 348422 308624 348478 308680
rect 349250 306312 349306 306368
rect 349986 306176 350042 306232
rect 350630 305496 350686 305552
rect 310518 244704 310574 244760
rect 298098 243480 298154 243536
rect 278134 159840 278190 159896
rect 271050 159568 271106 159624
rect 275834 159568 275890 159624
rect 220818 158616 220874 158672
rect 238114 158652 238116 158672
rect 238116 158652 238168 158672
rect 238168 158652 238170 158672
rect 219438 157800 219494 157856
rect 238114 158616 238170 158652
rect 239586 158616 239642 158672
rect 240690 158616 240746 158672
rect 248326 158616 248382 158672
rect 250442 158616 250498 158672
rect 252374 158616 252430 158672
rect 254950 158616 255006 158672
rect 255870 158616 255926 158672
rect 224958 158480 225014 158536
rect 223578 158344 223634 158400
rect 219254 3440 219310 3496
rect 227718 158208 227774 158264
rect 231858 158072 231914 158128
rect 238758 157936 238814 157992
rect 246854 158072 246910 158128
rect 246854 155896 246910 155952
rect 248694 157936 248750 157992
rect 252282 157936 252338 157992
rect 251270 155488 251326 155544
rect 253570 157936 253626 157992
rect 253662 157392 253718 157448
rect 256238 157392 256294 157448
rect 257250 158616 257306 158672
rect 259090 158616 259146 158672
rect 259550 158616 259606 158672
rect 261482 158616 261538 158672
rect 262862 158616 262918 158672
rect 263598 158616 263654 158672
rect 260654 157936 260710 157992
rect 261758 157800 261814 157856
rect 268750 158616 268806 158672
rect 269854 158616 269910 158672
rect 267646 158208 267702 158264
rect 264518 157800 264574 157856
rect 266910 157800 266966 157856
rect 265990 157664 266046 157720
rect 268934 157800 268990 157856
rect 300950 159704 301006 159760
rect 279238 159568 279294 159624
rect 288346 159568 288402 159624
rect 295890 159568 295946 159624
rect 271142 158616 271198 158672
rect 272246 158616 272302 158672
rect 274454 158616 274510 158672
rect 277030 158616 277086 158672
rect 298558 158652 298560 158672
rect 298560 158652 298612 158672
rect 298612 158652 298614 158672
rect 298558 158616 298614 158652
rect 303526 158616 303582 158672
rect 306102 158652 306104 158672
rect 306104 158652 306156 158672
rect 306156 158652 306158 158672
rect 306102 158616 306158 158652
rect 308770 158636 308826 158672
rect 308770 158616 308772 158636
rect 308772 158616 308824 158636
rect 308824 158616 308826 158636
rect 274454 158344 274510 158400
rect 276110 158344 276166 158400
rect 281354 158344 281410 158400
rect 286322 158344 286378 158400
rect 293682 158344 293738 158400
rect 274546 157664 274602 157720
rect 269118 155352 269174 155408
rect 270498 155216 270554 155272
rect 278686 157664 278742 157720
rect 283930 157528 283986 157584
rect 291014 157528 291070 157584
rect 313462 158616 313518 158672
rect 315854 158616 315910 158672
rect 318614 158616 318670 158672
rect 311070 158208 311126 158264
rect 299478 157936 299534 157992
rect 292578 153720 292634 153776
rect 290186 3304 290242 3360
rect 321006 158616 321062 158672
rect 323398 158616 323454 158672
rect 325974 158616 326030 158672
rect 354126 158208 354182 158264
rect 353942 158072 353998 158128
rect 352562 156848 352618 156904
rect 348422 156712 348478 156768
rect 345662 156576 345718 156632
rect 320914 6160 320970 6216
rect 326802 6432 326858 6488
rect 323306 6296 323362 6352
rect 325606 3576 325662 3632
rect 324410 3440 324466 3496
rect 327998 3712 328054 3768
rect 331586 3848 331642 3904
rect 335082 3984 335138 4040
rect 339866 3168 339922 3224
rect 348054 6568 348110 6624
rect 351642 6704 351698 6760
rect 357438 303320 357494 303376
rect 356886 243480 356942 243536
rect 357346 159568 357402 159624
rect 357346 158888 357402 158944
rect 356794 156848 356850 156904
rect 355966 3712 356022 3768
rect 356334 3576 356390 3632
rect 355966 3168 356022 3224
rect 358358 306448 358414 306504
rect 357622 304272 357678 304328
rect 358266 305904 358322 305960
rect 358266 160112 358322 160168
rect 358358 158888 358414 158944
rect 359646 243616 359702 243672
rect 359646 156576 359702 156632
rect 362130 309032 362186 309088
rect 361578 6704 361634 6760
rect 358726 3440 358782 3496
rect 359922 3440 359978 3496
rect 361118 3440 361174 3496
rect 364982 308896 365038 308952
rect 364890 308760 364946 308816
rect 362130 159568 362186 159624
rect 362498 158888 362554 158944
rect 362406 156712 362462 156768
rect 362314 3440 362370 3496
rect 363878 160112 363934 160168
rect 363694 157936 363750 157992
rect 363786 157392 363842 157448
rect 363510 3440 363566 3496
rect 364982 158888 365038 158944
rect 364890 158752 364946 158808
rect 365166 158208 365222 158264
rect 367006 3576 367062 3632
rect 364614 3440 364670 3496
rect 365810 3440 365866 3496
rect 370134 308624 370190 308680
rect 367650 157120 367706 157176
rect 367926 159160 367982 159216
rect 368662 306312 368718 306368
rect 368662 155896 368718 155952
rect 368846 305496 368902 305552
rect 369214 158072 369270 158128
rect 370318 306176 370374 306232
rect 370134 157256 370190 157312
rect 370318 156984 370374 157040
rect 370594 159296 370650 159352
rect 368202 3440 368258 3496
rect 369398 3440 369454 3496
rect 370594 3440 370650 3496
rect 374366 159432 374422 159488
rect 374274 158480 374330 158536
rect 577502 443128 577558 443184
rect 379978 3304 380034 3360
rect 462962 308352 463018 308408
rect 396722 303184 396778 303240
rect 476762 305768 476818 305824
rect 489182 303048 489238 303104
rect 520922 302912 520978 302968
rect 539690 302776 539746 302832
rect 570602 305632 570658 305688
rect 580354 442992 580410 443048
rect 579802 431568 579858 431624
rect 579986 418240 580042 418296
rect 579802 404912 579858 404968
rect 580078 378392 580134 378448
rect 580078 365064 580134 365120
rect 579986 351872 580042 351928
rect 580078 325216 580134 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 578882 245520 578938 245576
rect 579618 205672 579674 205728
rect 580170 165824 580226 165880
rect 580170 59608 580226 59664
rect 580906 232328 580962 232384
rect 580814 219000 580870 219056
rect 580814 192480 580870 192536
rect 580722 152632 580778 152688
rect 580630 139304 580686 139360
rect 580538 112784 580594 112840
rect 580446 72936 580502 72992
rect 580354 33088 580410 33144
rect 580262 19760 580318 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 217593 516898 217659 516901
rect 219390 516898 220064 516924
rect 217593 516896 220064 516898
rect 217593 516840 217598 516896
rect 217654 516864 220064 516896
rect 217654 516840 219450 516864
rect 217593 516838 219450 516840
rect 217593 516835 217659 516838
rect 217685 515946 217751 515949
rect 219390 515946 220064 515972
rect 217685 515944 220064 515946
rect 217685 515888 217690 515944
rect 217746 515912 220064 515944
rect 217746 515888 219450 515912
rect 217685 515886 219450 515888
rect 217685 515883 217751 515886
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 217501 513770 217567 513773
rect 219390 513770 220064 513796
rect 217501 513768 220064 513770
rect 217501 513712 217506 513768
rect 217562 513736 220064 513768
rect 217562 513712 219450 513736
rect 217501 513710 219450 513712
rect 217501 513707 217567 513710
rect 219157 512818 219223 512821
rect 219390 512818 220064 512844
rect 219157 512816 220064 512818
rect 219157 512760 219162 512816
rect 219218 512784 220064 512816
rect 219218 512760 219450 512784
rect 219157 512758 219450 512760
rect 219157 512755 219223 512758
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 219249 511050 219315 511053
rect 219390 511050 220064 511076
rect 219249 511048 220064 511050
rect 219249 510992 219254 511048
rect 219310 511016 220064 511048
rect 219310 510992 219450 511016
rect 219249 510990 219450 510992
rect 219249 510987 219315 510990
rect 219065 509962 219131 509965
rect 219390 509962 220064 509988
rect 219065 509960 220064 509962
rect 219065 509904 219070 509960
rect 219126 509928 220064 509960
rect 219126 509904 219450 509928
rect 219065 509902 219450 509904
rect 219065 509899 219131 509902
rect 218973 508194 219039 508197
rect 219390 508194 220064 508220
rect 218973 508192 220064 508194
rect 218973 508136 218978 508192
rect 219034 508160 220064 508192
rect 219034 508136 219450 508160
rect 218973 508134 219450 508136
rect 218973 508131 219039 508134
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 217409 489970 217475 489973
rect 219390 489970 220064 489996
rect 217409 489968 220064 489970
rect 217409 489912 217414 489968
rect 217470 489936 220064 489968
rect 217470 489912 219450 489936
rect 217409 489910 219450 489912
rect 217409 489907 217475 489910
rect -960 488596 480 488836
rect 218881 488338 218947 488341
rect 219390 488338 220064 488364
rect 218881 488336 220064 488338
rect 218881 488280 218886 488336
rect 218942 488304 220064 488336
rect 218942 488280 219450 488304
rect 218881 488278 219450 488280
rect 218881 488275 218947 488278
rect 217317 488066 217383 488069
rect 219390 488066 220064 488092
rect 217317 488064 220064 488066
rect 217317 488008 217322 488064
rect 217378 488032 220064 488064
rect 217378 488008 219450 488032
rect 217317 488006 219450 488008
rect 217317 488003 217383 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 238334 477260 238340 477324
rect 238404 477322 238410 477324
rect 238477 477322 238543 477325
rect 238404 477320 238543 477322
rect 238404 477264 238482 477320
rect 238538 477264 238543 477320
rect 238404 477262 238543 477264
rect 238404 477260 238410 477262
rect 238477 477259 238543 477262
rect 241830 477124 241836 477188
rect 241900 477186 241906 477188
rect 242801 477186 242867 477189
rect 241900 477184 242867 477186
rect 241900 477128 242806 477184
rect 242862 477128 242867 477184
rect 241900 477126 242867 477128
rect 241900 477124 241906 477126
rect 242801 477123 242867 477126
rect 256182 476988 256188 477052
rect 256252 477050 256258 477052
rect 256601 477050 256667 477053
rect 256252 477048 256667 477050
rect 256252 476992 256606 477048
rect 256662 476992 256667 477048
rect 256252 476990 256667 476992
rect 256252 476988 256258 476990
rect 256601 476987 256667 476990
rect 239622 476852 239628 476916
rect 239692 476914 239698 476916
rect 240041 476914 240107 476917
rect 239692 476912 240107 476914
rect 239692 476856 240046 476912
rect 240102 476856 240107 476912
rect 239692 476854 240107 476856
rect 239692 476852 239698 476854
rect 240041 476851 240107 476854
rect 240542 476852 240548 476916
rect 240612 476914 240618 476916
rect 241421 476914 241487 476917
rect 240612 476912 241487 476914
rect 240612 476856 241426 476912
rect 241482 476856 241487 476912
rect 240612 476854 241487 476856
rect 240612 476852 240618 476854
rect 241421 476851 241487 476854
rect 236126 476716 236132 476780
rect 236196 476778 236202 476780
rect 237281 476778 237347 476781
rect 236196 476776 237347 476778
rect 236196 476720 237286 476776
rect 237342 476720 237347 476776
rect 236196 476718 237347 476720
rect 236196 476716 236202 476718
rect 237281 476715 237347 476718
rect 258022 476716 258028 476780
rect 258092 476778 258098 476780
rect 259361 476778 259427 476781
rect 258092 476776 259427 476778
rect 258092 476720 259366 476776
rect 259422 476720 259427 476776
rect 258092 476718 259427 476720
rect 258092 476716 258098 476718
rect 259361 476715 259427 476718
rect 263542 476716 263548 476780
rect 263612 476778 263618 476780
rect 264789 476778 264855 476781
rect 263612 476776 264855 476778
rect 263612 476720 264794 476776
rect 264850 476720 264855 476776
rect 263612 476718 264855 476720
rect 263612 476716 263618 476718
rect 264789 476715 264855 476718
rect 308622 476716 308628 476780
rect 308692 476778 308698 476780
rect 309041 476778 309107 476781
rect 308692 476776 309107 476778
rect 308692 476720 309046 476776
rect 309102 476720 309107 476776
rect 308692 476718 309107 476720
rect 308692 476716 308698 476718
rect 309041 476715 309107 476718
rect 313406 476716 313412 476780
rect 313476 476778 313482 476780
rect 314561 476778 314627 476781
rect 313476 476776 314627 476778
rect 313476 476720 314566 476776
rect 314622 476720 314627 476776
rect 313476 476718 314627 476720
rect 313476 476716 313482 476718
rect 314561 476715 314627 476718
rect 265934 476580 265940 476644
rect 266004 476642 266010 476644
rect 266261 476642 266327 476645
rect 266004 476640 266327 476642
rect 266004 476584 266266 476640
rect 266322 476584 266327 476640
rect 266004 476582 266327 476584
rect 266004 476580 266010 476582
rect 266261 476579 266327 476582
rect 270902 476580 270908 476644
rect 270972 476642 270978 476644
rect 271781 476642 271847 476645
rect 270972 476640 271847 476642
rect 270972 476584 271786 476640
rect 271842 476584 271847 476640
rect 270972 476582 271847 476584
rect 270972 476580 270978 476582
rect 271781 476579 271847 476582
rect 253422 476444 253428 476508
rect 253492 476506 253498 476508
rect 253749 476506 253815 476509
rect 253492 476504 253815 476506
rect 253492 476448 253754 476504
rect 253810 476448 253815 476504
rect 253492 476446 253815 476448
rect 253492 476444 253498 476446
rect 253749 476443 253815 476446
rect 261150 476444 261156 476508
rect 261220 476506 261226 476508
rect 262121 476506 262187 476509
rect 274449 476508 274515 476509
rect 261220 476504 262187 476506
rect 261220 476448 262126 476504
rect 262182 476448 262187 476504
rect 261220 476446 262187 476448
rect 261220 476444 261226 476446
rect 262121 476443 262187 476446
rect 274398 476444 274404 476508
rect 274468 476506 274515 476508
rect 274468 476504 274560 476506
rect 274510 476448 274560 476504
rect 274468 476446 274560 476448
rect 274468 476444 274515 476446
rect 318558 476444 318564 476508
rect 318628 476506 318634 476508
rect 318701 476506 318767 476509
rect 318628 476504 318767 476506
rect 318628 476448 318706 476504
rect 318762 476448 318767 476504
rect 318628 476446 318767 476448
rect 318628 476444 318634 476446
rect 274449 476443 274515 476444
rect 318701 476443 318767 476446
rect 325918 476444 325924 476508
rect 325988 476506 325994 476508
rect 326981 476506 327047 476509
rect 325988 476504 327047 476506
rect 325988 476448 326986 476504
rect 327042 476448 327047 476504
rect 325988 476446 327047 476448
rect 325988 476444 325994 476446
rect 326981 476443 327047 476446
rect 244222 476308 244228 476372
rect 244292 476370 244298 476372
rect 245469 476370 245535 476373
rect 244292 476368 245535 476370
rect 244292 476312 245474 476368
rect 245530 476312 245535 476368
rect 244292 476310 245535 476312
rect 244292 476308 244298 476310
rect 245469 476307 245535 476310
rect 247718 476308 247724 476372
rect 247788 476370 247794 476372
rect 248321 476370 248387 476373
rect 247788 476368 248387 476370
rect 247788 476312 248326 476368
rect 248382 476312 248387 476368
rect 247788 476310 248387 476312
rect 247788 476308 247794 476310
rect 248321 476307 248387 476310
rect 250110 476308 250116 476372
rect 250180 476370 250186 476372
rect 251081 476370 251147 476373
rect 250180 476368 251147 476370
rect 250180 476312 251086 476368
rect 251142 476312 251147 476368
rect 250180 476310 251147 476312
rect 250180 476308 250186 476310
rect 251081 476307 251147 476310
rect 251398 476308 251404 476372
rect 251468 476370 251474 476372
rect 252369 476370 252435 476373
rect 251468 476368 252435 476370
rect 251468 476312 252374 476368
rect 252430 476312 252435 476368
rect 251468 476310 252435 476312
rect 251468 476308 251474 476310
rect 252369 476307 252435 476310
rect 259494 476308 259500 476372
rect 259564 476370 259570 476372
rect 260741 476370 260807 476373
rect 259564 476368 260807 476370
rect 259564 476312 260746 476368
rect 260802 476312 260807 476368
rect 259564 476310 260807 476312
rect 259564 476308 259570 476310
rect 260741 476307 260807 476310
rect 266486 476308 266492 476372
rect 266556 476370 266562 476372
rect 267641 476370 267707 476373
rect 266556 476368 267707 476370
rect 266556 476312 267646 476368
rect 267702 476312 267707 476368
rect 266556 476310 267707 476312
rect 266556 476308 266562 476310
rect 267641 476307 267707 476310
rect 268326 476308 268332 476372
rect 268396 476370 268402 476372
rect 268929 476370 268995 476373
rect 268396 476368 268995 476370
rect 268396 476312 268934 476368
rect 268990 476312 268995 476368
rect 268396 476310 268995 476312
rect 268396 476308 268402 476310
rect 268929 476307 268995 476310
rect 273662 476308 273668 476372
rect 273732 476370 273738 476372
rect 274541 476370 274607 476373
rect 273732 476368 274607 476370
rect 273732 476312 274546 476368
rect 274602 476312 274607 476368
rect 273732 476310 274607 476312
rect 273732 476308 273738 476310
rect 274541 476307 274607 476310
rect 276054 476308 276060 476372
rect 276124 476370 276130 476372
rect 277301 476370 277367 476373
rect 276124 476368 277367 476370
rect 276124 476312 277306 476368
rect 277362 476312 277367 476368
rect 276124 476310 277367 476312
rect 276124 476308 276130 476310
rect 277301 476307 277367 476310
rect 278078 476308 278084 476372
rect 278148 476370 278154 476372
rect 278589 476370 278655 476373
rect 278148 476368 278655 476370
rect 278148 476312 278594 476368
rect 278650 476312 278655 476368
rect 278148 476310 278655 476312
rect 278148 476308 278154 476310
rect 278589 476307 278655 476310
rect 311014 476308 311020 476372
rect 311084 476370 311090 476372
rect 311801 476370 311867 476373
rect 311084 476368 311867 476370
rect 311084 476312 311806 476368
rect 311862 476312 311867 476368
rect 311084 476310 311867 476312
rect 311084 476308 311090 476310
rect 311801 476307 311867 476310
rect 237189 476236 237255 476237
rect 237189 476234 237236 476236
rect 237144 476232 237236 476234
rect 237144 476176 237194 476232
rect 237144 476174 237236 476176
rect 237189 476172 237236 476174
rect 237300 476172 237306 476236
rect 243118 476172 243124 476236
rect 243188 476234 243194 476236
rect 244181 476234 244247 476237
rect 245561 476236 245627 476237
rect 243188 476232 244247 476234
rect 243188 476176 244186 476232
rect 244242 476176 244247 476232
rect 243188 476174 244247 476176
rect 243188 476172 243194 476174
rect 237189 476171 237255 476172
rect 244181 476171 244247 476174
rect 245510 476172 245516 476236
rect 245580 476234 245627 476236
rect 245580 476232 245672 476234
rect 245622 476176 245672 476232
rect 245580 476174 245672 476176
rect 245580 476172 245627 476174
rect 246614 476172 246620 476236
rect 246684 476234 246690 476236
rect 246941 476234 247007 476237
rect 248229 476236 248295 476237
rect 248229 476234 248276 476236
rect 246684 476232 247007 476234
rect 246684 476176 246946 476232
rect 247002 476176 247007 476232
rect 246684 476174 247007 476176
rect 248184 476232 248276 476234
rect 248184 476176 248234 476232
rect 248184 476174 248276 476176
rect 246684 476172 246690 476174
rect 245561 476171 245627 476172
rect 246941 476171 247007 476174
rect 248229 476172 248276 476174
rect 248340 476172 248346 476236
rect 248638 476172 248644 476236
rect 248708 476234 248714 476236
rect 249701 476234 249767 476237
rect 248708 476232 249767 476234
rect 248708 476176 249706 476232
rect 249762 476176 249767 476232
rect 248708 476174 249767 476176
rect 248708 476172 248714 476174
rect 248229 476171 248295 476172
rect 249701 476171 249767 476174
rect 250846 476172 250852 476236
rect 250916 476234 250922 476236
rect 250989 476234 251055 476237
rect 250916 476232 251055 476234
rect 250916 476176 250994 476232
rect 251050 476176 251055 476232
rect 250916 476174 251055 476176
rect 250916 476172 250922 476174
rect 250989 476171 251055 476174
rect 252318 476172 252324 476236
rect 252388 476234 252394 476236
rect 252461 476234 252527 476237
rect 252388 476232 252527 476234
rect 252388 476176 252466 476232
rect 252522 476176 252527 476232
rect 252388 476174 252527 476176
rect 252388 476172 252394 476174
rect 252461 476171 252527 476174
rect 253606 476172 253612 476236
rect 253676 476234 253682 476236
rect 253841 476234 253907 476237
rect 253676 476232 253907 476234
rect 253676 476176 253846 476232
rect 253902 476176 253907 476232
rect 253676 476174 253907 476176
rect 253676 476172 253682 476174
rect 253841 476171 253907 476174
rect 254526 476172 254532 476236
rect 254596 476234 254602 476236
rect 255221 476234 255287 476237
rect 254596 476232 255287 476234
rect 254596 476176 255226 476232
rect 255282 476176 255287 476232
rect 254596 476174 255287 476176
rect 254596 476172 254602 476174
rect 255221 476171 255287 476174
rect 255814 476172 255820 476236
rect 255884 476234 255890 476236
rect 256509 476234 256575 476237
rect 255884 476232 256575 476234
rect 255884 476176 256514 476232
rect 256570 476176 256575 476232
rect 255884 476174 256575 476176
rect 255884 476172 255890 476174
rect 256509 476171 256575 476174
rect 257102 476172 257108 476236
rect 257172 476234 257178 476236
rect 257981 476234 258047 476237
rect 257172 476232 258047 476234
rect 257172 476176 257986 476232
rect 258042 476176 258047 476232
rect 257172 476174 258047 476176
rect 257172 476172 257178 476174
rect 257981 476171 258047 476174
rect 258574 476172 258580 476236
rect 258644 476234 258650 476236
rect 259269 476234 259335 476237
rect 260649 476236 260715 476237
rect 258644 476232 259335 476234
rect 258644 476176 259274 476232
rect 259330 476176 259335 476232
rect 258644 476174 259335 476176
rect 258644 476172 258650 476174
rect 259269 476171 259335 476174
rect 260598 476172 260604 476236
rect 260668 476234 260715 476236
rect 260668 476232 260760 476234
rect 260710 476176 260760 476232
rect 260668 476174 260760 476176
rect 260668 476172 260715 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262029 476234 262095 476237
rect 261772 476232 262095 476234
rect 261772 476176 262034 476232
rect 262090 476176 262095 476232
rect 261772 476174 262095 476176
rect 261772 476172 261778 476174
rect 260649 476171 260715 476172
rect 262029 476171 262095 476174
rect 262806 476172 262812 476236
rect 262876 476234 262882 476236
rect 263501 476234 263567 476237
rect 262876 476232 263567 476234
rect 262876 476176 263506 476232
rect 263562 476176 263567 476232
rect 262876 476174 263567 476176
rect 262876 476172 262882 476174
rect 263501 476171 263567 476174
rect 263910 476172 263916 476236
rect 263980 476234 263986 476236
rect 264881 476234 264947 476237
rect 263980 476232 264947 476234
rect 263980 476176 264886 476232
rect 264942 476176 264947 476232
rect 263980 476174 264947 476176
rect 263980 476172 263986 476174
rect 264881 476171 264947 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266169 476234 266235 476237
rect 267549 476236 267615 476237
rect 267549 476234 267596 476236
rect 265452 476232 266235 476234
rect 265452 476176 266174 476232
rect 266230 476176 266235 476232
rect 265452 476174 266235 476176
rect 267504 476232 267596 476234
rect 267504 476176 267554 476232
rect 267504 476174 267596 476176
rect 265452 476172 265458 476174
rect 266169 476171 266235 476174
rect 267549 476172 267596 476174
rect 267660 476172 267666 476236
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 267549 476171 267615 476172
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271689 476234 271755 476237
rect 271340 476232 271755 476234
rect 271340 476176 271694 476232
rect 271750 476176 271755 476232
rect 271340 476174 271755 476176
rect 271340 476172 271346 476174
rect 271689 476171 271755 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 273294 476172 273300 476236
rect 273364 476234 273370 476236
rect 274357 476234 274423 476237
rect 275921 476236 275987 476237
rect 273364 476232 274423 476234
rect 273364 476176 274362 476232
rect 274418 476176 274423 476232
rect 273364 476174 274423 476176
rect 273364 476172 273370 476174
rect 274357 476171 274423 476174
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277209 476234 277275 476237
rect 277044 476232 277275 476234
rect 277044 476176 277214 476232
rect 277270 476176 277275 476232
rect 277044 476174 277275 476176
rect 277044 476172 277050 476174
rect 275921 476171 275987 476172
rect 277209 476171 277275 476174
rect 278446 476172 278452 476236
rect 278516 476234 278522 476236
rect 278681 476234 278747 476237
rect 278516 476232 278747 476234
rect 278516 476176 278686 476232
rect 278742 476176 278747 476232
rect 278516 476174 278747 476176
rect 278516 476172 278522 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 281022 476172 281028 476236
rect 281092 476234 281098 476236
rect 281441 476234 281507 476237
rect 281092 476232 281507 476234
rect 281092 476176 281446 476232
rect 281502 476176 281507 476232
rect 281092 476174 281507 476176
rect 281092 476172 281098 476174
rect 281441 476171 281507 476174
rect 283598 476172 283604 476236
rect 283668 476234 283674 476236
rect 284201 476234 284267 476237
rect 283668 476232 284267 476234
rect 283668 476176 284206 476232
rect 284262 476176 284267 476232
rect 283668 476174 284267 476176
rect 283668 476172 283674 476174
rect 284201 476171 284267 476174
rect 285990 476172 285996 476236
rect 286060 476234 286066 476236
rect 286501 476234 286567 476237
rect 286060 476232 286567 476234
rect 286060 476176 286506 476232
rect 286562 476176 286567 476232
rect 286060 476174 286567 476176
rect 286060 476172 286066 476174
rect 286501 476171 286567 476174
rect 288198 476172 288204 476236
rect 288268 476234 288274 476236
rect 288341 476234 288407 476237
rect 288268 476232 288407 476234
rect 288268 476176 288346 476232
rect 288402 476176 288407 476232
rect 288268 476174 288407 476176
rect 288268 476172 288274 476174
rect 288341 476171 288407 476174
rect 290958 476172 290964 476236
rect 291028 476234 291034 476236
rect 291101 476234 291167 476237
rect 291028 476232 291167 476234
rect 291028 476176 291106 476232
rect 291162 476176 291167 476232
rect 291028 476174 291167 476176
rect 291028 476172 291034 476174
rect 291101 476171 291167 476174
rect 293534 476172 293540 476236
rect 293604 476234 293610 476236
rect 293861 476234 293927 476237
rect 293604 476232 293927 476234
rect 293604 476176 293866 476232
rect 293922 476176 293927 476232
rect 293604 476174 293927 476176
rect 293604 476172 293610 476174
rect 293861 476171 293927 476174
rect 295926 476172 295932 476236
rect 295996 476234 296002 476236
rect 296621 476234 296687 476237
rect 295996 476232 296687 476234
rect 295996 476176 296626 476232
rect 296682 476176 296687 476232
rect 295996 476174 296687 476176
rect 295996 476172 296002 476174
rect 296621 476171 296687 476174
rect 298502 476172 298508 476236
rect 298572 476234 298578 476236
rect 299381 476234 299447 476237
rect 298572 476232 299447 476234
rect 298572 476176 299386 476232
rect 299442 476176 299447 476232
rect 298572 476174 299447 476176
rect 298572 476172 298578 476174
rect 299381 476171 299447 476174
rect 300894 476172 300900 476236
rect 300964 476234 300970 476236
rect 302141 476234 302207 476237
rect 303521 476236 303587 476237
rect 300964 476232 302207 476234
rect 300964 476176 302146 476232
rect 302202 476176 302207 476232
rect 300964 476174 302207 476176
rect 300964 476172 300970 476174
rect 302141 476171 302207 476174
rect 303470 476172 303476 476236
rect 303540 476234 303587 476236
rect 303540 476232 303632 476234
rect 303582 476176 303632 476232
rect 303540 476174 303632 476176
rect 303540 476172 303587 476174
rect 306046 476172 306052 476236
rect 306116 476234 306122 476236
rect 306281 476234 306347 476237
rect 306116 476232 306347 476234
rect 306116 476176 306286 476232
rect 306342 476176 306347 476232
rect 306116 476174 306347 476176
rect 306116 476172 306122 476174
rect 303521 476171 303587 476172
rect 306281 476171 306347 476174
rect 315798 476172 315804 476236
rect 315868 476234 315874 476236
rect 315941 476234 316007 476237
rect 315868 476232 316007 476234
rect 315868 476176 315946 476232
rect 316002 476176 316007 476232
rect 315868 476174 316007 476176
rect 315868 476172 315874 476174
rect 315941 476171 316007 476174
rect 320950 476172 320956 476236
rect 321020 476234 321026 476236
rect 321461 476234 321527 476237
rect 321020 476232 321527 476234
rect 321020 476176 321466 476232
rect 321522 476176 321527 476232
rect 321020 476174 321527 476176
rect 321020 476172 321026 476174
rect 321461 476171 321527 476174
rect 323342 476172 323348 476236
rect 323412 476234 323418 476236
rect 324221 476234 324287 476237
rect 323412 476232 324287 476234
rect 323412 476176 324226 476232
rect 324282 476176 324287 476232
rect 323412 476174 324287 476176
rect 323412 476172 323418 476174
rect 324221 476171 324287 476174
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 4061 449578 4127 449581
rect -960 449576 4127 449578
rect -960 449520 4066 449576
rect 4122 449520 4127 449576
rect -960 449518 4127 449520
rect -960 449428 480 449518
rect 4061 449515 4127 449518
rect 241789 445906 241855 445909
rect 367870 445906 367876 445908
rect 241789 445904 367876 445906
rect 241789 445848 241794 445904
rect 241850 445848 367876 445904
rect 241789 445846 367876 445848
rect 241789 445843 241855 445846
rect 367870 445844 367876 445846
rect 367940 445844 367946 445908
rect 237833 445770 237899 445773
rect 365110 445770 365116 445772
rect 237833 445768 365116 445770
rect 237833 445712 237838 445768
rect 237894 445712 365116 445768
rect 237833 445710 365116 445712
rect 237833 445707 237899 445710
rect 365110 445708 365116 445710
rect 365180 445708 365186 445772
rect 214598 444756 214604 444820
rect 214668 444818 214674 444820
rect 299381 444818 299447 444821
rect 214668 444816 299447 444818
rect 214668 444760 299386 444816
rect 299442 444760 299447 444816
rect 214668 444758 299447 444760
rect 214668 444756 214674 444758
rect 299381 444755 299447 444758
rect 234613 444682 234679 444685
rect 364926 444682 364932 444684
rect 234613 444680 364932 444682
rect 234613 444624 234618 444680
rect 234674 444624 364932 444680
rect 234613 444622 364932 444624
rect 234613 444619 234679 444622
rect 364926 444620 364932 444622
rect 364996 444620 365002 444684
rect 583520 444668 584960 444908
rect 238569 444546 238635 444549
rect 368974 444546 368980 444548
rect 238569 444544 368980 444546
rect 238569 444488 238574 444544
rect 238630 444488 368980 444544
rect 238569 444486 368980 444488
rect 238569 444483 238635 444486
rect 368974 444484 368980 444486
rect 369044 444484 369050 444548
rect 236545 444410 236611 444413
rect 367686 444410 367692 444412
rect 236545 444408 367692 444410
rect 236545 444352 236550 444408
rect 236606 444352 367692 444408
rect 236545 444350 367692 444352
rect 236545 444347 236611 444350
rect 367686 444348 367692 444350
rect 367756 444348 367762 444412
rect 233969 443458 234035 443461
rect 279969 443458 280035 443461
rect 233969 443456 280035 443458
rect 233969 443400 233974 443456
rect 234030 443400 279974 443456
rect 280030 443400 280035 443456
rect 233969 443398 280035 443400
rect 233969 443395 234035 443398
rect 279969 443395 280035 443398
rect 239857 443322 239923 443325
rect 300853 443322 300919 443325
rect 239857 443320 300919 443322
rect 239857 443264 239862 443320
rect 239918 443264 300858 443320
rect 300914 443264 300919 443320
rect 239857 443262 300919 443264
rect 239857 443259 239923 443262
rect 300853 443259 300919 443262
rect 232681 443186 232747 443189
rect 577497 443186 577563 443189
rect 232681 443184 577563 443186
rect 232681 443128 232686 443184
rect 232742 443128 577502 443184
rect 577558 443128 577563 443184
rect 232681 443126 577563 443128
rect 232681 443123 232747 443126
rect 577497 443123 577563 443126
rect 233325 443050 233391 443053
rect 580349 443050 580415 443053
rect 233325 443048 580415 443050
rect 233325 442992 233330 443048
rect 233386 442992 580354 443048
rect 580410 442992 580415 443048
rect 233325 442990 580415 442992
rect 233325 442987 233391 442990
rect 580349 442987 580415 442990
rect 216070 441628 216076 441692
rect 216140 441690 216146 441692
rect 298093 441690 298159 441693
rect 216140 441688 298159 441690
rect 216140 441632 298098 441688
rect 298154 441632 298159 441688
rect 216140 441630 298159 441632
rect 216140 441628 216146 441630
rect 298093 441627 298159 441630
rect 283557 441146 283623 441149
rect 304993 441146 305059 441149
rect 283557 441144 305059 441146
rect 283557 441088 283562 441144
rect 283618 441088 304998 441144
rect 305054 441088 305059 441144
rect 283557 441086 305059 441088
rect 283557 441083 283623 441086
rect 304993 441083 305059 441086
rect 283097 441010 283163 441013
rect 298645 441010 298711 441013
rect 283097 441008 298711 441010
rect 283097 440952 283102 441008
rect 283158 440952 298650 441008
rect 298706 440952 298711 441008
rect 283097 440950 298711 440952
rect 283097 440947 283163 440950
rect 298645 440947 298711 440950
rect -960 436508 480 436748
rect 579797 431626 579863 431629
rect 583520 431626 584960 431716
rect 579797 431624 584960 431626
rect 579797 431568 579802 431624
rect 579858 431568 584960 431624
rect 579797 431566 584960 431568
rect 579797 431563 579863 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579981 418298 580047 418301
rect 583520 418298 584960 418388
rect 579981 418296 584960 418298
rect 579981 418240 579986 418296
rect 580042 418240 584960 418296
rect 579981 418238 584960 418240
rect 579981 418235 580047 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 579797 404970 579863 404973
rect 583520 404970 584960 405060
rect 579797 404968 584960 404970
rect 579797 404912 579802 404968
rect 579858 404912 584960 404968
rect 579797 404910 584960 404912
rect 579797 404907 579863 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect 159909 374098 159975 374101
rect 232078 374098 232084 374100
rect 159909 374096 232084 374098
rect 159909 374040 159914 374096
rect 159970 374040 232084 374096
rect 159909 374038 232084 374040
rect 159909 374035 159975 374038
rect 232078 374036 232084 374038
rect 232148 374036 232154 374100
rect 134149 372738 134215 372741
rect 232078 372738 232084 372740
rect 134149 372736 232084 372738
rect 134149 372680 134154 372736
rect 134210 372680 232084 372736
rect 134149 372678 232084 372680
rect 134149 372675 134215 372678
rect 232078 372676 232084 372678
rect 232148 372676 232154 372740
rect 133873 371650 133939 371653
rect 135161 371650 135227 371653
rect 133873 371648 135227 371650
rect 133873 371592 133878 371648
rect 133934 371592 135166 371648
rect 135222 371592 135227 371648
rect 133873 371590 135227 371592
rect 133873 371587 133939 371590
rect 135161 371587 135227 371590
rect 143257 371650 143323 371653
rect 153009 371650 153075 371653
rect 143257 371648 153075 371650
rect 143257 371592 143262 371648
rect 143318 371592 153014 371648
rect 153070 371592 153075 371648
rect 143257 371590 153075 371592
rect 143257 371587 143323 371590
rect 153009 371587 153075 371590
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 99833 370698 99899 370701
rect 99833 370696 100218 370698
rect 99833 370640 99838 370696
rect 99894 370640 100218 370696
rect 99833 370638 100218 370640
rect 99833 370635 99899 370638
rect 100158 370124 100218 370638
rect 172329 369474 172395 369477
rect 169924 369472 172395 369474
rect 169924 369416 172334 369472
rect 172390 369416 172395 369472
rect 169924 369414 172395 369416
rect 172329 369411 172395 369414
rect 97901 367434 97967 367437
rect 97901 367432 100188 367434
rect 97901 367376 97906 367432
rect 97962 367376 100188 367432
rect 97901 367374 100188 367376
rect 97901 367371 97967 367374
rect 172421 366754 172487 366757
rect 169924 366752 172487 366754
rect 169924 366696 172426 366752
rect 172482 366696 172487 366752
rect 169924 366694 172487 366696
rect 172421 366691 172487 366694
rect 580073 365122 580139 365125
rect 583520 365122 584960 365212
rect 580073 365120 584960 365122
rect 580073 365064 580078 365120
rect 580134 365064 584960 365120
rect 580073 365062 584960 365064
rect 580073 365059 580139 365062
rect 583520 364972 584960 365062
rect 97809 364714 97875 364717
rect 97809 364712 100188 364714
rect 97809 364656 97814 364712
rect 97870 364656 100188 364712
rect 97809 364654 100188 364656
rect 97809 364651 97875 364654
rect 171869 364034 171935 364037
rect 169924 364032 171935 364034
rect 169924 363976 171874 364032
rect 171930 363976 171935 364032
rect 169924 363974 171935 363976
rect 171869 363971 171935 363974
rect 97717 361994 97783 361997
rect 97717 361992 100188 361994
rect 97717 361936 97722 361992
rect 97778 361936 100188 361992
rect 97717 361934 100188 361936
rect 97717 361931 97783 361934
rect 171961 361314 172027 361317
rect 169924 361312 172027 361314
rect 169924 361256 171966 361312
rect 172022 361256 172027 361312
rect 169924 361254 172027 361256
rect 171961 361251 172027 361254
rect 99281 359274 99347 359277
rect 99281 359272 100188 359274
rect 99281 359216 99286 359272
rect 99342 359216 100188 359272
rect 99281 359214 100188 359216
rect 99281 359211 99347 359214
rect 171685 358594 171751 358597
rect 169924 358592 171751 358594
rect -960 358458 480 358548
rect 169924 358536 171690 358592
rect 171746 358536 171751 358592
rect 169924 358534 171751 358536
rect 171685 358531 171751 358534
rect 3693 358458 3759 358461
rect -960 358456 3759 358458
rect -960 358400 3698 358456
rect 3754 358400 3759 358456
rect -960 358398 3759 358400
rect -960 358308 480 358398
rect 3693 358395 3759 358398
rect 99189 356554 99255 356557
rect 99189 356552 100188 356554
rect 99189 356496 99194 356552
rect 99250 356496 100188 356552
rect 99189 356494 100188 356496
rect 99189 356491 99255 356494
rect 172421 355874 172487 355877
rect 169924 355872 172487 355874
rect 169924 355816 172426 355872
rect 172482 355816 172487 355872
rect 169924 355814 172487 355816
rect 172421 355811 172487 355814
rect 97901 353834 97967 353837
rect 97901 353832 100188 353834
rect 97901 353776 97906 353832
rect 97962 353776 100188 353832
rect 97901 353774 100188 353776
rect 97901 353771 97967 353774
rect 172421 353154 172487 353157
rect 169924 353152 172487 353154
rect 169924 353096 172426 353152
rect 172482 353096 172487 353152
rect 169924 353094 172487 353096
rect 172421 353091 172487 353094
rect 579981 351930 580047 351933
rect 583520 351930 584960 352020
rect 579981 351928 584960 351930
rect 579981 351872 579986 351928
rect 580042 351872 584960 351928
rect 579981 351870 584960 351872
rect 579981 351867 580047 351870
rect 583520 351780 584960 351870
rect 97625 351114 97691 351117
rect 97625 351112 100188 351114
rect 97625 351056 97630 351112
rect 97686 351056 100188 351112
rect 97625 351054 100188 351056
rect 97625 351051 97691 351054
rect 171869 350434 171935 350437
rect 169924 350432 171935 350434
rect 169924 350376 171874 350432
rect 171930 350376 171935 350432
rect 169924 350374 171935 350376
rect 171869 350371 171935 350374
rect 99097 348394 99163 348397
rect 99097 348392 100188 348394
rect 99097 348336 99102 348392
rect 99158 348336 100188 348392
rect 99097 348334 100188 348336
rect 99097 348331 99163 348334
rect 172421 347714 172487 347717
rect 169924 347712 172487 347714
rect 169924 347656 172426 347712
rect 172482 347656 172487 347712
rect 169924 347654 172487 347656
rect 172421 347651 172487 347654
rect 97809 345674 97875 345677
rect 97809 345672 100188 345674
rect 97809 345616 97814 345672
rect 97870 345616 100188 345672
rect 97809 345614 100188 345616
rect 97809 345611 97875 345614
rect -960 345402 480 345492
rect 3601 345402 3667 345405
rect -960 345400 3667 345402
rect -960 345344 3606 345400
rect 3662 345344 3667 345400
rect -960 345342 3667 345344
rect -960 345252 480 345342
rect 3601 345339 3667 345342
rect 172053 344994 172119 344997
rect 169924 344992 172119 344994
rect 169924 344936 172058 344992
rect 172114 344936 172119 344992
rect 169924 344934 172119 344936
rect 172053 344931 172119 344934
rect 99005 342954 99071 342957
rect 99005 342952 100188 342954
rect 99005 342896 99010 342952
rect 99066 342896 100188 342952
rect 99005 342894 100188 342896
rect 99005 342891 99071 342894
rect 172421 342274 172487 342277
rect 169924 342272 172487 342274
rect 169924 342216 172426 342272
rect 172482 342216 172487 342272
rect 169924 342214 172487 342216
rect 172421 342211 172487 342214
rect 97717 340234 97783 340237
rect 97717 340232 100188 340234
rect 97717 340176 97722 340232
rect 97778 340176 100188 340232
rect 97717 340174 100188 340176
rect 97717 340171 97783 340174
rect 172145 339554 172211 339557
rect 169924 339552 172211 339554
rect 169924 339496 172150 339552
rect 172206 339496 172211 339552
rect 169924 339494 172211 339496
rect 172145 339491 172211 339494
rect 583520 338452 584960 338692
rect 98913 337514 98979 337517
rect 98913 337512 100188 337514
rect 98913 337456 98918 337512
rect 98974 337456 100188 337512
rect 98913 337454 100188 337456
rect 98913 337451 98979 337454
rect 172421 336834 172487 336837
rect 169924 336832 172487 336834
rect 169924 336776 172426 336832
rect 172482 336776 172487 336832
rect 169924 336774 172487 336776
rect 172421 336771 172487 336774
rect 97625 334794 97691 334797
rect 97625 334792 100188 334794
rect 97625 334736 97630 334792
rect 97686 334736 100188 334792
rect 97625 334734 100188 334736
rect 97625 334731 97691 334734
rect 172421 334114 172487 334117
rect 169924 334112 172487 334114
rect 169924 334056 172426 334112
rect 172482 334056 172487 334112
rect 169924 334054 172487 334056
rect 172421 334051 172487 334054
rect -960 332196 480 332436
rect 97533 332074 97599 332077
rect 97533 332072 100188 332074
rect 97533 332016 97538 332072
rect 97594 332016 100188 332072
rect 97533 332014 100188 332016
rect 97533 332011 97599 332014
rect 172421 331394 172487 331397
rect 169924 331392 172487 331394
rect 169924 331336 172426 331392
rect 172482 331336 172487 331392
rect 169924 331334 172487 331336
rect 172421 331331 172487 331334
rect 98821 329354 98887 329357
rect 98821 329352 100188 329354
rect 98821 329296 98826 329352
rect 98882 329296 100188 329352
rect 98821 329294 100188 329296
rect 98821 329291 98887 329294
rect 172421 328674 172487 328677
rect 169924 328672 172487 328674
rect 169924 328616 172426 328672
rect 172482 328616 172487 328672
rect 169924 328614 172487 328616
rect 172421 328611 172487 328614
rect 97441 326634 97507 326637
rect 97441 326632 100188 326634
rect 97441 326576 97446 326632
rect 97502 326576 100188 326632
rect 97441 326574 100188 326576
rect 97441 326571 97507 326574
rect 171409 325954 171475 325957
rect 169924 325952 171475 325954
rect 169924 325896 171414 325952
rect 171470 325896 171475 325952
rect 169924 325894 171475 325896
rect 171409 325891 171475 325894
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect 97349 323914 97415 323917
rect 97349 323912 100188 323914
rect 97349 323856 97354 323912
rect 97410 323856 100188 323912
rect 97349 323854 100188 323856
rect 97349 323851 97415 323854
rect 172237 323234 172303 323237
rect 169924 323232 172303 323234
rect 169924 323176 172242 323232
rect 172298 323176 172303 323232
rect 169924 323174 172303 323176
rect 172237 323171 172303 323174
rect 98729 321194 98795 321197
rect 98729 321192 100188 321194
rect 98729 321136 98734 321192
rect 98790 321136 100188 321192
rect 98729 321134 100188 321136
rect 98729 321131 98795 321134
rect 172421 320514 172487 320517
rect 169924 320512 172487 320514
rect 169924 320456 172426 320512
rect 172482 320456 172487 320512
rect 169924 320454 172487 320456
rect 172421 320451 172487 320454
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 99373 318474 99439 318477
rect 99373 318472 100188 318474
rect 99373 318416 99378 318472
rect 99434 318416 100188 318472
rect 99373 318414 100188 318416
rect 99373 318411 99439 318414
rect 172421 317794 172487 317797
rect 169924 317792 172487 317794
rect 169924 317736 172426 317792
rect 172482 317736 172487 317792
rect 169924 317734 172487 317736
rect 172421 317731 172487 317734
rect 98637 315754 98703 315757
rect 98637 315752 100188 315754
rect 98637 315696 98642 315752
rect 98698 315696 100188 315752
rect 98637 315694 100188 315696
rect 98637 315691 98703 315694
rect 172421 315074 172487 315077
rect 169924 315072 172487 315074
rect 169924 315016 172426 315072
rect 172482 315016 172487 315072
rect 169924 315014 172487 315016
rect 172421 315011 172487 315014
rect 99465 313034 99531 313037
rect 99465 313032 100188 313034
rect 99465 312976 99470 313032
rect 99526 312976 100188 313032
rect 99465 312974 100188 312976
rect 99465 312971 99531 312974
rect 172421 312354 172487 312357
rect 169924 312352 172487 312354
rect 169924 312296 172426 312352
rect 172482 312296 172487 312352
rect 169924 312294 172487 312296
rect 172421 312291 172487 312294
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect 172053 310858 172119 310861
rect 172053 310856 234630 310858
rect 172053 310800 172058 310856
rect 172114 310800 234630 310856
rect 172053 310798 234630 310800
rect 172053 310795 172119 310798
rect 232313 310722 232379 310725
rect 232814 310722 232820 310724
rect 232313 310720 232820 310722
rect 232313 310664 232318 310720
rect 232374 310664 232820 310720
rect 232313 310662 232820 310664
rect 232313 310659 232379 310662
rect 232814 310660 232820 310662
rect 232884 310660 232890 310724
rect 225689 310586 225755 310589
rect 234429 310586 234495 310589
rect 225689 310584 234495 310586
rect 225689 310528 225694 310584
rect 225750 310528 234434 310584
rect 234490 310528 234495 310584
rect 225689 310526 234495 310528
rect 234570 310586 234630 310798
rect 235809 310586 235875 310589
rect 234570 310584 235875 310586
rect 234570 310528 235814 310584
rect 235870 310528 235875 310584
rect 234570 310526 235875 310528
rect 225689 310523 225755 310526
rect 234429 310523 234495 310526
rect 235809 310523 235875 310526
rect 232814 310388 232820 310452
rect 232884 310450 232890 310452
rect 232957 310450 233023 310453
rect 232884 310448 233023 310450
rect 232884 310392 232962 310448
rect 233018 310392 233023 310448
rect 232884 310390 233023 310392
rect 232884 310388 232890 310390
rect 232957 310387 233023 310390
rect 97257 310314 97323 310317
rect 97257 310312 100188 310314
rect 97257 310256 97262 310312
rect 97318 310256 100188 310312
rect 97257 310254 100188 310256
rect 97257 310251 97323 310254
rect 231117 309906 231183 309909
rect 244641 309906 244707 309909
rect 231117 309904 244707 309906
rect 231117 309848 231122 309904
rect 231178 309848 244646 309904
rect 244702 309848 244707 309904
rect 231117 309846 244707 309848
rect 231117 309843 231183 309846
rect 244641 309843 244707 309846
rect 232630 309708 232636 309772
rect 232700 309770 232706 309772
rect 247309 309770 247375 309773
rect 232700 309768 247375 309770
rect 232700 309712 247314 309768
rect 247370 309712 247375 309768
rect 232700 309710 247375 309712
rect 232700 309708 232706 309710
rect 247309 309707 247375 309710
rect 172421 309634 172487 309637
rect 169924 309632 172487 309634
rect 169924 309576 172426 309632
rect 172482 309576 172487 309632
rect 169924 309574 172487 309576
rect 172421 309571 172487 309574
rect 227069 309634 227135 309637
rect 249057 309634 249123 309637
rect 227069 309632 249123 309634
rect 227069 309576 227074 309632
rect 227130 309576 249062 309632
rect 249118 309576 249123 309632
rect 227069 309574 249123 309576
rect 227069 309571 227135 309574
rect 249057 309571 249123 309574
rect 170765 309498 170831 309501
rect 241237 309498 241303 309501
rect 170765 309496 241303 309498
rect 170765 309440 170770 309496
rect 170826 309440 241242 309496
rect 241298 309440 241303 309496
rect 170765 309438 241303 309440
rect 170765 309435 170831 309438
rect 241237 309435 241303 309438
rect 170949 309362 171015 309365
rect 246389 309362 246455 309365
rect 170949 309360 246455 309362
rect 170949 309304 170954 309360
rect 171010 309304 246394 309360
rect 246450 309304 246455 309360
rect 170949 309302 246455 309304
rect 170949 309299 171015 309302
rect 246389 309299 246455 309302
rect 174721 309226 174787 309229
rect 250621 309226 250687 309229
rect 174721 309224 250687 309226
rect 174721 309168 174726 309224
rect 174782 309168 250626 309224
rect 250682 309168 250687 309224
rect 174721 309166 250687 309168
rect 174721 309163 174787 309166
rect 250621 309163 250687 309166
rect 231301 309090 231367 309093
rect 248321 309090 248387 309093
rect 231301 309088 248387 309090
rect 231301 309032 231306 309088
rect 231362 309032 248326 309088
rect 248382 309032 248387 309088
rect 231301 309030 248387 309032
rect 231301 309027 231367 309030
rect 248321 309027 248387 309030
rect 346761 309090 346827 309093
rect 362125 309090 362191 309093
rect 346761 309088 362191 309090
rect 346761 309032 346766 309088
rect 346822 309032 362130 309088
rect 362186 309032 362191 309088
rect 346761 309030 362191 309032
rect 346761 309027 346827 309030
rect 362125 309027 362191 309030
rect 174629 308954 174695 308957
rect 244273 308954 244339 308957
rect 174629 308952 244339 308954
rect 174629 308896 174634 308952
rect 174690 308896 244278 308952
rect 244334 308896 244339 308952
rect 174629 308894 244339 308896
rect 174629 308891 174695 308894
rect 244273 308891 244339 308894
rect 346945 308954 347011 308957
rect 364977 308954 365043 308957
rect 346945 308952 365043 308954
rect 346945 308896 346950 308952
rect 347006 308896 364982 308952
rect 365038 308896 365043 308952
rect 346945 308894 365043 308896
rect 346945 308891 347011 308894
rect 364977 308891 365043 308894
rect 228633 308818 228699 308821
rect 246573 308818 246639 308821
rect 228633 308816 246639 308818
rect 228633 308760 228638 308816
rect 228694 308760 246578 308816
rect 246634 308760 246639 308816
rect 228633 308758 246639 308760
rect 228633 308755 228699 308758
rect 246573 308755 246639 308758
rect 347497 308818 347563 308821
rect 364885 308818 364951 308821
rect 347497 308816 364951 308818
rect 347497 308760 347502 308816
rect 347558 308760 364890 308816
rect 364946 308760 364951 308816
rect 347497 308758 364951 308760
rect 347497 308755 347563 308758
rect 364885 308755 364951 308758
rect 232446 308620 232452 308684
rect 232516 308682 232522 308684
rect 243353 308682 243419 308685
rect 232516 308680 243419 308682
rect 232516 308624 243358 308680
rect 243414 308624 243419 308680
rect 232516 308622 243419 308624
rect 232516 308620 232522 308622
rect 243353 308619 243419 308622
rect 348417 308682 348483 308685
rect 370129 308682 370195 308685
rect 348417 308680 370195 308682
rect 348417 308624 348422 308680
rect 348478 308624 370134 308680
rect 370190 308624 370195 308680
rect 348417 308622 370195 308624
rect 348417 308619 348483 308622
rect 370129 308619 370195 308622
rect 169334 308484 169340 308548
rect 169404 308546 169410 308548
rect 238017 308546 238083 308549
rect 169404 308544 238083 308546
rect 169404 308488 238022 308544
rect 238078 308488 238083 308544
rect 169404 308486 238083 308488
rect 169404 308484 169410 308486
rect 238017 308483 238083 308486
rect 306097 308546 306163 308549
rect 359958 308546 359964 308548
rect 306097 308544 359964 308546
rect 306097 308488 306102 308544
rect 306158 308488 359964 308544
rect 306097 308486 359964 308488
rect 306097 308483 306163 308486
rect 359958 308484 359964 308486
rect 360028 308484 360034 308548
rect 216581 308410 216647 308413
rect 298461 308410 298527 308413
rect 216581 308408 298527 308410
rect 216581 308352 216586 308408
rect 216642 308352 298466 308408
rect 298522 308352 298527 308408
rect 216581 308350 298527 308352
rect 216581 308347 216647 308350
rect 298461 308347 298527 308350
rect 329925 308410 329991 308413
rect 462957 308410 463023 308413
rect 329925 308408 463023 308410
rect 329925 308352 329930 308408
rect 329986 308352 462962 308408
rect 463018 308352 463023 308408
rect 329925 308350 463023 308352
rect 329925 308347 329991 308350
rect 462957 308347 463023 308350
rect 173249 308274 173315 308277
rect 252645 308274 252711 308277
rect 173249 308272 252711 308274
rect 173249 308216 173254 308272
rect 173310 308216 252650 308272
rect 252706 308216 252711 308272
rect 173249 308214 252711 308216
rect 173249 308211 173315 308214
rect 252645 308211 252711 308214
rect 98545 307594 98611 307597
rect 98545 307592 100188 307594
rect 98545 307536 98550 307592
rect 98606 307536 100188 307592
rect 98545 307534 100188 307536
rect 98545 307531 98611 307534
rect 172421 306914 172487 306917
rect 169924 306912 172487 306914
rect 169924 306856 172426 306912
rect 172482 306856 172487 306912
rect 169924 306854 172487 306856
rect 172421 306851 172487 306854
rect 263961 306506 264027 306509
rect 263918 306504 264027 306506
rect 263918 306448 263966 306504
rect 264022 306448 264027 306504
rect 263918 306443 264027 306448
rect 358118 306444 358124 306508
rect 358188 306506 358194 306508
rect 358353 306506 358419 306509
rect 358188 306504 358419 306506
rect 358188 306448 358358 306504
rect 358414 306448 358419 306504
rect 358188 306446 358419 306448
rect 358188 306444 358194 306446
rect 358353 306443 358419 306446
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 263777 306234 263843 306237
rect 263918 306234 263978 306443
rect 349245 306370 349311 306373
rect 368657 306370 368723 306373
rect 349245 306368 368723 306370
rect 349245 306312 349250 306368
rect 349306 306312 368662 306368
rect 368718 306312 368723 306368
rect 349245 306310 368723 306312
rect 349245 306307 349311 306310
rect 368657 306307 368723 306310
rect 263777 306232 263978 306234
rect 263777 306176 263782 306232
rect 263838 306176 263978 306232
rect 263777 306174 263978 306176
rect 282545 306234 282611 306237
rect 283649 306234 283715 306237
rect 282545 306232 283715 306234
rect 282545 306176 282550 306232
rect 282606 306176 283654 306232
rect 283710 306176 283715 306232
rect 282545 306174 283715 306176
rect 263777 306171 263843 306174
rect 282545 306171 282611 306174
rect 283649 306171 283715 306174
rect 349981 306234 350047 306237
rect 370313 306234 370379 306237
rect 349981 306232 370379 306234
rect 349981 306176 349986 306232
rect 350042 306176 370318 306232
rect 370374 306176 370379 306232
rect 349981 306174 370379 306176
rect 349981 306171 350047 306174
rect 370313 306171 370379 306174
rect 218830 306036 218836 306100
rect 218900 306098 218906 306100
rect 288341 306098 288407 306101
rect 218900 306096 288407 306098
rect 218900 306040 288346 306096
rect 288402 306040 288407 306096
rect 218900 306038 288407 306040
rect 218900 306036 218906 306038
rect 288341 306035 288407 306038
rect 312445 306098 312511 306101
rect 367134 306098 367140 306100
rect 312445 306096 367140 306098
rect 312445 306040 312450 306096
rect 312506 306040 367140 306096
rect 312445 306038 367140 306040
rect 312445 306035 312511 306038
rect 367134 306036 367140 306038
rect 367204 306036 367210 306100
rect 219014 305900 219020 305964
rect 219084 305962 219090 305964
rect 288893 305962 288959 305965
rect 219084 305960 288959 305962
rect 219084 305904 288898 305960
rect 288954 305904 288959 305960
rect 219084 305902 288959 305904
rect 219084 305900 219090 305902
rect 288893 305899 288959 305902
rect 299381 305962 299447 305965
rect 358261 305962 358327 305965
rect 299381 305960 358327 305962
rect 299381 305904 299386 305960
rect 299442 305904 358266 305960
rect 358322 305904 358327 305960
rect 299381 305902 358327 305904
rect 299381 305899 299447 305902
rect 358261 305899 358327 305902
rect 217174 305764 217180 305828
rect 217244 305826 217250 305828
rect 290089 305826 290155 305829
rect 217244 305824 290155 305826
rect 217244 305768 290094 305824
rect 290150 305768 290155 305824
rect 217244 305766 290155 305768
rect 217244 305764 217250 305766
rect 290089 305763 290155 305766
rect 330753 305826 330819 305829
rect 476757 305826 476823 305829
rect 330753 305824 476823 305826
rect 330753 305768 330758 305824
rect 330814 305768 476762 305824
rect 476818 305768 476823 305824
rect 330753 305766 476823 305768
rect 330753 305763 330819 305766
rect 476757 305763 476823 305766
rect 217358 305628 217364 305692
rect 217428 305690 217434 305692
rect 291193 305690 291259 305693
rect 217428 305688 291259 305690
rect 217428 305632 291198 305688
rect 291254 305632 291259 305688
rect 217428 305630 291259 305632
rect 217428 305628 217434 305630
rect 291193 305627 291259 305630
rect 345473 305690 345539 305693
rect 570597 305690 570663 305693
rect 345473 305688 570663 305690
rect 345473 305632 345478 305688
rect 345534 305632 570602 305688
rect 570658 305632 570663 305688
rect 345473 305630 570663 305632
rect 345473 305627 345539 305630
rect 570597 305627 570663 305630
rect 350625 305554 350691 305557
rect 368841 305554 368907 305557
rect 350625 305552 368907 305554
rect 350625 305496 350630 305552
rect 350686 305496 368846 305552
rect 368902 305496 368907 305552
rect 350625 305494 368907 305496
rect 350625 305491 350691 305494
rect 368841 305491 368907 305494
rect 97901 304874 97967 304877
rect 97901 304872 100188 304874
rect 97901 304816 97906 304872
rect 97962 304816 100188 304872
rect 97901 304814 100188 304816
rect 97901 304811 97967 304814
rect 357617 304330 357683 304333
rect 358118 304330 358124 304332
rect 357617 304328 358124 304330
rect 357617 304272 357622 304328
rect 357678 304272 358124 304328
rect 357617 304270 358124 304272
rect 357617 304267 357683 304270
rect 358118 304268 358124 304270
rect 358188 304268 358194 304332
rect 172329 304194 172395 304197
rect 169924 304192 172395 304194
rect 169924 304136 172334 304192
rect 172390 304136 172395 304192
rect 169924 304134 172395 304136
rect 172329 304131 172395 304134
rect 312353 303514 312419 303517
rect 369894 303514 369900 303516
rect 312353 303512 369900 303514
rect 312353 303456 312358 303512
rect 312414 303456 369900 303512
rect 312353 303454 369900 303456
rect 312353 303451 312419 303454
rect 369894 303452 369900 303454
rect 369964 303452 369970 303516
rect 298277 303378 298343 303381
rect 357433 303378 357499 303381
rect 298277 303376 357499 303378
rect 298277 303320 298282 303376
rect 298338 303320 357438 303376
rect 357494 303320 357499 303376
rect 298277 303318 357499 303320
rect 298277 303315 298343 303318
rect 357433 303315 357499 303318
rect 215150 303180 215156 303244
rect 215220 303242 215226 303244
rect 287053 303242 287119 303245
rect 215220 303240 287119 303242
rect 215220 303184 287058 303240
rect 287114 303184 287119 303240
rect 215220 303182 287119 303184
rect 215220 303180 215226 303182
rect 287053 303179 287119 303182
rect 317873 303242 317939 303245
rect 396717 303242 396783 303245
rect 317873 303240 396783 303242
rect 317873 303184 317878 303240
rect 317934 303184 396722 303240
rect 396778 303184 396783 303240
rect 317873 303182 396783 303184
rect 317873 303179 317939 303182
rect 396717 303179 396783 303182
rect 216254 303044 216260 303108
rect 216324 303106 216330 303108
rect 288709 303106 288775 303109
rect 216324 303104 288775 303106
rect 216324 303048 288714 303104
rect 288770 303048 288775 303104
rect 216324 303046 288775 303048
rect 216324 303044 216330 303046
rect 288709 303043 288775 303046
rect 331857 303106 331923 303109
rect 489177 303106 489243 303109
rect 331857 303104 489243 303106
rect 331857 303048 331862 303104
rect 331918 303048 489182 303104
rect 489238 303048 489243 303104
rect 331857 303046 489243 303048
rect 331857 303043 331923 303046
rect 489177 303043 489243 303046
rect 170489 302970 170555 302973
rect 260189 302970 260255 302973
rect 170489 302968 260255 302970
rect 170489 302912 170494 302968
rect 170550 302912 260194 302968
rect 260250 302912 260255 302968
rect 170489 302910 260255 302912
rect 170489 302907 170555 302910
rect 260189 302907 260255 302910
rect 337285 302970 337351 302973
rect 520917 302970 520983 302973
rect 337285 302968 520983 302970
rect 337285 302912 337290 302968
rect 337346 302912 520922 302968
rect 520978 302912 520983 302968
rect 337285 302910 520983 302912
rect 337285 302907 337351 302910
rect 520917 302907 520983 302910
rect 182173 302834 182239 302837
rect 282177 302834 282243 302837
rect 182173 302832 282243 302834
rect 182173 302776 182178 302832
rect 182234 302776 282182 302832
rect 282238 302776 282243 302832
rect 182173 302774 282243 302776
rect 182173 302771 182239 302774
rect 282177 302771 282243 302774
rect 339953 302834 340019 302837
rect 539685 302834 539751 302837
rect 339953 302832 539751 302834
rect 339953 302776 339958 302832
rect 340014 302776 539690 302832
rect 539746 302776 539751 302832
rect 339953 302774 539751 302776
rect 339953 302771 340019 302774
rect 539685 302771 539751 302774
rect 99833 302154 99899 302157
rect 99833 302152 100188 302154
rect 99833 302096 99838 302152
rect 99894 302096 100188 302152
rect 99833 302094 100188 302096
rect 99833 302091 99899 302094
rect 219198 301684 219204 301748
rect 219268 301746 219274 301748
rect 287421 301746 287487 301749
rect 219268 301744 287487 301746
rect 219268 301688 287426 301744
rect 287482 301688 287487 301744
rect 219268 301686 287487 301688
rect 219268 301684 219274 301686
rect 287421 301683 287487 301686
rect 169702 301548 169708 301612
rect 169772 301610 169778 301612
rect 239029 301610 239095 301613
rect 169772 301608 239095 301610
rect 169772 301552 239034 301608
rect 239090 301552 239095 301608
rect 169772 301550 239095 301552
rect 169772 301548 169778 301550
rect 239029 301547 239095 301550
rect 172421 301474 172487 301477
rect 169924 301472 172487 301474
rect 169924 301416 172426 301472
rect 172482 301416 172487 301472
rect 169924 301414 172487 301416
rect 172421 301411 172487 301414
rect 216990 301412 216996 301476
rect 217060 301474 217066 301476
rect 292941 301474 293007 301477
rect 217060 301472 293007 301474
rect 217060 301416 292946 301472
rect 293002 301416 293007 301472
rect 217060 301414 293007 301416
rect 217060 301412 217066 301414
rect 292941 301411 293007 301414
rect 169150 301140 169156 301204
rect 169220 301202 169226 301204
rect 248505 301202 248571 301205
rect 169220 301200 248571 301202
rect 169220 301144 248510 301200
rect 248566 301144 248571 301200
rect 169220 301142 248571 301144
rect 169220 301140 169226 301142
rect 248505 301139 248571 301142
rect 99281 300794 99347 300797
rect 245837 300794 245903 300797
rect 99281 300792 245903 300794
rect 99281 300736 99286 300792
rect 99342 300736 245842 300792
rect 245898 300736 245903 300792
rect 99281 300734 245903 300736
rect 99281 300731 99347 300734
rect 245837 300731 245903 300734
rect 164233 300386 164299 300389
rect 279325 300386 279391 300389
rect 164233 300384 279391 300386
rect 164233 300328 164238 300384
rect 164294 300328 279330 300384
rect 279386 300328 279391 300384
rect 164233 300326 279391 300328
rect 164233 300323 164299 300326
rect 279325 300323 279391 300326
rect 160093 300250 160159 300253
rect 278589 300250 278655 300253
rect 160093 300248 278655 300250
rect 160093 300192 160098 300248
rect 160154 300192 278594 300248
rect 278650 300192 278655 300248
rect 160093 300190 278655 300192
rect 160093 300187 160159 300190
rect 278589 300187 278655 300190
rect 34513 300114 34579 300117
rect 258533 300114 258599 300117
rect 34513 300112 258599 300114
rect 34513 300056 34518 300112
rect 34574 300056 258538 300112
rect 258594 300056 258599 300112
rect 34513 300054 258599 300056
rect 34513 300051 34579 300054
rect 258533 300051 258599 300054
rect 300025 300114 300091 300117
rect 368606 300114 368612 300116
rect 300025 300112 368612 300114
rect 300025 300056 300030 300112
rect 300086 300056 368612 300112
rect 300025 300054 368612 300056
rect 300025 300051 300091 300054
rect 368606 300052 368612 300054
rect 368676 300052 368682 300116
rect 97533 299434 97599 299437
rect 249885 299434 249951 299437
rect 97533 299432 249951 299434
rect 97533 299376 97538 299432
rect 97594 299376 249890 299432
rect 249946 299376 249951 299432
rect 97533 299374 249951 299376
rect 97533 299371 97599 299374
rect 249885 299371 249951 299374
rect 99189 299298 99255 299301
rect 234337 299298 234403 299301
rect 99189 299296 234403 299298
rect 99189 299240 99194 299296
rect 99250 299240 234342 299296
rect 234398 299240 234403 299296
rect 99189 299238 234403 299240
rect 99189 299235 99255 299238
rect 234337 299235 234403 299238
rect 97257 299162 97323 299165
rect 169334 299162 169340 299164
rect 97257 299160 169340 299162
rect 97257 299104 97262 299160
rect 97318 299104 169340 299160
rect 97257 299102 169340 299104
rect 97257 299099 97323 299102
rect 169334 299100 169340 299102
rect 169404 299100 169410 299164
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 97349 298074 97415 298077
rect 237649 298074 237715 298077
rect 97349 298072 237715 298074
rect 97349 298016 97354 298072
rect 97410 298016 237654 298072
rect 237710 298016 237715 298072
rect 97349 298014 237715 298016
rect 97349 298011 97415 298014
rect 237649 298011 237715 298014
rect 109677 297938 109743 297941
rect 169150 297938 169156 297940
rect 109677 297936 169156 297938
rect 109677 297880 109682 297936
rect 109738 297880 169156 297936
rect 109677 297878 169156 297880
rect 109677 297875 109743 297878
rect 169150 297876 169156 297878
rect 169220 297876 169226 297940
rect 150893 297802 150959 297805
rect 169702 297802 169708 297804
rect 150893 297800 169708 297802
rect 150893 297744 150898 297800
rect 150954 297744 169708 297800
rect 150893 297742 169708 297744
rect 150893 297739 150959 297742
rect 169702 297740 169708 297742
rect 169772 297740 169778 297804
rect 213545 297666 213611 297669
rect 291653 297666 291719 297669
rect 213545 297664 291719 297666
rect 213545 297608 213550 297664
rect 213606 297608 291658 297664
rect 291714 297608 291719 297664
rect 213545 297606 291719 297608
rect 213545 297603 213611 297606
rect 291653 297603 291719 297606
rect 211981 297530 212047 297533
rect 290181 297530 290247 297533
rect 211981 297528 290247 297530
rect 211981 297472 211986 297528
rect 212042 297472 290186 297528
rect 290242 297472 290247 297528
rect 211981 297470 290247 297472
rect 211981 297467 212047 297470
rect 290181 297467 290247 297470
rect 212349 297394 212415 297397
rect 291561 297394 291627 297397
rect 212349 297392 291627 297394
rect 212349 297336 212354 297392
rect 212410 297336 291566 297392
rect 291622 297336 291627 297392
rect 212349 297334 291627 297336
rect 212349 297331 212415 297334
rect 291561 297331 291627 297334
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect 214414 284820 214420 284884
rect 214484 284882 214490 284884
rect 285949 284882 286015 284885
rect 214484 284880 286015 284882
rect 214484 284824 285954 284880
rect 286010 284824 286015 284880
rect 214484 284822 286015 284824
rect 214484 284820 214490 284822
rect 285949 284819 286015 284822
rect 312077 280802 312143 280805
rect 368422 280802 368428 280804
rect 312077 280800 368428 280802
rect 312077 280744 312082 280800
rect 312138 280744 368428 280800
rect 312077 280742 368428 280744
rect 312077 280739 312143 280742
rect 368422 280740 368428 280742
rect 368492 280740 368498 280804
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 215886 269724 215892 269788
rect 215956 269786 215962 269788
rect 286133 269786 286199 269789
rect 215956 269784 286199 269786
rect 215956 269728 286138 269784
rect 286194 269728 286199 269784
rect 215956 269726 286199 269728
rect 215956 269724 215962 269726
rect 286133 269723 286199 269726
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 313365 265570 313431 265573
rect 369158 265570 369164 265572
rect 313365 265568 369164 265570
rect 313365 265512 313370 265568
rect 313426 265512 369164 265568
rect 313365 265510 369164 265512
rect 313365 265507 313431 265510
rect 369158 265508 369164 265510
rect 369228 265508 369234 265572
rect 311249 260266 311315 260269
rect 361614 260266 361620 260268
rect 311249 260264 361620 260266
rect 311249 260208 311254 260264
rect 311310 260208 361620 260264
rect 311249 260206 361620 260208
rect 311249 260203 311315 260206
rect 361614 260204 361620 260206
rect 361684 260204 361690 260268
rect 311065 260130 311131 260133
rect 365662 260130 365668 260132
rect 311065 260128 365668 260130
rect 311065 260072 311070 260128
rect 311126 260072 365668 260128
rect 311065 260070 365668 260072
rect 311065 260067 311131 260070
rect 365662 260068 365668 260070
rect 365732 260068 365738 260132
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 216438 254492 216444 254556
rect 216508 254554 216514 254556
rect 287145 254554 287211 254557
rect 216508 254552 287211 254554
rect 216508 254496 287150 254552
rect 287206 254496 287211 254552
rect 216508 254494 287211 254496
rect 216508 254492 216514 254494
rect 287145 254491 287211 254494
rect 310973 254554 311039 254557
rect 364374 254554 364380 254556
rect 310973 254552 364380 254554
rect 310973 254496 310978 254552
rect 311034 254496 364380 254552
rect 310973 254494 364380 254496
rect 310973 254491 311039 254494
rect 364374 254492 364380 254494
rect 364444 254492 364450 254556
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 310789 251834 310855 251837
rect 365846 251834 365852 251836
rect 310789 251832 365852 251834
rect 310789 251776 310794 251832
rect 310850 251776 365852 251832
rect 310789 251774 365852 251776
rect 310789 251771 310855 251774
rect 365846 251772 365852 251774
rect 365916 251772 365922 251836
rect 310881 251018 310947 251021
rect 358854 251018 358860 251020
rect 310881 251016 358860 251018
rect 310881 250960 310886 251016
rect 310942 250960 358860 251016
rect 310881 250958 358860 250960
rect 310881 250955 310947 250958
rect 358854 250956 358860 250958
rect 358924 250956 358930 251020
rect 310697 250882 310763 250885
rect 362902 250882 362908 250884
rect 310697 250880 362908 250882
rect 310697 250824 310702 250880
rect 310758 250824 362908 250880
rect 310697 250822 362908 250824
rect 310697 250819 310763 250822
rect 362902 250820 362908 250822
rect 362972 250820 362978 250884
rect 305545 250746 305611 250749
rect 359038 250746 359044 250748
rect 305545 250744 359044 250746
rect 305545 250688 305550 250744
rect 305606 250688 359044 250744
rect 305545 250686 359044 250688
rect 305545 250683 305611 250686
rect 359038 250684 359044 250686
rect 359108 250684 359114 250748
rect 303797 250610 303863 250613
rect 358302 250610 358308 250612
rect 303797 250608 358308 250610
rect 303797 250552 303802 250608
rect 303858 250552 358308 250608
rect 303797 250550 358308 250552
rect 303797 250547 303863 250550
rect 358302 250548 358308 250550
rect 358372 250548 358378 250612
rect 217542 250412 217548 250476
rect 217612 250474 217618 250476
rect 287513 250474 287579 250477
rect 217612 250472 287579 250474
rect 217612 250416 287518 250472
rect 287574 250416 287579 250472
rect 217612 250414 287579 250416
rect 217612 250412 217618 250414
rect 287513 250411 287579 250414
rect 308305 250474 308371 250477
rect 364558 250474 364564 250476
rect 308305 250472 364564 250474
rect 308305 250416 308310 250472
rect 308366 250416 364564 250472
rect 308305 250414 364564 250416
rect 308305 250411 308371 250414
rect 364558 250412 364564 250414
rect 364628 250412 364634 250476
rect 310605 248162 310671 248165
rect 360326 248162 360332 248164
rect 310605 248160 360332 248162
rect 310605 248104 310610 248160
rect 310666 248104 360332 248160
rect 310605 248102 360332 248104
rect 310605 248099 310671 248102
rect 360326 248100 360332 248102
rect 360396 248100 360402 248164
rect 305269 248026 305335 248029
rect 358118 248026 358124 248028
rect 305269 248024 358124 248026
rect 305269 247968 305274 248024
rect 305330 247968 358124 248024
rect 305269 247966 358124 247968
rect 305269 247963 305335 247966
rect 358118 247964 358124 247966
rect 358188 247964 358194 248028
rect 309225 247890 309291 247893
rect 363270 247890 363276 247892
rect 309225 247888 363276 247890
rect 309225 247832 309230 247888
rect 309286 247832 363276 247888
rect 309225 247830 363276 247832
rect 309225 247827 309291 247830
rect 363270 247828 363276 247830
rect 363340 247828 363346 247892
rect 308029 247754 308095 247757
rect 363454 247754 363460 247756
rect 308029 247752 363460 247754
rect 308029 247696 308034 247752
rect 308090 247696 363460 247752
rect 308029 247694 363460 247696
rect 308029 247691 308095 247694
rect 363454 247692 363460 247694
rect 363524 247692 363530 247756
rect 306557 247618 306623 247621
rect 363086 247618 363092 247620
rect 306557 247616 363092 247618
rect 306557 247560 306562 247616
rect 306618 247560 363092 247616
rect 306557 247558 363092 247560
rect 306557 247555 306623 247558
rect 363086 247556 363092 247558
rect 363156 247556 363162 247620
rect 309317 245578 309383 245581
rect 360694 245578 360700 245580
rect 309317 245576 360700 245578
rect 309317 245520 309322 245576
rect 309378 245520 360700 245576
rect 309317 245518 360700 245520
rect 309317 245515 309383 245518
rect 360694 245516 360700 245518
rect 360764 245516 360770 245580
rect 578877 245578 578943 245581
rect 583520 245578 584960 245668
rect 578877 245576 584960 245578
rect 578877 245520 578882 245576
rect 578938 245520 584960 245576
rect 578877 245518 584960 245520
rect 578877 245515 578943 245518
rect 306465 245442 306531 245445
rect 359406 245442 359412 245444
rect 306465 245440 359412 245442
rect 306465 245384 306470 245440
rect 306526 245384 359412 245440
rect 306465 245382 359412 245384
rect 306465 245379 306531 245382
rect 359406 245380 359412 245382
rect 359476 245380 359482 245444
rect 583520 245428 584960 245518
rect 309133 245306 309199 245309
rect 362534 245306 362540 245308
rect 309133 245304 362540 245306
rect 309133 245248 309138 245304
rect 309194 245248 362540 245304
rect 309133 245246 362540 245248
rect 309133 245243 309199 245246
rect 362534 245244 362540 245246
rect 362604 245244 362610 245308
rect 305177 245170 305243 245173
rect 359222 245170 359228 245172
rect 305177 245168 359228 245170
rect 305177 245112 305182 245168
rect 305238 245112 359228 245168
rect 305177 245110 359228 245112
rect 305177 245107 305243 245110
rect 359222 245108 359228 245110
rect 359292 245108 359298 245172
rect 304993 245034 305059 245037
rect 360510 245034 360516 245036
rect 304993 245032 360516 245034
rect 304993 244976 304998 245032
rect 305054 244976 360516 245032
rect 304993 244974 360516 244976
rect 304993 244971 305059 244974
rect 360510 244972 360516 244974
rect 360580 244972 360586 245036
rect 303705 244898 303771 244901
rect 367318 244898 367324 244900
rect 303705 244896 367324 244898
rect 303705 244840 303710 244896
rect 303766 244840 367324 244896
rect 303705 244838 367324 244840
rect 303705 244835 303771 244838
rect 367318 244836 367324 244838
rect 367388 244836 367394 244900
rect 310513 244762 310579 244765
rect 358486 244762 358492 244764
rect 310513 244760 358492 244762
rect 310513 244704 310518 244760
rect 310574 244704 358492 244760
rect 310513 244702 358492 244704
rect 310513 244699 310579 244702
rect 358486 244700 358492 244702
rect 358556 244700 358562 244764
rect 359641 243674 359707 243677
rect 354630 243672 359707 243674
rect 354630 243616 359646 243672
rect 359702 243616 359707 243672
rect 354630 243614 359707 243616
rect 218421 243538 218487 243541
rect 218646 243538 218652 243540
rect 218421 243536 218652 243538
rect 218421 243480 218426 243536
rect 218482 243480 218652 243536
rect 218421 243478 218652 243480
rect 218421 243475 218487 243478
rect 218646 243476 218652 243478
rect 218716 243476 218722 243540
rect 298093 243538 298159 243541
rect 354630 243538 354690 243614
rect 359641 243611 359707 243614
rect 298093 243536 354690 243538
rect 298093 243480 298098 243536
rect 298154 243480 354690 243536
rect 298093 243478 354690 243480
rect 356881 243538 356947 243541
rect 357566 243538 357572 243540
rect 356881 243536 357572 243538
rect 356881 243480 356886 243536
rect 356942 243480 357572 243536
rect 356881 243478 357572 243480
rect 298093 243475 298159 243478
rect 356881 243475 356947 243478
rect 357566 243476 357572 243478
rect 357636 243476 357642 243540
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580901 232386 580967 232389
rect 583520 232386 584960 232476
rect 580901 232384 584960 232386
rect 580901 232328 580906 232384
rect 580962 232328 584960 232384
rect 580901 232326 584960 232328
rect 580901 232323 580967 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580809 219058 580875 219061
rect 583520 219058 584960 219148
rect 580809 219056 584960 219058
rect 580809 219000 580814 219056
rect 580870 219000 584960 219056
rect 580809 218998 584960 219000
rect 580809 218995 580875 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 217685 196890 217751 196893
rect 219390 196890 220064 196924
rect 217685 196888 220064 196890
rect 217685 196832 217690 196888
rect 217746 196864 220064 196888
rect 217746 196832 219450 196864
rect 217685 196830 219450 196832
rect 217685 196827 217751 196830
rect 217225 195938 217291 195941
rect 219390 195938 220064 195972
rect 217225 195936 220064 195938
rect 217225 195880 217230 195936
rect 217286 195912 220064 195936
rect 217286 195880 219450 195912
rect 217225 195878 219450 195880
rect 217225 195875 217291 195878
rect 217593 193762 217659 193765
rect 219390 193762 220064 193796
rect 217593 193760 220064 193762
rect 217593 193704 217598 193760
rect 217654 193736 220064 193760
rect 217654 193704 219450 193736
rect 217593 193702 219450 193704
rect 217593 193699 217659 193702
rect 217133 192810 217199 192813
rect 219390 192810 220064 192844
rect 217133 192808 220064 192810
rect 217133 192752 217138 192808
rect 217194 192784 220064 192808
rect 217194 192752 219450 192784
rect 217133 192750 219450 192752
rect 217133 192747 217199 192750
rect 580809 192538 580875 192541
rect 583520 192538 584960 192628
rect 580809 192536 584960 192538
rect 580809 192480 580814 192536
rect 580870 192480 584960 192536
rect 580809 192478 584960 192480
rect 580809 192475 580875 192478
rect 583520 192388 584960 192478
rect 218697 191042 218763 191045
rect 219390 191042 220064 191076
rect 218697 191040 220064 191042
rect 218697 190984 218702 191040
rect 218758 191016 220064 191040
rect 218758 190984 219450 191016
rect 218697 190982 219450 190984
rect 218697 190979 218763 190982
rect 218513 189954 218579 189957
rect 219390 189954 220064 189988
rect 218513 189952 220064 189954
rect 218513 189896 218518 189952
rect 218574 189928 220064 189952
rect 218574 189896 219450 189928
rect 218513 189894 219450 189896
rect 218513 189891 218579 189894
rect -960 188866 480 188956
rect -960 188806 674 188866
rect -960 188730 480 188806
rect 614 188730 674 188806
rect -960 188716 674 188730
rect 246 188670 674 188716
rect 246 188186 306 188670
rect 218605 188186 218671 188189
rect 219390 188186 220064 188220
rect 246 188126 6930 188186
rect 6870 187778 6930 188126
rect 218605 188184 220064 188186
rect 218605 188128 218610 188184
rect 218666 188160 220064 188184
rect 218666 188128 219450 188160
rect 218605 188126 219450 188128
rect 218605 188123 218671 188126
rect 216070 187778 216076 187780
rect 6870 187718 216076 187778
rect 216070 187716 216076 187718
rect 216140 187716 216146 187780
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 367870 178060 367876 178124
rect 367940 178122 367946 178124
rect 583526 178122 583586 179014
rect 367940 178062 583586 178122
rect 367940 178060 367946 178062
rect -960 175796 480 176036
rect 217501 169962 217567 169965
rect 219390 169962 220064 169996
rect 217501 169960 220064 169962
rect 217501 169904 217506 169960
rect 217562 169936 220064 169960
rect 217562 169904 219450 169936
rect 217501 169902 219450 169904
rect 217501 169899 217567 169902
rect 217777 168330 217843 168333
rect 219390 168330 220064 168364
rect 217777 168328 220064 168330
rect 217777 168272 217782 168328
rect 217838 168304 220064 168328
rect 217838 168272 219450 168304
rect 217777 168270 219450 168272
rect 217777 168267 217843 168270
rect 217317 168058 217383 168061
rect 219390 168058 220064 168092
rect 217317 168056 220064 168058
rect 217317 168000 217322 168056
rect 217378 168032 220064 168056
rect 217378 168000 219450 168032
rect 217317 167998 219450 168000
rect 217317 167995 217383 167998
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 214598 162890 214604 162892
rect -960 162830 214604 162890
rect -960 162740 480 162830
rect 214598 162828 214604 162830
rect 214668 162828 214674 162892
rect 356830 160108 356836 160172
rect 356900 160170 356906 160172
rect 358261 160170 358327 160173
rect 356900 160168 358327 160170
rect 356900 160112 358266 160168
rect 358322 160112 358327 160168
rect 356900 160110 358327 160112
rect 356900 160108 356906 160110
rect 358261 160107 358327 160110
rect 363454 160108 363460 160172
rect 363524 160170 363530 160172
rect 363873 160170 363939 160173
rect 363524 160168 363939 160170
rect 363524 160112 363878 160168
rect 363934 160112 363939 160168
rect 363524 160110 363939 160112
rect 363524 160108 363530 160110
rect 363873 160107 363939 160110
rect 278129 159900 278195 159901
rect 278072 159898 278078 159900
rect 278038 159838 278078 159898
rect 278142 159896 278195 159900
rect 278190 159840 278195 159896
rect 278072 159836 278078 159838
rect 278142 159836 278195 159840
rect 278129 159835 278195 159836
rect 300945 159764 301011 159765
rect 300920 159762 300926 159764
rect 300854 159702 300926 159762
rect 300990 159760 301011 159764
rect 301006 159704 301011 159760
rect 300920 159700 300926 159702
rect 300990 159700 301011 159704
rect 300945 159699 301011 159700
rect 271045 159628 271111 159629
rect 275829 159628 275895 159629
rect 279233 159628 279299 159629
rect 288341 159628 288407 159629
rect 258488 159564 258494 159628
rect 258558 159564 258564 159628
rect 271000 159626 271006 159628
rect 270954 159566 271006 159626
rect 271070 159624 271111 159628
rect 275760 159626 275766 159628
rect 271106 159568 271111 159624
rect 271000 159564 271006 159566
rect 271070 159564 271111 159568
rect 275738 159566 275766 159626
rect 275760 159564 275766 159566
rect 275830 159624 275895 159628
rect 279160 159626 279166 159628
rect 275830 159568 275834 159624
rect 275890 159568 275895 159624
rect 275830 159564 275895 159568
rect 279142 159566 279166 159626
rect 279160 159564 279166 159566
rect 279230 159624 279299 159628
rect 288272 159626 288278 159628
rect 279230 159568 279238 159624
rect 279294 159568 279299 159624
rect 279230 159564 279299 159568
rect 288250 159566 288278 159626
rect 288272 159564 288278 159566
rect 288342 159624 288407 159628
rect 288342 159568 288346 159624
rect 288402 159568 288407 159624
rect 288342 159564 288407 159568
rect 258496 159354 258556 159564
rect 271045 159563 271111 159564
rect 275829 159563 275895 159564
rect 279233 159563 279299 159564
rect 288341 159563 288407 159564
rect 295885 159628 295951 159629
rect 295885 159624 295894 159628
rect 295958 159626 295964 159628
rect 357341 159626 357407 159629
rect 362125 159626 362191 159629
rect 295885 159568 295890 159624
rect 295885 159564 295894 159568
rect 295958 159566 296042 159626
rect 357341 159624 362191 159626
rect 357341 159568 357346 159624
rect 357402 159568 362130 159624
rect 362186 159568 362191 159624
rect 357341 159566 362191 159568
rect 295958 159564 295964 159566
rect 295885 159563 295951 159564
rect 357341 159563 357407 159566
rect 362125 159563 362191 159566
rect 265934 159428 265940 159492
rect 266004 159490 266010 159492
rect 374361 159490 374427 159493
rect 266004 159488 374427 159490
rect 266004 159432 374366 159488
rect 374422 159432 374427 159488
rect 266004 159430 374427 159432
rect 266004 159428 266010 159430
rect 374361 159427 374427 159430
rect 370589 159354 370655 159357
rect 258496 159352 370655 159354
rect 258496 159296 370594 159352
rect 370650 159296 370655 159352
rect 258496 159294 370655 159296
rect 370589 159291 370655 159294
rect 250846 159156 250852 159220
rect 250916 159218 250922 159220
rect 367921 159218 367987 159221
rect 250916 159216 367987 159218
rect 250916 159160 367926 159216
rect 367982 159160 367987 159216
rect 250916 159158 367987 159160
rect 250916 159156 250922 159158
rect 367921 159155 367987 159158
rect 243118 159020 243124 159084
rect 243188 159082 243194 159084
rect 243188 159022 364350 159082
rect 243188 159020 243194 159022
rect 236126 158884 236132 158948
rect 236196 158946 236202 158948
rect 357341 158946 357407 158949
rect 236196 158944 357407 158946
rect 236196 158888 357346 158944
rect 357402 158888 357407 158944
rect 236196 158886 357407 158888
rect 236196 158884 236202 158886
rect 357341 158883 357407 158886
rect 357566 158884 357572 158948
rect 357636 158946 357642 158948
rect 358353 158946 358419 158949
rect 362493 158948 362559 158949
rect 362493 158946 362540 158948
rect 357636 158944 358419 158946
rect 357636 158888 358358 158944
rect 358414 158888 358419 158944
rect 357636 158886 358419 158888
rect 362448 158944 362540 158946
rect 362448 158888 362498 158944
rect 362448 158886 362540 158888
rect 357636 158884 357642 158886
rect 358353 158883 358419 158886
rect 362493 158884 362540 158886
rect 362604 158884 362610 158948
rect 364290 158946 364350 159022
rect 364977 158946 365043 158949
rect 364290 158944 365043 158946
rect 364290 158888 364982 158944
rect 365038 158888 365043 158944
rect 364290 158886 365043 158888
rect 362493 158883 362559 158884
rect 364977 158883 365043 158886
rect 237230 158748 237236 158812
rect 237300 158810 237306 158812
rect 364885 158810 364951 158813
rect 237300 158808 364951 158810
rect 237300 158752 364890 158808
rect 364946 158752 364951 158808
rect 237300 158750 364951 158752
rect 237300 158748 237306 158750
rect 364885 158747 364951 158750
rect 218830 158612 218836 158676
rect 218900 158674 218906 158676
rect 220813 158674 220879 158677
rect 218900 158672 220879 158674
rect 218900 158616 220818 158672
rect 220874 158616 220879 158672
rect 218900 158614 220879 158616
rect 218900 158612 218906 158614
rect 220813 158611 220879 158614
rect 238109 158676 238175 158677
rect 239581 158676 239647 158677
rect 238109 158672 238156 158676
rect 238220 158674 238226 158676
rect 238109 158616 238114 158672
rect 238109 158612 238156 158616
rect 238220 158614 238266 158674
rect 239581 158672 239628 158676
rect 239692 158674 239698 158676
rect 239581 158616 239586 158672
rect 238220 158612 238226 158614
rect 239581 158612 239628 158616
rect 239692 158614 239738 158674
rect 239692 158612 239698 158614
rect 240542 158612 240548 158676
rect 240612 158674 240618 158676
rect 240685 158674 240751 158677
rect 248321 158676 248387 158677
rect 248270 158674 248276 158676
rect 240612 158672 240751 158674
rect 240612 158616 240690 158672
rect 240746 158616 240751 158672
rect 240612 158614 240751 158616
rect 248230 158614 248276 158674
rect 248340 158672 248387 158676
rect 248382 158616 248387 158672
rect 240612 158612 240618 158614
rect 238109 158611 238175 158612
rect 239581 158611 239647 158612
rect 240685 158611 240751 158614
rect 248270 158612 248276 158614
rect 248340 158612 248387 158616
rect 250110 158612 250116 158676
rect 250180 158674 250186 158676
rect 250437 158674 250503 158677
rect 252369 158676 252435 158677
rect 252318 158674 252324 158676
rect 250180 158672 250503 158674
rect 250180 158616 250442 158672
rect 250498 158616 250503 158672
rect 250180 158614 250503 158616
rect 252278 158614 252324 158674
rect 252388 158672 252435 158676
rect 252430 158616 252435 158672
rect 250180 158612 250186 158614
rect 248321 158611 248387 158612
rect 250437 158611 250503 158614
rect 252318 158612 252324 158614
rect 252388 158612 252435 158616
rect 254526 158612 254532 158676
rect 254596 158674 254602 158676
rect 254945 158674 255011 158677
rect 255865 158676 255931 158677
rect 255814 158674 255820 158676
rect 254596 158672 255011 158674
rect 254596 158616 254950 158672
rect 255006 158616 255011 158672
rect 254596 158614 255011 158616
rect 255774 158614 255820 158674
rect 255884 158672 255931 158676
rect 255926 158616 255931 158672
rect 254596 158612 254602 158614
rect 252369 158611 252435 158612
rect 254945 158611 255011 158614
rect 255814 158612 255820 158614
rect 255884 158612 255931 158616
rect 257102 158612 257108 158676
rect 257172 158674 257178 158676
rect 257245 158674 257311 158677
rect 257172 158672 257311 158674
rect 257172 158616 257250 158672
rect 257306 158616 257311 158672
rect 257172 158614 257311 158616
rect 257172 158612 257178 158614
rect 255865 158611 255931 158612
rect 257245 158611 257311 158614
rect 258206 158612 258212 158676
rect 258276 158674 258282 158676
rect 259085 158674 259151 158677
rect 259545 158676 259611 158677
rect 259494 158674 259500 158676
rect 258276 158672 259151 158674
rect 258276 158616 259090 158672
rect 259146 158616 259151 158672
rect 258276 158614 259151 158616
rect 259454 158614 259500 158674
rect 259564 158672 259611 158676
rect 259606 158616 259611 158672
rect 258276 158612 258282 158614
rect 259085 158611 259151 158614
rect 259494 158612 259500 158614
rect 259564 158612 259611 158616
rect 261150 158612 261156 158676
rect 261220 158674 261226 158676
rect 261477 158674 261543 158677
rect 262857 158676 262923 158677
rect 263593 158676 263659 158677
rect 268745 158676 268811 158677
rect 269849 158676 269915 158677
rect 271137 158676 271203 158677
rect 272241 158676 272307 158677
rect 274449 158676 274515 158677
rect 277025 158676 277091 158677
rect 298553 158676 298619 158677
rect 303521 158676 303587 158677
rect 306097 158676 306163 158677
rect 262806 158674 262812 158676
rect 261220 158672 261543 158674
rect 261220 158616 261482 158672
rect 261538 158616 261543 158672
rect 261220 158614 261543 158616
rect 262766 158614 262812 158674
rect 262876 158672 262923 158676
rect 263542 158674 263548 158676
rect 262918 158616 262923 158672
rect 261220 158612 261226 158614
rect 259545 158611 259611 158612
rect 261477 158611 261543 158614
rect 262806 158612 262812 158614
rect 262876 158612 262923 158616
rect 263502 158614 263548 158674
rect 263612 158672 263659 158676
rect 268694 158674 268700 158676
rect 263654 158616 263659 158672
rect 263542 158612 263548 158614
rect 263612 158612 263659 158616
rect 268654 158614 268700 158674
rect 268764 158672 268811 158676
rect 269798 158674 269804 158676
rect 268806 158616 268811 158672
rect 268694 158612 268700 158614
rect 268764 158612 268811 158616
rect 269758 158614 269804 158674
rect 269868 158672 269915 158676
rect 271086 158674 271092 158676
rect 269910 158616 269915 158672
rect 269798 158612 269804 158614
rect 269868 158612 269915 158616
rect 271046 158614 271092 158674
rect 271156 158672 271203 158676
rect 272190 158674 272196 158676
rect 271198 158616 271203 158672
rect 271086 158612 271092 158614
rect 271156 158612 271203 158616
rect 272150 158614 272196 158674
rect 272260 158672 272307 158676
rect 274398 158674 274404 158676
rect 272302 158616 272307 158672
rect 272190 158612 272196 158614
rect 272260 158612 272307 158616
rect 274358 158614 274404 158674
rect 274468 158672 274515 158676
rect 276974 158674 276980 158676
rect 274510 158616 274515 158672
rect 274398 158612 274404 158614
rect 274468 158612 274515 158616
rect 276934 158614 276980 158674
rect 277044 158672 277091 158676
rect 298502 158674 298508 158676
rect 277086 158616 277091 158672
rect 276974 158612 276980 158614
rect 277044 158612 277091 158616
rect 298462 158614 298508 158674
rect 298572 158672 298619 158676
rect 303470 158674 303476 158676
rect 298614 158616 298619 158672
rect 298502 158612 298508 158614
rect 298572 158612 298619 158616
rect 303430 158614 303476 158674
rect 303540 158672 303587 158676
rect 306046 158674 306052 158676
rect 303582 158616 303587 158672
rect 303470 158612 303476 158614
rect 303540 158612 303587 158616
rect 306006 158614 306052 158674
rect 306116 158672 306163 158676
rect 306158 158616 306163 158672
rect 306046 158612 306052 158614
rect 306116 158612 306163 158616
rect 308622 158612 308628 158676
rect 308692 158674 308698 158676
rect 308765 158674 308831 158677
rect 313457 158676 313523 158677
rect 315849 158676 315915 158677
rect 318609 158676 318675 158677
rect 321001 158676 321067 158677
rect 323393 158676 323459 158677
rect 325969 158676 326035 158677
rect 313406 158674 313412 158676
rect 308692 158672 308831 158674
rect 308692 158616 308770 158672
rect 308826 158616 308831 158672
rect 308692 158614 308831 158616
rect 313366 158614 313412 158674
rect 313476 158672 313523 158676
rect 315798 158674 315804 158676
rect 313518 158616 313523 158672
rect 308692 158612 308698 158614
rect 262857 158611 262923 158612
rect 263593 158611 263659 158612
rect 268745 158611 268811 158612
rect 269849 158611 269915 158612
rect 271137 158611 271203 158612
rect 272241 158611 272307 158612
rect 274449 158611 274515 158612
rect 277025 158611 277091 158612
rect 298553 158611 298619 158612
rect 303521 158611 303587 158612
rect 306097 158611 306163 158612
rect 308765 158611 308831 158614
rect 313406 158612 313412 158614
rect 313476 158612 313523 158616
rect 315758 158614 315804 158674
rect 315868 158672 315915 158676
rect 318558 158674 318564 158676
rect 315910 158616 315915 158672
rect 315798 158612 315804 158614
rect 315868 158612 315915 158616
rect 318518 158614 318564 158674
rect 318628 158672 318675 158676
rect 320950 158674 320956 158676
rect 318670 158616 318675 158672
rect 318558 158612 318564 158614
rect 318628 158612 318675 158616
rect 320910 158614 320956 158674
rect 321020 158672 321067 158676
rect 323342 158674 323348 158676
rect 321062 158616 321067 158672
rect 320950 158612 320956 158614
rect 321020 158612 321067 158616
rect 323302 158614 323348 158674
rect 323412 158672 323459 158676
rect 325918 158674 325924 158676
rect 323454 158616 323459 158672
rect 323342 158612 323348 158614
rect 323412 158612 323459 158616
rect 325878 158614 325924 158674
rect 325988 158672 326035 158676
rect 326030 158616 326035 158672
rect 325918 158612 325924 158614
rect 325988 158612 326035 158616
rect 313457 158611 313523 158612
rect 315849 158611 315915 158612
rect 318609 158611 318675 158612
rect 321001 158611 321067 158612
rect 323393 158611 323459 158612
rect 325969 158611 326035 158612
rect 219014 158476 219020 158540
rect 219084 158538 219090 158540
rect 224953 158538 225019 158541
rect 219084 158536 225019 158538
rect 219084 158480 224958 158536
rect 225014 158480 225019 158536
rect 219084 158478 225019 158480
rect 219084 158476 219090 158478
rect 224953 158475 225019 158478
rect 241830 158476 241836 158540
rect 241900 158538 241906 158540
rect 374269 158538 374335 158541
rect 241900 158536 374335 158538
rect 241900 158480 374274 158536
rect 374330 158480 374335 158536
rect 241900 158478 374335 158480
rect 241900 158476 241906 158478
rect 374269 158475 374335 158478
rect 216254 158340 216260 158404
rect 216324 158402 216330 158404
rect 223573 158402 223639 158405
rect 216324 158400 223639 158402
rect 216324 158344 223578 158400
rect 223634 158344 223639 158400
rect 216324 158342 223639 158344
rect 216324 158340 216330 158342
rect 223573 158339 223639 158342
rect 273294 158340 273300 158404
rect 273364 158402 273370 158404
rect 274449 158402 274515 158405
rect 276105 158404 276171 158405
rect 276054 158402 276060 158404
rect 273364 158400 274515 158402
rect 273364 158344 274454 158400
rect 274510 158344 274515 158400
rect 273364 158342 274515 158344
rect 276014 158342 276060 158402
rect 276124 158400 276171 158404
rect 276166 158344 276171 158400
rect 273364 158340 273370 158342
rect 274449 158339 274515 158342
rect 276054 158340 276060 158342
rect 276124 158340 276171 158344
rect 281022 158340 281028 158404
rect 281092 158402 281098 158404
rect 281349 158402 281415 158405
rect 281092 158400 281415 158402
rect 281092 158344 281354 158400
rect 281410 158344 281415 158400
rect 281092 158342 281415 158344
rect 281092 158340 281098 158342
rect 276105 158339 276171 158340
rect 281349 158339 281415 158342
rect 285990 158340 285996 158404
rect 286060 158402 286066 158404
rect 286317 158402 286383 158405
rect 286060 158400 286383 158402
rect 286060 158344 286322 158400
rect 286378 158344 286383 158400
rect 286060 158342 286383 158344
rect 286060 158340 286066 158342
rect 286317 158339 286383 158342
rect 293534 158340 293540 158404
rect 293604 158402 293610 158404
rect 293677 158402 293743 158405
rect 293604 158400 293743 158402
rect 293604 158344 293682 158400
rect 293738 158344 293743 158400
rect 293604 158342 293743 158344
rect 293604 158340 293610 158342
rect 293677 158339 293743 158342
rect 218881 158266 218947 158269
rect 227713 158266 227779 158269
rect 267641 158268 267707 158269
rect 311065 158268 311131 158269
rect 267590 158266 267596 158268
rect 218881 158264 227779 158266
rect 218881 158208 218886 158264
rect 218942 158208 227718 158264
rect 227774 158208 227779 158264
rect 218881 158206 227779 158208
rect 267550 158206 267596 158266
rect 267660 158264 267707 158268
rect 311014 158266 311020 158268
rect 267702 158208 267707 158264
rect 218881 158203 218947 158206
rect 227713 158203 227779 158206
rect 267590 158204 267596 158206
rect 267660 158204 267707 158208
rect 310974 158206 311020 158266
rect 311084 158264 311131 158268
rect 311126 158208 311131 158264
rect 311014 158204 311020 158206
rect 311084 158204 311131 158208
rect 267641 158203 267707 158204
rect 311065 158203 311131 158204
rect 354121 158266 354187 158269
rect 365161 158266 365227 158269
rect 354121 158264 365227 158266
rect 354121 158208 354126 158264
rect 354182 158208 365166 158264
rect 365222 158208 365227 158264
rect 354121 158206 365227 158208
rect 354121 158203 354187 158206
rect 365161 158203 365227 158206
rect 217174 158068 217180 158132
rect 217244 158130 217250 158132
rect 231853 158130 231919 158133
rect 217244 158128 231919 158130
rect 217244 158072 231858 158128
rect 231914 158072 231919 158128
rect 217244 158070 231919 158072
rect 217244 158068 217250 158070
rect 231853 158067 231919 158070
rect 246614 158068 246620 158132
rect 246684 158130 246690 158132
rect 246849 158130 246915 158133
rect 246684 158128 246915 158130
rect 246684 158072 246854 158128
rect 246910 158072 246915 158128
rect 246684 158070 246915 158072
rect 246684 158068 246690 158070
rect 246849 158067 246915 158070
rect 353937 158130 354003 158133
rect 369209 158130 369275 158133
rect 353937 158128 369275 158130
rect 353937 158072 353942 158128
rect 353998 158072 369214 158128
rect 369270 158072 369275 158128
rect 353937 158070 369275 158072
rect 353937 158067 354003 158070
rect 369209 158067 369275 158070
rect 217358 157932 217364 157996
rect 217428 157994 217434 157996
rect 238753 157994 238819 157997
rect 248689 157996 248755 157997
rect 248638 157994 248644 157996
rect 217428 157992 238819 157994
rect 217428 157936 238758 157992
rect 238814 157936 238819 157992
rect 217428 157934 238819 157936
rect 248598 157934 248644 157994
rect 248708 157992 248755 157996
rect 248750 157936 248755 157992
rect 217428 157932 217434 157934
rect 238753 157931 238819 157934
rect 248638 157932 248644 157934
rect 248708 157932 248755 157936
rect 251398 157932 251404 157996
rect 251468 157994 251474 157996
rect 252277 157994 252343 157997
rect 251468 157992 252343 157994
rect 251468 157936 252282 157992
rect 252338 157936 252343 157992
rect 251468 157934 252343 157936
rect 251468 157932 251474 157934
rect 248689 157931 248755 157932
rect 252277 157931 252343 157934
rect 253422 157932 253428 157996
rect 253492 157994 253498 157996
rect 253565 157994 253631 157997
rect 260649 157996 260715 157997
rect 260598 157994 260604 157996
rect 253492 157992 253631 157994
rect 253492 157936 253570 157992
rect 253626 157936 253631 157992
rect 253492 157934 253631 157936
rect 260558 157934 260604 157994
rect 260668 157992 260715 157996
rect 260710 157936 260715 157992
rect 253492 157932 253498 157934
rect 253565 157931 253631 157934
rect 260598 157932 260604 157934
rect 260668 157932 260715 157936
rect 260649 157931 260715 157932
rect 299473 157994 299539 157997
rect 363689 157994 363755 157997
rect 299473 157992 363755 157994
rect 299473 157936 299478 157992
rect 299534 157936 363694 157992
rect 363750 157936 363755 157992
rect 299473 157934 363755 157936
rect 299473 157931 299539 157934
rect 363689 157931 363755 157934
rect 214741 157858 214807 157861
rect 219433 157858 219499 157861
rect 261753 157860 261819 157861
rect 261702 157858 261708 157860
rect 214741 157856 219499 157858
rect 214741 157800 214746 157856
rect 214802 157800 219438 157856
rect 219494 157800 219499 157856
rect 214741 157798 219499 157800
rect 261662 157798 261708 157858
rect 261772 157856 261819 157860
rect 261814 157800 261819 157856
rect 214741 157795 214807 157798
rect 219433 157795 219499 157798
rect 261702 157796 261708 157798
rect 261772 157796 261819 157800
rect 263910 157796 263916 157860
rect 263980 157858 263986 157860
rect 264513 157858 264579 157861
rect 263980 157856 264579 157858
rect 263980 157800 264518 157856
rect 264574 157800 264579 157856
rect 263980 157798 264579 157800
rect 263980 157796 263986 157798
rect 261753 157795 261819 157796
rect 264513 157795 264579 157798
rect 266486 157796 266492 157860
rect 266556 157858 266562 157860
rect 266905 157858 266971 157861
rect 266556 157856 266971 157858
rect 266556 157800 266910 157856
rect 266966 157800 266971 157856
rect 266556 157798 266971 157800
rect 266556 157796 266562 157798
rect 266905 157795 266971 157798
rect 268326 157796 268332 157860
rect 268396 157858 268402 157860
rect 268929 157858 268995 157861
rect 268396 157856 268995 157858
rect 268396 157800 268934 157856
rect 268990 157800 268995 157856
rect 268396 157798 268995 157800
rect 268396 157796 268402 157798
rect 268929 157795 268995 157798
rect 265382 157660 265388 157724
rect 265452 157722 265458 157724
rect 265985 157722 266051 157725
rect 265452 157720 266051 157722
rect 265452 157664 265990 157720
rect 266046 157664 266051 157720
rect 265452 157662 266051 157664
rect 265452 157660 265458 157662
rect 265985 157659 266051 157662
rect 273662 157660 273668 157724
rect 273732 157722 273738 157724
rect 274541 157722 274607 157725
rect 273732 157720 274607 157722
rect 273732 157664 274546 157720
rect 274602 157664 274607 157720
rect 273732 157662 274607 157664
rect 273732 157660 273738 157662
rect 274541 157659 274607 157662
rect 278446 157660 278452 157724
rect 278516 157722 278522 157724
rect 278681 157722 278747 157725
rect 278516 157720 278747 157722
rect 278516 157664 278686 157720
rect 278742 157664 278747 157720
rect 278516 157662 278747 157664
rect 278516 157660 278522 157662
rect 278681 157659 278747 157662
rect 283598 157524 283604 157588
rect 283668 157586 283674 157588
rect 283925 157586 283991 157589
rect 291009 157588 291075 157589
rect 290958 157586 290964 157588
rect 283668 157584 283991 157586
rect 283668 157528 283930 157584
rect 283986 157528 283991 157584
rect 283668 157526 283991 157528
rect 290918 157526 290964 157586
rect 291028 157584 291075 157588
rect 291070 157528 291075 157584
rect 283668 157524 283674 157526
rect 283925 157523 283991 157526
rect 290958 157524 290964 157526
rect 291028 157524 291075 157528
rect 291009 157523 291075 157524
rect 253657 157452 253723 157453
rect 256233 157452 256299 157453
rect 244222 157388 244228 157452
rect 244292 157450 244298 157452
rect 244292 157390 244474 157450
rect 244292 157388 244298 157390
rect 244414 157178 244474 157390
rect 245510 157388 245516 157452
rect 245580 157388 245586 157452
rect 253606 157450 253612 157452
rect 253566 157390 253612 157450
rect 253676 157448 253723 157452
rect 256182 157450 256188 157452
rect 253718 157392 253723 157448
rect 253606 157388 253612 157390
rect 253676 157388 253723 157392
rect 256142 157390 256188 157450
rect 256252 157448 256299 157452
rect 256294 157392 256299 157448
rect 256182 157388 256188 157390
rect 256252 157388 256299 157392
rect 363270 157388 363276 157452
rect 363340 157450 363346 157452
rect 363781 157450 363847 157453
rect 363340 157448 363847 157450
rect 363340 157392 363786 157448
rect 363842 157392 363847 157448
rect 363340 157390 363847 157392
rect 363340 157388 363346 157390
rect 245518 157314 245578 157388
rect 253657 157387 253723 157388
rect 256233 157387 256299 157388
rect 363781 157387 363847 157390
rect 370129 157314 370195 157317
rect 245518 157312 370195 157314
rect 245518 157256 370134 157312
rect 370190 157256 370195 157312
rect 245518 157254 370195 157256
rect 370129 157251 370195 157254
rect 367645 157178 367711 157181
rect 244414 157176 367711 157178
rect 244414 157120 367650 157176
rect 367706 157120 367711 157176
rect 244414 157118 367711 157120
rect 367645 157115 367711 157118
rect 247718 156980 247724 157044
rect 247788 157042 247794 157044
rect 370313 157042 370379 157045
rect 247788 157040 370379 157042
rect 247788 156984 370318 157040
rect 370374 156984 370379 157040
rect 247788 156982 370379 156984
rect 247788 156980 247794 156982
rect 370313 156979 370379 156982
rect 352557 156906 352623 156909
rect 356789 156906 356855 156909
rect 352557 156904 356855 156906
rect 352557 156848 352562 156904
rect 352618 156848 356794 156904
rect 356850 156848 356855 156904
rect 352557 156846 356855 156848
rect 352557 156843 352623 156846
rect 356789 156843 356855 156846
rect 348417 156770 348483 156773
rect 362401 156770 362467 156773
rect 348417 156768 362467 156770
rect 348417 156712 348422 156768
rect 348478 156712 362406 156768
rect 362462 156712 362467 156768
rect 348417 156710 362467 156712
rect 348417 156707 348483 156710
rect 362401 156707 362467 156710
rect 345657 156634 345723 156637
rect 359641 156634 359707 156637
rect 345657 156632 359707 156634
rect 345657 156576 345662 156632
rect 345718 156576 359646 156632
rect 359702 156576 359707 156632
rect 345657 156574 359707 156576
rect 345657 156571 345723 156574
rect 359641 156571 359707 156574
rect 246849 155954 246915 155957
rect 368657 155954 368723 155957
rect 246849 155952 368723 155954
rect 246849 155896 246854 155952
rect 246910 155896 368662 155952
rect 368718 155896 368723 155952
rect 246849 155894 368723 155896
rect 246849 155891 246915 155894
rect 368657 155891 368723 155894
rect 216990 155484 216996 155548
rect 217060 155546 217066 155548
rect 251265 155546 251331 155549
rect 217060 155544 251331 155546
rect 217060 155488 251270 155544
rect 251326 155488 251331 155544
rect 217060 155486 251331 155488
rect 217060 155484 217066 155486
rect 251265 155483 251331 155486
rect 210969 155410 211035 155413
rect 269113 155410 269179 155413
rect 210969 155408 269179 155410
rect 210969 155352 210974 155408
rect 211030 155352 269118 155408
rect 269174 155352 269179 155408
rect 210969 155350 269179 155352
rect 210969 155347 211035 155350
rect 269113 155347 269179 155350
rect 210785 155274 210851 155277
rect 270493 155274 270559 155277
rect 210785 155272 270559 155274
rect 210785 155216 210790 155272
rect 210846 155216 270498 155272
rect 270554 155216 270559 155272
rect 210785 155214 270559 155216
rect 210785 155211 210851 155214
rect 270493 155211 270559 155214
rect 292573 153778 292639 153781
rect 368606 153778 368612 153780
rect 292573 153776 368612 153778
rect 292573 153720 292578 153776
rect 292634 153720 368612 153776
rect 292573 153718 368612 153720
rect 292573 153715 292639 153718
rect 368606 153716 368612 153718
rect 368676 153716 368682 153780
rect 580717 152690 580783 152693
rect 583520 152690 584960 152780
rect 580717 152688 584960 152690
rect 580717 152632 580722 152688
rect 580778 152632 584960 152688
rect 580717 152630 584960 152632
rect 580717 152627 580783 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580625 139362 580691 139365
rect 583520 139362 584960 139452
rect 580625 139360 584960 139362
rect 580625 139304 580630 139360
rect 580686 139304 584960 139360
rect 580625 139302 584960 139304
rect 580625 139299 580691 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 368974 125564 368980 125628
rect 369044 125626 369050 125628
rect 583526 125626 583586 125838
rect 369044 125566 583586 125626
rect 369044 125564 369050 125566
rect -960 123572 480 123812
rect 580533 112842 580599 112845
rect 583520 112842 584960 112932
rect 580533 112840 584960 112842
rect 580533 112784 580538 112840
rect 580594 112784 584960 112840
rect 580533 112782 584960 112784
rect 580533 112779 580599 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 365110 99452 365116 99516
rect 365180 99514 365186 99516
rect 583520 99514 584960 99604
rect 365180 99454 584960 99514
rect 365180 99452 365186 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 367686 85580 367692 85644
rect 367756 85642 367762 85644
rect 583526 85642 583586 85990
rect 367756 85582 583586 85642
rect 367756 85580 367762 85582
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580441 72994 580507 72997
rect 583520 72994 584960 73084
rect 580441 72992 584960 72994
rect 580441 72936 580446 72992
rect 580502 72936 584960 72992
rect 580441 72934 584960 72936
rect 580441 72931 580507 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 364926 45596 364932 45660
rect 364996 45658 365002 45660
rect 583526 45658 583586 46142
rect 364996 45598 583586 45658
rect 364996 45596 365002 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 351637 6762 351703 6765
rect 361573 6762 361639 6765
rect 351637 6760 361639 6762
rect 351637 6704 351642 6760
rect 351698 6704 361578 6760
rect 361634 6704 361639 6760
rect 351637 6702 361639 6704
rect 351637 6699 351703 6702
rect 361573 6699 361639 6702
rect 348049 6626 348115 6629
rect 364558 6626 364564 6628
rect 348049 6624 364564 6626
rect -960 6490 480 6580
rect 348049 6568 348054 6624
rect 348110 6568 364564 6624
rect 348049 6566 364564 6568
rect 348049 6563 348115 6566
rect 364558 6564 364564 6566
rect 364628 6564 364634 6628
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 326797 6490 326863 6493
rect 359038 6490 359044 6492
rect 326797 6488 359044 6490
rect 326797 6432 326802 6488
rect 326858 6432 359044 6488
rect 326797 6430 359044 6432
rect 326797 6427 326863 6430
rect 359038 6428 359044 6430
rect 359108 6428 359114 6492
rect 583520 6476 584960 6566
rect 323301 6354 323367 6357
rect 358302 6354 358308 6356
rect 323301 6352 358308 6354
rect 323301 6296 323306 6352
rect 323362 6296 358308 6352
rect 323301 6294 358308 6296
rect 323301 6291 323367 6294
rect 358302 6292 358308 6294
rect 358372 6292 358378 6356
rect 320909 6218 320975 6221
rect 367318 6218 367324 6220
rect 320909 6216 367324 6218
rect 320909 6160 320914 6216
rect 320970 6160 367324 6216
rect 320909 6158 367324 6160
rect 320909 6155 320975 6158
rect 367318 6156 367324 6158
rect 367388 6156 367394 6220
rect 335077 4042 335143 4045
rect 359406 4042 359412 4044
rect 335077 4040 359412 4042
rect 335077 3984 335082 4040
rect 335138 3984 359412 4040
rect 335077 3982 359412 3984
rect 335077 3979 335143 3982
rect 359406 3980 359412 3982
rect 359476 3980 359482 4044
rect 331581 3906 331647 3909
rect 360142 3906 360148 3908
rect 331581 3904 360148 3906
rect 331581 3848 331586 3904
rect 331642 3848 360148 3904
rect 331581 3846 360148 3848
rect 331581 3843 331647 3846
rect 360142 3844 360148 3846
rect 360212 3844 360218 3908
rect 327993 3770 328059 3773
rect 355961 3770 356027 3773
rect 358118 3770 358124 3772
rect 327993 3768 356027 3770
rect 327993 3712 327998 3768
rect 328054 3712 355966 3768
rect 356022 3712 356027 3768
rect 327993 3710 356027 3712
rect 327993 3707 328059 3710
rect 355961 3707 356027 3710
rect 356102 3710 358124 3770
rect 212165 3634 212231 3637
rect 215886 3634 215892 3636
rect 212165 3632 215892 3634
rect 212165 3576 212170 3632
rect 212226 3576 215892 3632
rect 212165 3574 215892 3576
rect 212165 3571 212231 3574
rect 215886 3572 215892 3574
rect 215956 3572 215962 3636
rect 218053 3634 218119 3637
rect 219198 3634 219204 3636
rect 218053 3632 219204 3634
rect 218053 3576 218058 3632
rect 218114 3576 219204 3632
rect 218053 3574 219204 3576
rect 218053 3571 218119 3574
rect 219198 3572 219204 3574
rect 219268 3572 219274 3636
rect 325601 3634 325667 3637
rect 356102 3634 356162 3710
rect 358118 3708 358124 3710
rect 358188 3708 358194 3772
rect 325601 3632 356162 3634
rect 325601 3576 325606 3632
rect 325662 3576 356162 3632
rect 325601 3574 356162 3576
rect 356329 3634 356395 3637
rect 360694 3634 360700 3636
rect 356329 3632 360700 3634
rect 356329 3576 356334 3632
rect 356390 3576 360700 3632
rect 356329 3574 360700 3576
rect 325601 3571 325667 3574
rect 356329 3571 356395 3574
rect 360694 3572 360700 3574
rect 360764 3572 360770 3636
rect 365846 3572 365852 3636
rect 365916 3634 365922 3636
rect 367001 3634 367067 3637
rect 365916 3632 367067 3634
rect 365916 3576 367006 3632
rect 367062 3576 367067 3632
rect 365916 3574 367067 3576
rect 365916 3572 365922 3574
rect 367001 3571 367067 3574
rect 214465 3498 214531 3501
rect 215150 3498 215156 3500
rect 214465 3496 215156 3498
rect 214465 3440 214470 3496
rect 214526 3440 215156 3496
rect 214465 3438 215156 3440
rect 214465 3435 214531 3438
rect 215150 3436 215156 3438
rect 215220 3436 215226 3500
rect 215661 3498 215727 3501
rect 216438 3498 216444 3500
rect 215661 3496 216444 3498
rect 215661 3440 215666 3496
rect 215722 3440 216444 3496
rect 215661 3438 216444 3440
rect 215661 3435 215727 3438
rect 216438 3436 216444 3438
rect 216508 3436 216514 3500
rect 216857 3498 216923 3501
rect 217542 3498 217548 3500
rect 216857 3496 217548 3498
rect 216857 3440 216862 3496
rect 216918 3440 217548 3496
rect 216857 3438 217548 3440
rect 216857 3435 216923 3438
rect 217542 3436 217548 3438
rect 217612 3436 217618 3500
rect 218646 3436 218652 3500
rect 218716 3498 218722 3500
rect 219249 3498 219315 3501
rect 218716 3496 219315 3498
rect 218716 3440 219254 3496
rect 219310 3440 219315 3496
rect 218716 3438 219315 3440
rect 218716 3436 218722 3438
rect 219249 3435 219315 3438
rect 324405 3498 324471 3501
rect 324405 3496 357082 3498
rect 324405 3440 324410 3496
rect 324466 3440 357082 3496
rect 324405 3438 357082 3440
rect 324405 3435 324471 3438
rect 205081 3362 205147 3365
rect 214414 3362 214420 3364
rect 205081 3360 214420 3362
rect 205081 3304 205086 3360
rect 205142 3304 214420 3360
rect 205081 3302 214420 3304
rect 205081 3299 205147 3302
rect 214414 3300 214420 3302
rect 214484 3300 214490 3364
rect 290181 3362 290247 3365
rect 356830 3362 356836 3364
rect 290181 3360 356836 3362
rect 290181 3304 290186 3360
rect 290242 3304 356836 3360
rect 290181 3302 356836 3304
rect 290181 3299 290247 3302
rect 356830 3300 356836 3302
rect 356900 3300 356906 3364
rect 357022 3362 357082 3438
rect 358486 3436 358492 3500
rect 358556 3498 358562 3500
rect 358721 3498 358787 3501
rect 358556 3496 358787 3498
rect 358556 3440 358726 3496
rect 358782 3440 358787 3496
rect 358556 3438 358787 3440
rect 358556 3436 358562 3438
rect 358721 3435 358787 3438
rect 358854 3436 358860 3500
rect 358924 3498 358930 3500
rect 359917 3498 359983 3501
rect 358924 3496 359983 3498
rect 358924 3440 359922 3496
rect 359978 3440 359983 3496
rect 358924 3438 359983 3440
rect 358924 3436 358930 3438
rect 359917 3435 359983 3438
rect 360326 3436 360332 3500
rect 360396 3498 360402 3500
rect 361113 3498 361179 3501
rect 360396 3496 361179 3498
rect 360396 3440 361118 3496
rect 361174 3440 361179 3496
rect 360396 3438 361179 3440
rect 360396 3436 360402 3438
rect 361113 3435 361179 3438
rect 361614 3436 361620 3500
rect 361684 3498 361690 3500
rect 362309 3498 362375 3501
rect 361684 3496 362375 3498
rect 361684 3440 362314 3496
rect 362370 3440 362375 3496
rect 361684 3438 362375 3440
rect 361684 3436 361690 3438
rect 362309 3435 362375 3438
rect 362902 3436 362908 3500
rect 362972 3498 362978 3500
rect 363505 3498 363571 3501
rect 362972 3496 363571 3498
rect 362972 3440 363510 3496
rect 363566 3440 363571 3496
rect 362972 3438 363571 3440
rect 362972 3436 362978 3438
rect 363505 3435 363571 3438
rect 364374 3436 364380 3500
rect 364444 3498 364450 3500
rect 364609 3498 364675 3501
rect 364444 3496 364675 3498
rect 364444 3440 364614 3496
rect 364670 3440 364675 3496
rect 364444 3438 364675 3440
rect 364444 3436 364450 3438
rect 364609 3435 364675 3438
rect 365662 3436 365668 3500
rect 365732 3498 365738 3500
rect 365805 3498 365871 3501
rect 365732 3496 365871 3498
rect 365732 3440 365810 3496
rect 365866 3440 365871 3496
rect 365732 3438 365871 3440
rect 365732 3436 365738 3438
rect 365805 3435 365871 3438
rect 367134 3436 367140 3500
rect 367204 3498 367210 3500
rect 368197 3498 368263 3501
rect 367204 3496 368263 3498
rect 367204 3440 368202 3496
rect 368258 3440 368263 3496
rect 367204 3438 368263 3440
rect 367204 3436 367210 3438
rect 368197 3435 368263 3438
rect 368422 3436 368428 3500
rect 368492 3498 368498 3500
rect 369393 3498 369459 3501
rect 368492 3496 369459 3498
rect 368492 3440 369398 3496
rect 369454 3440 369459 3496
rect 368492 3438 369459 3440
rect 368492 3436 368498 3438
rect 369393 3435 369459 3438
rect 369894 3436 369900 3500
rect 369964 3498 369970 3500
rect 370589 3498 370655 3501
rect 369964 3496 370655 3498
rect 369964 3440 370594 3496
rect 370650 3440 370655 3496
rect 369964 3438 370655 3440
rect 369964 3436 369970 3438
rect 370589 3435 370655 3438
rect 359222 3362 359228 3364
rect 357022 3302 359228 3362
rect 359222 3300 359228 3302
rect 359292 3300 359298 3364
rect 369158 3300 369164 3364
rect 369228 3362 369234 3364
rect 379973 3362 380039 3365
rect 369228 3360 380039 3362
rect 369228 3304 379978 3360
rect 380034 3304 380039 3360
rect 369228 3302 380039 3304
rect 369228 3300 369234 3302
rect 379973 3299 380039 3302
rect 339861 3226 339927 3229
rect 355961 3226 356027 3229
rect 360510 3226 360516 3228
rect 339861 3224 354690 3226
rect 339861 3168 339866 3224
rect 339922 3168 354690 3224
rect 339861 3166 354690 3168
rect 339861 3163 339927 3166
rect 354630 3090 354690 3166
rect 355961 3224 360516 3226
rect 355961 3168 355966 3224
rect 356022 3168 360516 3224
rect 355961 3166 360516 3168
rect 355961 3163 356027 3166
rect 360510 3164 360516 3166
rect 360580 3164 360586 3228
rect 363086 3090 363092 3092
rect 354630 3030 363092 3090
rect 363086 3028 363092 3030
rect 363156 3028 363162 3092
<< via3 >>
rect 238340 477260 238404 477324
rect 241836 477124 241900 477188
rect 256188 476988 256252 477052
rect 239628 476852 239692 476916
rect 240548 476852 240612 476916
rect 236132 476716 236196 476780
rect 258028 476716 258092 476780
rect 263548 476716 263612 476780
rect 308628 476716 308692 476780
rect 313412 476716 313476 476780
rect 265940 476580 266004 476644
rect 270908 476580 270972 476644
rect 253428 476444 253492 476508
rect 261156 476444 261220 476508
rect 274404 476504 274468 476508
rect 274404 476448 274454 476504
rect 274454 476448 274468 476504
rect 274404 476444 274468 476448
rect 318564 476444 318628 476508
rect 325924 476444 325988 476508
rect 244228 476308 244292 476372
rect 247724 476308 247788 476372
rect 250116 476308 250180 476372
rect 251404 476308 251468 476372
rect 259500 476308 259564 476372
rect 266492 476308 266556 476372
rect 268332 476308 268396 476372
rect 273668 476308 273732 476372
rect 276060 476308 276124 476372
rect 278084 476308 278148 476372
rect 311020 476308 311084 476372
rect 237236 476232 237300 476236
rect 237236 476176 237250 476232
rect 237250 476176 237300 476232
rect 237236 476172 237300 476176
rect 243124 476172 243188 476236
rect 245516 476232 245580 476236
rect 245516 476176 245566 476232
rect 245566 476176 245580 476232
rect 245516 476172 245580 476176
rect 246620 476172 246684 476236
rect 248276 476232 248340 476236
rect 248276 476176 248290 476232
rect 248290 476176 248340 476232
rect 248276 476172 248340 476176
rect 248644 476172 248708 476236
rect 250852 476172 250916 476236
rect 252324 476172 252388 476236
rect 253612 476172 253676 476236
rect 254532 476172 254596 476236
rect 255820 476172 255884 476236
rect 257108 476172 257172 476236
rect 258580 476172 258644 476236
rect 260604 476232 260668 476236
rect 260604 476176 260654 476232
rect 260654 476176 260668 476232
rect 260604 476172 260668 476176
rect 261708 476172 261772 476236
rect 262812 476172 262876 476236
rect 263916 476172 263980 476236
rect 265388 476172 265452 476236
rect 267596 476232 267660 476236
rect 267596 476176 267610 476232
rect 267610 476176 267660 476232
rect 267596 476172 267660 476176
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 273300 476172 273364 476236
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278452 476172 278516 476236
rect 279188 476172 279252 476236
rect 281028 476172 281092 476236
rect 283604 476172 283668 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293540 476172 293604 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476172 300964 476236
rect 303476 476232 303540 476236
rect 303476 476176 303526 476232
rect 303526 476176 303540 476232
rect 303476 476172 303540 476176
rect 306052 476172 306116 476236
rect 315804 476172 315868 476236
rect 320956 476172 321020 476236
rect 323348 476172 323412 476236
rect 367876 445844 367940 445908
rect 365116 445708 365180 445772
rect 214604 444756 214668 444820
rect 364932 444620 364996 444684
rect 368980 444484 369044 444548
rect 367692 444348 367756 444412
rect 216076 441628 216140 441692
rect 232084 374036 232148 374100
rect 232084 372676 232148 372740
rect 232820 310660 232884 310724
rect 232820 310388 232884 310452
rect 232636 309708 232700 309772
rect 232452 308620 232516 308684
rect 169340 308484 169404 308548
rect 359964 308484 360028 308548
rect 358124 306444 358188 306508
rect 218836 306036 218900 306100
rect 367140 306036 367204 306100
rect 219020 305900 219084 305964
rect 217180 305764 217244 305828
rect 217364 305628 217428 305692
rect 358124 304268 358188 304332
rect 369900 303452 369964 303516
rect 215156 303180 215220 303244
rect 216260 303044 216324 303108
rect 219204 301684 219268 301748
rect 169708 301548 169772 301612
rect 216996 301412 217060 301476
rect 169156 301140 169220 301204
rect 368612 300052 368676 300116
rect 169340 299100 169404 299164
rect 169156 297876 169220 297940
rect 169708 297740 169772 297804
rect 214420 284820 214484 284884
rect 368428 280740 368492 280804
rect 215892 269724 215956 269788
rect 369164 265508 369228 265572
rect 361620 260204 361684 260268
rect 365668 260068 365732 260132
rect 216444 254492 216508 254556
rect 364380 254492 364444 254556
rect 365852 251772 365916 251836
rect 358860 250956 358924 251020
rect 362908 250820 362972 250884
rect 359044 250684 359108 250748
rect 358308 250548 358372 250612
rect 217548 250412 217612 250476
rect 364564 250412 364628 250476
rect 360332 248100 360396 248164
rect 358124 247964 358188 248028
rect 363276 247828 363340 247892
rect 363460 247692 363524 247756
rect 363092 247556 363156 247620
rect 360700 245516 360764 245580
rect 359412 245380 359476 245444
rect 362540 245244 362604 245308
rect 359228 245108 359292 245172
rect 360516 244972 360580 245036
rect 367324 244836 367388 244900
rect 358492 244700 358556 244764
rect 218652 243476 218716 243540
rect 357572 243476 357636 243540
rect 216076 187716 216140 187780
rect 367876 178060 367940 178124
rect 214604 162828 214668 162892
rect 356836 160108 356900 160172
rect 363460 160108 363524 160172
rect 278078 159896 278142 159900
rect 278078 159840 278134 159896
rect 278134 159840 278142 159896
rect 278078 159836 278142 159840
rect 300926 159760 300990 159764
rect 300926 159704 300950 159760
rect 300950 159704 300990 159760
rect 300926 159700 300990 159704
rect 258494 159564 258558 159628
rect 271006 159624 271070 159628
rect 271006 159568 271050 159624
rect 271050 159568 271070 159624
rect 271006 159564 271070 159568
rect 275766 159564 275830 159628
rect 279166 159564 279230 159628
rect 288278 159564 288342 159628
rect 295894 159624 295958 159628
rect 295894 159568 295946 159624
rect 295946 159568 295958 159624
rect 295894 159564 295958 159568
rect 265940 159428 266004 159492
rect 250852 159156 250916 159220
rect 243124 159020 243188 159084
rect 236132 158884 236196 158948
rect 357572 158884 357636 158948
rect 362540 158944 362604 158948
rect 362540 158888 362554 158944
rect 362554 158888 362604 158944
rect 362540 158884 362604 158888
rect 237236 158748 237300 158812
rect 218836 158612 218900 158676
rect 238156 158672 238220 158676
rect 238156 158616 238170 158672
rect 238170 158616 238220 158672
rect 238156 158612 238220 158616
rect 239628 158672 239692 158676
rect 239628 158616 239642 158672
rect 239642 158616 239692 158672
rect 239628 158612 239692 158616
rect 240548 158612 240612 158676
rect 248276 158672 248340 158676
rect 248276 158616 248326 158672
rect 248326 158616 248340 158672
rect 248276 158612 248340 158616
rect 250116 158612 250180 158676
rect 252324 158672 252388 158676
rect 252324 158616 252374 158672
rect 252374 158616 252388 158672
rect 252324 158612 252388 158616
rect 254532 158612 254596 158676
rect 255820 158672 255884 158676
rect 255820 158616 255870 158672
rect 255870 158616 255884 158672
rect 255820 158612 255884 158616
rect 257108 158612 257172 158676
rect 258212 158612 258276 158676
rect 259500 158672 259564 158676
rect 259500 158616 259550 158672
rect 259550 158616 259564 158672
rect 259500 158612 259564 158616
rect 261156 158612 261220 158676
rect 262812 158672 262876 158676
rect 262812 158616 262862 158672
rect 262862 158616 262876 158672
rect 262812 158612 262876 158616
rect 263548 158672 263612 158676
rect 263548 158616 263598 158672
rect 263598 158616 263612 158672
rect 263548 158612 263612 158616
rect 268700 158672 268764 158676
rect 268700 158616 268750 158672
rect 268750 158616 268764 158672
rect 268700 158612 268764 158616
rect 269804 158672 269868 158676
rect 269804 158616 269854 158672
rect 269854 158616 269868 158672
rect 269804 158612 269868 158616
rect 271092 158672 271156 158676
rect 271092 158616 271142 158672
rect 271142 158616 271156 158672
rect 271092 158612 271156 158616
rect 272196 158672 272260 158676
rect 272196 158616 272246 158672
rect 272246 158616 272260 158672
rect 272196 158612 272260 158616
rect 274404 158672 274468 158676
rect 274404 158616 274454 158672
rect 274454 158616 274468 158672
rect 274404 158612 274468 158616
rect 276980 158672 277044 158676
rect 276980 158616 277030 158672
rect 277030 158616 277044 158672
rect 276980 158612 277044 158616
rect 298508 158672 298572 158676
rect 298508 158616 298558 158672
rect 298558 158616 298572 158672
rect 298508 158612 298572 158616
rect 303476 158672 303540 158676
rect 303476 158616 303526 158672
rect 303526 158616 303540 158672
rect 303476 158612 303540 158616
rect 306052 158672 306116 158676
rect 306052 158616 306102 158672
rect 306102 158616 306116 158672
rect 306052 158612 306116 158616
rect 308628 158612 308692 158676
rect 313412 158672 313476 158676
rect 313412 158616 313462 158672
rect 313462 158616 313476 158672
rect 313412 158612 313476 158616
rect 315804 158672 315868 158676
rect 315804 158616 315854 158672
rect 315854 158616 315868 158672
rect 315804 158612 315868 158616
rect 318564 158672 318628 158676
rect 318564 158616 318614 158672
rect 318614 158616 318628 158672
rect 318564 158612 318628 158616
rect 320956 158672 321020 158676
rect 320956 158616 321006 158672
rect 321006 158616 321020 158672
rect 320956 158612 321020 158616
rect 323348 158672 323412 158676
rect 323348 158616 323398 158672
rect 323398 158616 323412 158672
rect 323348 158612 323412 158616
rect 325924 158672 325988 158676
rect 325924 158616 325974 158672
rect 325974 158616 325988 158672
rect 325924 158612 325988 158616
rect 219020 158476 219084 158540
rect 241836 158476 241900 158540
rect 216260 158340 216324 158404
rect 273300 158340 273364 158404
rect 276060 158400 276124 158404
rect 276060 158344 276110 158400
rect 276110 158344 276124 158400
rect 276060 158340 276124 158344
rect 281028 158340 281092 158404
rect 285996 158340 286060 158404
rect 293540 158340 293604 158404
rect 267596 158264 267660 158268
rect 267596 158208 267646 158264
rect 267646 158208 267660 158264
rect 267596 158204 267660 158208
rect 311020 158264 311084 158268
rect 311020 158208 311070 158264
rect 311070 158208 311084 158264
rect 311020 158204 311084 158208
rect 217180 158068 217244 158132
rect 246620 158068 246684 158132
rect 217364 157932 217428 157996
rect 248644 157992 248708 157996
rect 248644 157936 248694 157992
rect 248694 157936 248708 157992
rect 248644 157932 248708 157936
rect 251404 157932 251468 157996
rect 253428 157932 253492 157996
rect 260604 157992 260668 157996
rect 260604 157936 260654 157992
rect 260654 157936 260668 157992
rect 260604 157932 260668 157936
rect 261708 157856 261772 157860
rect 261708 157800 261758 157856
rect 261758 157800 261772 157856
rect 261708 157796 261772 157800
rect 263916 157796 263980 157860
rect 266492 157796 266556 157860
rect 268332 157796 268396 157860
rect 265388 157660 265452 157724
rect 273668 157660 273732 157724
rect 278452 157660 278516 157724
rect 283604 157524 283668 157588
rect 290964 157584 291028 157588
rect 290964 157528 291014 157584
rect 291014 157528 291028 157584
rect 290964 157524 291028 157528
rect 244228 157388 244292 157452
rect 245516 157388 245580 157452
rect 253612 157448 253676 157452
rect 253612 157392 253662 157448
rect 253662 157392 253676 157448
rect 253612 157388 253676 157392
rect 256188 157448 256252 157452
rect 256188 157392 256238 157448
rect 256238 157392 256252 157448
rect 256188 157388 256252 157392
rect 363276 157388 363340 157452
rect 247724 156980 247788 157044
rect 216996 155484 217060 155548
rect 368612 153716 368676 153780
rect 368980 125564 369044 125628
rect 365116 99452 365180 99516
rect 367692 85580 367756 85644
rect 364932 45596 364996 45660
rect 364564 6564 364628 6628
rect 359044 6428 359108 6492
rect 358308 6292 358372 6356
rect 367324 6156 367388 6220
rect 359412 3980 359476 4044
rect 360148 3844 360212 3908
rect 215892 3572 215956 3636
rect 219204 3572 219268 3636
rect 358124 3708 358188 3772
rect 360700 3572 360764 3636
rect 365852 3572 365916 3636
rect 215156 3436 215220 3500
rect 216444 3436 216508 3500
rect 217548 3436 217612 3500
rect 218652 3436 218716 3500
rect 214420 3300 214484 3364
rect 356836 3300 356900 3364
rect 358492 3436 358556 3500
rect 358860 3436 358924 3500
rect 360332 3436 360396 3500
rect 361620 3436 361684 3500
rect 362908 3436 362972 3500
rect 364380 3436 364444 3500
rect 365668 3436 365732 3500
rect 367140 3436 367204 3500
rect 368428 3436 368492 3500
rect 369900 3436 369964 3500
rect 359228 3300 359292 3364
rect 369164 3300 369228 3364
rect 360516 3164 360580 3228
rect 363092 3028 363156 3092
<< metal4 >>
rect -9036 711868 -8416 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 -8416 711868
rect -9036 711548 -8416 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 -8416 711548
rect -9036 682954 -8416 711312
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 -8416 682954
rect -9036 682634 -8416 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 -8416 682634
rect -9036 646954 -8416 682398
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 -8416 646954
rect -9036 646634 -8416 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 -8416 646634
rect -9036 610954 -8416 646398
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 -8416 610954
rect -9036 610634 -8416 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 -8416 610634
rect -9036 574954 -8416 610398
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 -8416 574954
rect -9036 574634 -8416 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 -8416 574634
rect -9036 538954 -8416 574398
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 -8416 538954
rect -9036 538634 -8416 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 -8416 538634
rect -9036 502954 -8416 538398
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 -8416 502954
rect -9036 502634 -8416 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 -8416 502634
rect -9036 466954 -8416 502398
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 -8416 466954
rect -9036 466634 -8416 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 -8416 466634
rect -9036 430954 -8416 466398
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 -8416 430954
rect -9036 430634 -8416 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 -8416 430634
rect -9036 394954 -8416 430398
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 -8416 394954
rect -9036 394634 -8416 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 -8416 394634
rect -9036 358954 -8416 394398
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 -8416 358954
rect -9036 358634 -8416 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 -8416 358634
rect -9036 322954 -8416 358398
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 -8416 322954
rect -9036 322634 -8416 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 -8416 322634
rect -9036 286954 -8416 322398
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 -8416 286954
rect -9036 286634 -8416 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 -8416 286634
rect -9036 250954 -8416 286398
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 -8416 250954
rect -9036 250634 -8416 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 -8416 250634
rect -9036 214954 -8416 250398
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 -8416 214954
rect -9036 214634 -8416 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 -8416 214634
rect -9036 178954 -8416 214398
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 -8416 178954
rect -9036 178634 -8416 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 -8416 178634
rect -9036 142954 -8416 178398
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 -8416 142954
rect -9036 142634 -8416 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 -8416 142634
rect -9036 106954 -8416 142398
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 -8416 106954
rect -9036 106634 -8416 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 -8416 106634
rect -9036 70954 -8416 106398
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 -8416 70954
rect -9036 70634 -8416 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 -8416 70634
rect -9036 34954 -8416 70398
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 -8416 34954
rect -9036 34634 -8416 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 -8416 34634
rect -9036 -7376 -8416 34398
rect -8076 710908 -7456 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 -7456 710908
rect -8076 710588 -7456 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 -7456 710588
rect -8076 678454 -7456 710352
rect -8076 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 -7456 678454
rect -8076 678134 -7456 678218
rect -8076 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 -7456 678134
rect -8076 642454 -7456 677898
rect -8076 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 -7456 642454
rect -8076 642134 -7456 642218
rect -8076 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 -7456 642134
rect -8076 606454 -7456 641898
rect -8076 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 -7456 606454
rect -8076 606134 -7456 606218
rect -8076 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 -7456 606134
rect -8076 570454 -7456 605898
rect -8076 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 -7456 570454
rect -8076 570134 -7456 570218
rect -8076 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 -7456 570134
rect -8076 534454 -7456 569898
rect -8076 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 -7456 534454
rect -8076 534134 -7456 534218
rect -8076 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 -7456 534134
rect -8076 498454 -7456 533898
rect -8076 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 -7456 498454
rect -8076 498134 -7456 498218
rect -8076 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 -7456 498134
rect -8076 462454 -7456 497898
rect -8076 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 -7456 462454
rect -8076 462134 -7456 462218
rect -8076 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 -7456 462134
rect -8076 426454 -7456 461898
rect -8076 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 -7456 426454
rect -8076 426134 -7456 426218
rect -8076 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 -7456 426134
rect -8076 390454 -7456 425898
rect -8076 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 -7456 390454
rect -8076 390134 -7456 390218
rect -8076 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 -7456 390134
rect -8076 354454 -7456 389898
rect -8076 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 -7456 354454
rect -8076 354134 -7456 354218
rect -8076 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 -7456 354134
rect -8076 318454 -7456 353898
rect -8076 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 -7456 318454
rect -8076 318134 -7456 318218
rect -8076 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 -7456 318134
rect -8076 282454 -7456 317898
rect -8076 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 -7456 282454
rect -8076 282134 -7456 282218
rect -8076 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 -7456 282134
rect -8076 246454 -7456 281898
rect -8076 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 -7456 246454
rect -8076 246134 -7456 246218
rect -8076 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 -7456 246134
rect -8076 210454 -7456 245898
rect -8076 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 -7456 210454
rect -8076 210134 -7456 210218
rect -8076 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 -7456 210134
rect -8076 174454 -7456 209898
rect -8076 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 -7456 174454
rect -8076 174134 -7456 174218
rect -8076 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 -7456 174134
rect -8076 138454 -7456 173898
rect -8076 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 -7456 138454
rect -8076 138134 -7456 138218
rect -8076 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 -7456 138134
rect -8076 102454 -7456 137898
rect -8076 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 -7456 102454
rect -8076 102134 -7456 102218
rect -8076 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 -7456 102134
rect -8076 66454 -7456 101898
rect -8076 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 -7456 66454
rect -8076 66134 -7456 66218
rect -8076 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 -7456 66134
rect -8076 30454 -7456 65898
rect -8076 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 -7456 30454
rect -8076 30134 -7456 30218
rect -8076 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 -7456 30134
rect -8076 -6416 -7456 29898
rect -7116 709948 -6496 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 -6496 709948
rect -7116 709628 -6496 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 -6496 709628
rect -7116 673954 -6496 709392
rect -7116 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 -6496 673954
rect -7116 673634 -6496 673718
rect -7116 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 -6496 673634
rect -7116 637954 -6496 673398
rect -7116 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 -6496 637954
rect -7116 637634 -6496 637718
rect -7116 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 -6496 637634
rect -7116 601954 -6496 637398
rect -7116 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 -6496 601954
rect -7116 601634 -6496 601718
rect -7116 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 -6496 601634
rect -7116 565954 -6496 601398
rect -7116 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 -6496 565954
rect -7116 565634 -6496 565718
rect -7116 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 -6496 565634
rect -7116 529954 -6496 565398
rect -7116 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 -6496 529954
rect -7116 529634 -6496 529718
rect -7116 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 -6496 529634
rect -7116 493954 -6496 529398
rect -7116 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 -6496 493954
rect -7116 493634 -6496 493718
rect -7116 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 -6496 493634
rect -7116 457954 -6496 493398
rect -7116 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 -6496 457954
rect -7116 457634 -6496 457718
rect -7116 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 -6496 457634
rect -7116 421954 -6496 457398
rect -7116 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 -6496 421954
rect -7116 421634 -6496 421718
rect -7116 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 -6496 421634
rect -7116 385954 -6496 421398
rect -7116 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 -6496 385954
rect -7116 385634 -6496 385718
rect -7116 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 -6496 385634
rect -7116 349954 -6496 385398
rect -7116 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 -6496 349954
rect -7116 349634 -6496 349718
rect -7116 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 -6496 349634
rect -7116 313954 -6496 349398
rect -7116 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 -6496 313954
rect -7116 313634 -6496 313718
rect -7116 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 -6496 313634
rect -7116 277954 -6496 313398
rect -7116 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 -6496 277954
rect -7116 277634 -6496 277718
rect -7116 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 -6496 277634
rect -7116 241954 -6496 277398
rect -7116 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 -6496 241954
rect -7116 241634 -6496 241718
rect -7116 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 -6496 241634
rect -7116 205954 -6496 241398
rect -7116 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 -6496 205954
rect -7116 205634 -6496 205718
rect -7116 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 -6496 205634
rect -7116 169954 -6496 205398
rect -7116 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 -6496 169954
rect -7116 169634 -6496 169718
rect -7116 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 -6496 169634
rect -7116 133954 -6496 169398
rect -7116 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 -6496 133954
rect -7116 133634 -6496 133718
rect -7116 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 -6496 133634
rect -7116 97954 -6496 133398
rect -7116 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 -6496 97954
rect -7116 97634 -6496 97718
rect -7116 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 -6496 97634
rect -7116 61954 -6496 97398
rect -7116 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 -6496 61954
rect -7116 61634 -6496 61718
rect -7116 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 -6496 61634
rect -7116 25954 -6496 61398
rect -7116 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 -6496 25954
rect -7116 25634 -6496 25718
rect -7116 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 -6496 25634
rect -7116 -5456 -6496 25398
rect -6156 708988 -5536 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 -5536 708988
rect -6156 708668 -5536 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 -5536 708668
rect -6156 669454 -5536 708432
rect -6156 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 -5536 669454
rect -6156 669134 -5536 669218
rect -6156 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 -5536 669134
rect -6156 633454 -5536 668898
rect -6156 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 -5536 633454
rect -6156 633134 -5536 633218
rect -6156 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 -5536 633134
rect -6156 597454 -5536 632898
rect -6156 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 -5536 597454
rect -6156 597134 -5536 597218
rect -6156 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 -5536 597134
rect -6156 561454 -5536 596898
rect -6156 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 -5536 561454
rect -6156 561134 -5536 561218
rect -6156 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 -5536 561134
rect -6156 525454 -5536 560898
rect -6156 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 -5536 525454
rect -6156 525134 -5536 525218
rect -6156 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 -5536 525134
rect -6156 489454 -5536 524898
rect -6156 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 -5536 489454
rect -6156 489134 -5536 489218
rect -6156 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 -5536 489134
rect -6156 453454 -5536 488898
rect -6156 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 -5536 453454
rect -6156 453134 -5536 453218
rect -6156 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 -5536 453134
rect -6156 417454 -5536 452898
rect -6156 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 -5536 417454
rect -6156 417134 -5536 417218
rect -6156 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 -5536 417134
rect -6156 381454 -5536 416898
rect -6156 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 -5536 381454
rect -6156 381134 -5536 381218
rect -6156 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 -5536 381134
rect -6156 345454 -5536 380898
rect -6156 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 -5536 345454
rect -6156 345134 -5536 345218
rect -6156 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 -5536 345134
rect -6156 309454 -5536 344898
rect -6156 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 -5536 309454
rect -6156 309134 -5536 309218
rect -6156 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 -5536 309134
rect -6156 273454 -5536 308898
rect -6156 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 -5536 273454
rect -6156 273134 -5536 273218
rect -6156 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 -5536 273134
rect -6156 237454 -5536 272898
rect -6156 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 -5536 237454
rect -6156 237134 -5536 237218
rect -6156 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 -5536 237134
rect -6156 201454 -5536 236898
rect -6156 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 -5536 201454
rect -6156 201134 -5536 201218
rect -6156 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 -5536 201134
rect -6156 165454 -5536 200898
rect -6156 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 -5536 165454
rect -6156 165134 -5536 165218
rect -6156 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 -5536 165134
rect -6156 129454 -5536 164898
rect -6156 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 -5536 129454
rect -6156 129134 -5536 129218
rect -6156 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 -5536 129134
rect -6156 93454 -5536 128898
rect -6156 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 -5536 93454
rect -6156 93134 -5536 93218
rect -6156 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 -5536 93134
rect -6156 57454 -5536 92898
rect -6156 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 -5536 57454
rect -6156 57134 -5536 57218
rect -6156 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 -5536 57134
rect -6156 21454 -5536 56898
rect -6156 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 -5536 21454
rect -6156 21134 -5536 21218
rect -6156 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 -5536 21134
rect -6156 -4496 -5536 20898
rect -5196 708028 -4576 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 -4576 708028
rect -5196 707708 -4576 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 -4576 707708
rect -5196 700954 -4576 707472
rect -5196 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 -4576 700954
rect -5196 700634 -4576 700718
rect -5196 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 -4576 700634
rect -5196 664954 -4576 700398
rect -5196 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 -4576 664954
rect -5196 664634 -4576 664718
rect -5196 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 -4576 664634
rect -5196 628954 -4576 664398
rect -5196 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 -4576 628954
rect -5196 628634 -4576 628718
rect -5196 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 -4576 628634
rect -5196 592954 -4576 628398
rect -5196 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 -4576 592954
rect -5196 592634 -4576 592718
rect -5196 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 -4576 592634
rect -5196 556954 -4576 592398
rect -5196 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 -4576 556954
rect -5196 556634 -4576 556718
rect -5196 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 -4576 556634
rect -5196 520954 -4576 556398
rect -5196 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 -4576 520954
rect -5196 520634 -4576 520718
rect -5196 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 -4576 520634
rect -5196 484954 -4576 520398
rect -5196 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 -4576 484954
rect -5196 484634 -4576 484718
rect -5196 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 -4576 484634
rect -5196 448954 -4576 484398
rect -5196 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 -4576 448954
rect -5196 448634 -4576 448718
rect -5196 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 -4576 448634
rect -5196 412954 -4576 448398
rect -5196 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 -4576 412954
rect -5196 412634 -4576 412718
rect -5196 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 -4576 412634
rect -5196 376954 -4576 412398
rect -5196 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 -4576 376954
rect -5196 376634 -4576 376718
rect -5196 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 -4576 376634
rect -5196 340954 -4576 376398
rect -5196 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 -4576 340954
rect -5196 340634 -4576 340718
rect -5196 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 -4576 340634
rect -5196 304954 -4576 340398
rect -5196 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 -4576 304954
rect -5196 304634 -4576 304718
rect -5196 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 -4576 304634
rect -5196 268954 -4576 304398
rect -5196 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 -4576 268954
rect -5196 268634 -4576 268718
rect -5196 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 -4576 268634
rect -5196 232954 -4576 268398
rect -5196 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 -4576 232954
rect -5196 232634 -4576 232718
rect -5196 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 -4576 232634
rect -5196 196954 -4576 232398
rect -5196 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 -4576 196954
rect -5196 196634 -4576 196718
rect -5196 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 -4576 196634
rect -5196 160954 -4576 196398
rect -5196 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 -4576 160954
rect -5196 160634 -4576 160718
rect -5196 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 -4576 160634
rect -5196 124954 -4576 160398
rect -5196 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 -4576 124954
rect -5196 124634 -4576 124718
rect -5196 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 -4576 124634
rect -5196 88954 -4576 124398
rect -5196 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 -4576 88954
rect -5196 88634 -4576 88718
rect -5196 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 -4576 88634
rect -5196 52954 -4576 88398
rect -5196 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 -4576 52954
rect -5196 52634 -4576 52718
rect -5196 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 -4576 52634
rect -5196 16954 -4576 52398
rect -5196 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 -4576 16954
rect -5196 16634 -4576 16718
rect -5196 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 -4576 16634
rect -5196 -3536 -4576 16398
rect -4236 707068 -3616 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 -3616 707068
rect -4236 706748 -3616 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 -3616 706748
rect -4236 696454 -3616 706512
rect -4236 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 -3616 696454
rect -4236 696134 -3616 696218
rect -4236 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 -3616 696134
rect -4236 660454 -3616 695898
rect -4236 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 -3616 660454
rect -4236 660134 -3616 660218
rect -4236 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 -3616 660134
rect -4236 624454 -3616 659898
rect -4236 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 -3616 624454
rect -4236 624134 -3616 624218
rect -4236 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 -3616 624134
rect -4236 588454 -3616 623898
rect -4236 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 -3616 588454
rect -4236 588134 -3616 588218
rect -4236 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 -3616 588134
rect -4236 552454 -3616 587898
rect -4236 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 -3616 552454
rect -4236 552134 -3616 552218
rect -4236 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 -3616 552134
rect -4236 516454 -3616 551898
rect -4236 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 -3616 516454
rect -4236 516134 -3616 516218
rect -4236 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 -3616 516134
rect -4236 480454 -3616 515898
rect -4236 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 -3616 480454
rect -4236 480134 -3616 480218
rect -4236 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 -3616 480134
rect -4236 444454 -3616 479898
rect -4236 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 -3616 444454
rect -4236 444134 -3616 444218
rect -4236 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 -3616 444134
rect -4236 408454 -3616 443898
rect -4236 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 -3616 408454
rect -4236 408134 -3616 408218
rect -4236 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 -3616 408134
rect -4236 372454 -3616 407898
rect -4236 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 -3616 372454
rect -4236 372134 -3616 372218
rect -4236 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 -3616 372134
rect -4236 336454 -3616 371898
rect -4236 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 -3616 336454
rect -4236 336134 -3616 336218
rect -4236 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 -3616 336134
rect -4236 300454 -3616 335898
rect -4236 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 -3616 300454
rect -4236 300134 -3616 300218
rect -4236 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 -3616 300134
rect -4236 264454 -3616 299898
rect -4236 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 -3616 264454
rect -4236 264134 -3616 264218
rect -4236 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 -3616 264134
rect -4236 228454 -3616 263898
rect -4236 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 -3616 228454
rect -4236 228134 -3616 228218
rect -4236 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 -3616 228134
rect -4236 192454 -3616 227898
rect -4236 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 -3616 192454
rect -4236 192134 -3616 192218
rect -4236 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 -3616 192134
rect -4236 156454 -3616 191898
rect -4236 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 -3616 156454
rect -4236 156134 -3616 156218
rect -4236 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 -3616 156134
rect -4236 120454 -3616 155898
rect -4236 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 -3616 120454
rect -4236 120134 -3616 120218
rect -4236 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 -3616 120134
rect -4236 84454 -3616 119898
rect -4236 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 -3616 84454
rect -4236 84134 -3616 84218
rect -4236 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 -3616 84134
rect -4236 48454 -3616 83898
rect -4236 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 -3616 48454
rect -4236 48134 -3616 48218
rect -4236 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 -3616 48134
rect -4236 12454 -3616 47898
rect -4236 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 -3616 12454
rect -4236 12134 -3616 12218
rect -4236 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 -3616 12134
rect -4236 -2576 -3616 11898
rect -3276 706108 -2656 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 -2656 706108
rect -3276 705788 -2656 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 -2656 705788
rect -3276 691954 -2656 705552
rect -3276 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 -2656 691954
rect -3276 691634 -2656 691718
rect -3276 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 -2656 691634
rect -3276 655954 -2656 691398
rect -3276 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 -2656 655954
rect -3276 655634 -2656 655718
rect -3276 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 -2656 655634
rect -3276 619954 -2656 655398
rect -3276 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 -2656 619954
rect -3276 619634 -2656 619718
rect -3276 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 -2656 619634
rect -3276 583954 -2656 619398
rect -3276 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 -2656 583954
rect -3276 583634 -2656 583718
rect -3276 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 -2656 583634
rect -3276 547954 -2656 583398
rect -3276 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 -2656 547954
rect -3276 547634 -2656 547718
rect -3276 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 -2656 547634
rect -3276 511954 -2656 547398
rect -3276 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 -2656 511954
rect -3276 511634 -2656 511718
rect -3276 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 -2656 511634
rect -3276 475954 -2656 511398
rect -3276 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 -2656 475954
rect -3276 475634 -2656 475718
rect -3276 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 -2656 475634
rect -3276 439954 -2656 475398
rect -3276 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 -2656 439954
rect -3276 439634 -2656 439718
rect -3276 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 -2656 439634
rect -3276 403954 -2656 439398
rect -3276 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 -2656 403954
rect -3276 403634 -2656 403718
rect -3276 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 -2656 403634
rect -3276 367954 -2656 403398
rect -3276 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 -2656 367954
rect -3276 367634 -2656 367718
rect -3276 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 -2656 367634
rect -3276 331954 -2656 367398
rect -3276 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 -2656 331954
rect -3276 331634 -2656 331718
rect -3276 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 -2656 331634
rect -3276 295954 -2656 331398
rect -3276 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 -2656 295954
rect -3276 295634 -2656 295718
rect -3276 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 -2656 295634
rect -3276 259954 -2656 295398
rect -3276 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 -2656 259954
rect -3276 259634 -2656 259718
rect -3276 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 -2656 259634
rect -3276 223954 -2656 259398
rect -3276 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 -2656 223954
rect -3276 223634 -2656 223718
rect -3276 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 -2656 223634
rect -3276 187954 -2656 223398
rect -3276 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 -2656 187954
rect -3276 187634 -2656 187718
rect -3276 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 -2656 187634
rect -3276 151954 -2656 187398
rect -3276 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 -2656 151954
rect -3276 151634 -2656 151718
rect -3276 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 -2656 151634
rect -3276 115954 -2656 151398
rect -3276 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 -2656 115954
rect -3276 115634 -2656 115718
rect -3276 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 -2656 115634
rect -3276 79954 -2656 115398
rect -3276 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 -2656 79954
rect -3276 79634 -2656 79718
rect -3276 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 -2656 79634
rect -3276 43954 -2656 79398
rect -3276 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 -2656 43954
rect -3276 43634 -2656 43718
rect -3276 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 -2656 43634
rect -3276 7954 -2656 43398
rect -3276 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 -2656 7954
rect -3276 7634 -2656 7718
rect -3276 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 -2656 7634
rect -3276 -1616 -2656 7398
rect -2316 705148 -1696 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 -1696 705148
rect -2316 704828 -1696 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 -1696 704828
rect -2316 687454 -1696 704592
rect -2316 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 -1696 687454
rect -2316 687134 -1696 687218
rect -2316 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 -1696 687134
rect -2316 651454 -1696 686898
rect -2316 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 -1696 651454
rect -2316 651134 -1696 651218
rect -2316 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 -1696 651134
rect -2316 615454 -1696 650898
rect -2316 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 -1696 615454
rect -2316 615134 -1696 615218
rect -2316 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 -1696 615134
rect -2316 579454 -1696 614898
rect -2316 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 -1696 579454
rect -2316 579134 -1696 579218
rect -2316 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 -1696 579134
rect -2316 543454 -1696 578898
rect -2316 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 -1696 543454
rect -2316 543134 -1696 543218
rect -2316 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 -1696 543134
rect -2316 507454 -1696 542898
rect -2316 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 -1696 507454
rect -2316 507134 -1696 507218
rect -2316 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 -1696 507134
rect -2316 471454 -1696 506898
rect -2316 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 -1696 471454
rect -2316 471134 -1696 471218
rect -2316 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 -1696 471134
rect -2316 435454 -1696 470898
rect -2316 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 -1696 435454
rect -2316 435134 -1696 435218
rect -2316 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 -1696 435134
rect -2316 399454 -1696 434898
rect -2316 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 -1696 399454
rect -2316 399134 -1696 399218
rect -2316 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 -1696 399134
rect -2316 363454 -1696 398898
rect -2316 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 -1696 363454
rect -2316 363134 -1696 363218
rect -2316 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 -1696 363134
rect -2316 327454 -1696 362898
rect -2316 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 -1696 327454
rect -2316 327134 -1696 327218
rect -2316 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 -1696 327134
rect -2316 291454 -1696 326898
rect -2316 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 -1696 291454
rect -2316 291134 -1696 291218
rect -2316 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 -1696 291134
rect -2316 255454 -1696 290898
rect -2316 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 -1696 255454
rect -2316 255134 -1696 255218
rect -2316 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 -1696 255134
rect -2316 219454 -1696 254898
rect -2316 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 -1696 219454
rect -2316 219134 -1696 219218
rect -2316 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 -1696 219134
rect -2316 183454 -1696 218898
rect -2316 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 -1696 183454
rect -2316 183134 -1696 183218
rect -2316 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 -1696 183134
rect -2316 147454 -1696 182898
rect -2316 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 -1696 147454
rect -2316 147134 -1696 147218
rect -2316 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 -1696 147134
rect -2316 111454 -1696 146898
rect -2316 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 -1696 111454
rect -2316 111134 -1696 111218
rect -2316 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 -1696 111134
rect -2316 75454 -1696 110898
rect -2316 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 -1696 75454
rect -2316 75134 -1696 75218
rect -2316 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 -1696 75134
rect -2316 39454 -1696 74898
rect -2316 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 -1696 39454
rect -2316 39134 -1696 39218
rect -2316 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 -1696 39134
rect -2316 3454 -1696 38898
rect -2316 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 -1696 3454
rect -2316 3134 -1696 3218
rect -2316 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 -1696 3134
rect -2316 -656 -1696 2898
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 -1696 -656
rect -2316 -976 -1696 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 -1696 -976
rect -2316 -1244 -1696 -1212
rect 1794 705148 2414 711900
rect 1794 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 2414 705148
rect 1794 704828 2414 704912
rect 1794 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 2414 704828
rect 1794 687454 2414 704592
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -656 2414 2898
rect 1794 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 2414 -656
rect 1794 -976 2414 -892
rect 1794 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 2414 -976
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 -2656 -1616
rect -3276 -1936 -2656 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 -2656 -1936
rect -3276 -2204 -2656 -2172
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 -3616 -2576
rect -4236 -2896 -3616 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 -3616 -2896
rect -4236 -3164 -3616 -3132
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 -4576 -3536
rect -5196 -3856 -4576 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 -4576 -3856
rect -5196 -4124 -4576 -4092
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 -5536 -4496
rect -6156 -4816 -5536 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 -5536 -4816
rect -6156 -5084 -5536 -5052
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 -6496 -5456
rect -7116 -5776 -6496 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 -6496 -5776
rect -7116 -6044 -6496 -6012
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 -7456 -6416
rect -8076 -6736 -7456 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 -7456 -6736
rect -8076 -7004 -7456 -6972
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 -8416 -7376
rect -9036 -7696 -8416 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 -8416 -7696
rect -9036 -7964 -8416 -7932
rect 1794 -7964 2414 -1212
rect 6294 706108 6914 711900
rect 6294 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 6914 706108
rect 6294 705788 6914 705872
rect 6294 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 6914 705788
rect 6294 691954 6914 705552
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1616 6914 7398
rect 6294 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 6914 -1616
rect 6294 -1936 6914 -1852
rect 6294 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 6914 -1936
rect 6294 -7964 6914 -2172
rect 10794 707068 11414 711900
rect 10794 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 11414 707068
rect 10794 706748 11414 706832
rect 10794 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 11414 706748
rect 10794 696454 11414 706512
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2576 11414 11898
rect 10794 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 11414 -2576
rect 10794 -2896 11414 -2812
rect 10794 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 11414 -2896
rect 10794 -7964 11414 -3132
rect 15294 708028 15914 711900
rect 15294 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 15914 708028
rect 15294 707708 15914 707792
rect 15294 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 15914 707708
rect 15294 700954 15914 707472
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3536 15914 16398
rect 15294 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 15914 -3536
rect 15294 -3856 15914 -3772
rect 15294 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 15914 -3856
rect 15294 -7964 15914 -4092
rect 19794 708988 20414 711900
rect 19794 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 20414 708988
rect 19794 708668 20414 708752
rect 19794 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 20414 708668
rect 19794 669454 20414 708432
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4496 20414 20898
rect 19794 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 20414 -4496
rect 19794 -4816 20414 -4732
rect 19794 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 20414 -4816
rect 19794 -7964 20414 -5052
rect 24294 709948 24914 711900
rect 24294 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 24914 709948
rect 24294 709628 24914 709712
rect 24294 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 24914 709628
rect 24294 673954 24914 709392
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5456 24914 25398
rect 24294 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 24914 -5456
rect 24294 -5776 24914 -5692
rect 24294 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 24914 -5776
rect 24294 -7964 24914 -6012
rect 28794 710908 29414 711900
rect 28794 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 29414 710908
rect 28794 710588 29414 710672
rect 28794 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 29414 710588
rect 28794 678454 29414 710352
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6416 29414 29898
rect 28794 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 29414 -6416
rect 28794 -6736 29414 -6652
rect 28794 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 29414 -6736
rect 28794 -7964 29414 -6972
rect 33294 711868 33914 711900
rect 33294 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 33914 711868
rect 33294 711548 33914 711632
rect 33294 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 33914 711548
rect 33294 682954 33914 711312
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7376 33914 34398
rect 33294 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 33914 -7376
rect 33294 -7696 33914 -7612
rect 33294 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 33914 -7696
rect 33294 -7964 33914 -7932
rect 37794 705148 38414 711900
rect 37794 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 38414 705148
rect 37794 704828 38414 704912
rect 37794 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 38414 704828
rect 37794 687454 38414 704592
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -656 38414 2898
rect 37794 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 38414 -656
rect 37794 -976 38414 -892
rect 37794 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 38414 -976
rect 37794 -7964 38414 -1212
rect 42294 706108 42914 711900
rect 42294 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 42914 706108
rect 42294 705788 42914 705872
rect 42294 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 42914 705788
rect 42294 691954 42914 705552
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1616 42914 7398
rect 42294 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 42914 -1616
rect 42294 -1936 42914 -1852
rect 42294 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 42914 -1936
rect 42294 -7964 42914 -2172
rect 46794 707068 47414 711900
rect 46794 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 47414 707068
rect 46794 706748 47414 706832
rect 46794 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 47414 706748
rect 46794 696454 47414 706512
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2576 47414 11898
rect 46794 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 47414 -2576
rect 46794 -2896 47414 -2812
rect 46794 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 47414 -2896
rect 46794 -7964 47414 -3132
rect 51294 708028 51914 711900
rect 51294 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 51914 708028
rect 51294 707708 51914 707792
rect 51294 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 51914 707708
rect 51294 700954 51914 707472
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3536 51914 16398
rect 51294 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 51914 -3536
rect 51294 -3856 51914 -3772
rect 51294 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 51914 -3856
rect 51294 -7964 51914 -4092
rect 55794 708988 56414 711900
rect 55794 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 56414 708988
rect 55794 708668 56414 708752
rect 55794 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 56414 708668
rect 55794 669454 56414 708432
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4496 56414 20898
rect 55794 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 56414 -4496
rect 55794 -4816 56414 -4732
rect 55794 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 56414 -4816
rect 55794 -7964 56414 -5052
rect 60294 709948 60914 711900
rect 60294 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 60914 709948
rect 60294 709628 60914 709712
rect 60294 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 60914 709628
rect 60294 673954 60914 709392
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5456 60914 25398
rect 60294 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 60914 -5456
rect 60294 -5776 60914 -5692
rect 60294 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 60914 -5776
rect 60294 -7964 60914 -6012
rect 64794 710908 65414 711900
rect 64794 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 65414 710908
rect 64794 710588 65414 710672
rect 64794 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 65414 710588
rect 64794 678454 65414 710352
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6416 65414 29898
rect 64794 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 65414 -6416
rect 64794 -6736 65414 -6652
rect 64794 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 65414 -6736
rect 64794 -7964 65414 -6972
rect 69294 711868 69914 711900
rect 69294 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 69914 711868
rect 69294 711548 69914 711632
rect 69294 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 69914 711548
rect 69294 682954 69914 711312
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7376 69914 34398
rect 69294 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 69914 -7376
rect 69294 -7696 69914 -7612
rect 69294 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 69914 -7696
rect 69294 -7964 69914 -7932
rect 73794 705148 74414 711900
rect 73794 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 74414 705148
rect 73794 704828 74414 704912
rect 73794 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 74414 704828
rect 73794 687454 74414 704592
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -656 74414 2898
rect 73794 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 74414 -656
rect 73794 -976 74414 -892
rect 73794 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 74414 -976
rect 73794 -7964 74414 -1212
rect 78294 706108 78914 711900
rect 78294 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 78914 706108
rect 78294 705788 78914 705872
rect 78294 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 78914 705788
rect 78294 691954 78914 705552
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1616 78914 7398
rect 78294 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 78914 -1616
rect 78294 -1936 78914 -1852
rect 78294 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 78914 -1936
rect 78294 -7964 78914 -2172
rect 82794 707068 83414 711900
rect 82794 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 83414 707068
rect 82794 706748 83414 706832
rect 82794 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 83414 706748
rect 82794 696454 83414 706512
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2576 83414 11898
rect 82794 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 83414 -2576
rect 82794 -2896 83414 -2812
rect 82794 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 83414 -2896
rect 82794 -7964 83414 -3132
rect 87294 708028 87914 711900
rect 87294 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 87914 708028
rect 87294 707708 87914 707792
rect 87294 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 87914 707708
rect 87294 700954 87914 707472
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3536 87914 16398
rect 87294 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 87914 -3536
rect 87294 -3856 87914 -3772
rect 87294 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 87914 -3856
rect 87294 -7964 87914 -4092
rect 91794 708988 92414 711900
rect 91794 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 92414 708988
rect 91794 708668 92414 708752
rect 91794 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 92414 708668
rect 91794 669454 92414 708432
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4496 92414 20898
rect 91794 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 92414 -4496
rect 91794 -4816 92414 -4732
rect 91794 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 92414 -4816
rect 91794 -7964 92414 -5052
rect 96294 709948 96914 711900
rect 96294 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 96914 709948
rect 96294 709628 96914 709712
rect 96294 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 96914 709628
rect 96294 673954 96914 709392
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 100794 710908 101414 711900
rect 100794 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 101414 710908
rect 100794 710588 101414 710672
rect 100794 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 101414 710588
rect 100794 678454 101414 710352
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 374164 101414 389898
rect 105294 711868 105914 711900
rect 105294 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 105914 711868
rect 105294 711548 105914 711632
rect 105294 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 105914 711548
rect 105294 682954 105914 711312
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 374164 105914 394398
rect 109794 705148 110414 711900
rect 109794 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 110414 705148
rect 109794 704828 110414 704912
rect 109794 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 110414 704828
rect 109794 687454 110414 704592
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 374164 110414 398898
rect 114294 706108 114914 711900
rect 114294 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 114914 706108
rect 114294 705788 114914 705872
rect 114294 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 114914 705788
rect 114294 691954 114914 705552
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 374164 114914 403398
rect 118794 707068 119414 711900
rect 118794 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 119414 707068
rect 118794 706748 119414 706832
rect 118794 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 119414 706748
rect 118794 696454 119414 706512
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 374164 119414 407898
rect 123294 708028 123914 711900
rect 123294 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 123914 708028
rect 123294 707708 123914 707792
rect 123294 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 123914 707708
rect 123294 700954 123914 707472
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 374164 123914 376398
rect 127794 708988 128414 711900
rect 127794 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 128414 708988
rect 127794 708668 128414 708752
rect 127794 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 128414 708668
rect 127794 669454 128414 708432
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 374164 128414 380898
rect 132294 709948 132914 711900
rect 132294 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 132914 709948
rect 132294 709628 132914 709712
rect 132294 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 132914 709628
rect 132294 673954 132914 709392
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 374164 132914 385398
rect 136794 710908 137414 711900
rect 136794 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 137414 710908
rect 136794 710588 137414 710672
rect 136794 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 137414 710588
rect 136794 678454 137414 710352
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 374164 137414 389898
rect 141294 711868 141914 711900
rect 141294 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 141914 711868
rect 141294 711548 141914 711632
rect 141294 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 141914 711548
rect 141294 682954 141914 711312
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 374164 141914 394398
rect 145794 705148 146414 711900
rect 145794 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 146414 705148
rect 145794 704828 146414 704912
rect 145794 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 146414 704828
rect 145794 687454 146414 704592
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 374164 146414 398898
rect 150294 706108 150914 711900
rect 150294 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 150914 706108
rect 150294 705788 150914 705872
rect 150294 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 150914 705788
rect 150294 691954 150914 705552
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 374164 150914 403398
rect 154794 707068 155414 711900
rect 154794 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 155414 707068
rect 154794 706748 155414 706832
rect 154794 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 155414 706748
rect 154794 696454 155414 706512
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 374164 155414 407898
rect 159294 708028 159914 711900
rect 159294 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 159914 708028
rect 159294 707708 159914 707792
rect 159294 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 159914 707708
rect 159294 700954 159914 707472
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 374164 159914 376398
rect 163794 708988 164414 711900
rect 163794 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 164414 708988
rect 163794 708668 164414 708752
rect 163794 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 164414 708668
rect 163794 669454 164414 708432
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 374164 164414 380898
rect 168294 709948 168914 711900
rect 168294 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 168914 709948
rect 168294 709628 168914 709712
rect 168294 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 168914 709628
rect 168294 673954 168914 709392
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 374164 168914 385398
rect 172794 710908 173414 711900
rect 172794 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 173414 710908
rect 172794 710588 173414 710672
rect 172794 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 173414 710588
rect 172794 678454 173414 710352
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 119568 367954 119888 367986
rect 119568 367718 119610 367954
rect 119846 367718 119888 367954
rect 119568 367634 119888 367718
rect 119568 367398 119610 367634
rect 119846 367398 119888 367634
rect 119568 367366 119888 367398
rect 150288 367954 150608 367986
rect 150288 367718 150330 367954
rect 150566 367718 150608 367954
rect 150288 367634 150608 367718
rect 150288 367398 150330 367634
rect 150566 367398 150608 367634
rect 150288 367366 150608 367398
rect 104208 363454 104528 363486
rect 104208 363218 104250 363454
rect 104486 363218 104528 363454
rect 104208 363134 104528 363218
rect 104208 362898 104250 363134
rect 104486 362898 104528 363134
rect 104208 362866 104528 362898
rect 134928 363454 135248 363486
rect 134928 363218 134970 363454
rect 135206 363218 135248 363454
rect 134928 363134 135248 363218
rect 134928 362898 134970 363134
rect 135206 362898 135248 363134
rect 134928 362866 135248 362898
rect 165648 363454 165968 363486
rect 165648 363218 165690 363454
rect 165926 363218 165968 363454
rect 165648 363134 165968 363218
rect 165648 362898 165690 363134
rect 165926 362898 165968 363134
rect 165648 362866 165968 362898
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 119568 331954 119888 331986
rect 119568 331718 119610 331954
rect 119846 331718 119888 331954
rect 119568 331634 119888 331718
rect 119568 331398 119610 331634
rect 119846 331398 119888 331634
rect 119568 331366 119888 331398
rect 150288 331954 150608 331986
rect 150288 331718 150330 331954
rect 150566 331718 150608 331954
rect 150288 331634 150608 331718
rect 150288 331398 150330 331634
rect 150566 331398 150608 331634
rect 150288 331366 150608 331398
rect 104208 327454 104528 327486
rect 104208 327218 104250 327454
rect 104486 327218 104528 327454
rect 104208 327134 104528 327218
rect 104208 326898 104250 327134
rect 104486 326898 104528 327134
rect 104208 326866 104528 326898
rect 134928 327454 135248 327486
rect 134928 327218 134970 327454
rect 135206 327218 135248 327454
rect 134928 327134 135248 327218
rect 134928 326898 134970 327134
rect 135206 326898 135248 327134
rect 134928 326866 135248 326898
rect 165648 327454 165968 327486
rect 165648 327218 165690 327454
rect 165926 327218 165968 327454
rect 165648 327134 165968 327218
rect 165648 326898 165690 327134
rect 165926 326898 165968 327134
rect 165648 326866 165968 326898
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 169339 308548 169405 308549
rect 169339 308484 169340 308548
rect 169404 308484 169405 308548
rect 169339 308483 169405 308484
rect 169155 301204 169221 301205
rect 169155 301140 169156 301204
rect 169220 301140 169221 301204
rect 169155 301139 169221 301140
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5456 96914 25398
rect 96294 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 96914 -5456
rect 96294 -5776 96914 -5692
rect 96294 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 96914 -5776
rect 96294 -7964 96914 -6012
rect 100794 282454 101414 298000
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6416 101414 29898
rect 100794 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 101414 -6416
rect 100794 -6736 101414 -6652
rect 100794 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 101414 -6736
rect 100794 -7964 101414 -6972
rect 105294 286954 105914 298000
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7376 105914 34398
rect 105294 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 105914 -7376
rect 105294 -7696 105914 -7612
rect 105294 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 105914 -7696
rect 105294 -7964 105914 -7932
rect 109794 291454 110414 298000
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -656 110414 2898
rect 109794 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 110414 -656
rect 109794 -976 110414 -892
rect 109794 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 110414 -976
rect 109794 -7964 110414 -1212
rect 114294 295954 114914 298000
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1616 114914 7398
rect 114294 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 114914 -1616
rect 114294 -1936 114914 -1852
rect 114294 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 114914 -1936
rect 114294 -7964 114914 -2172
rect 118794 264454 119414 298000
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2576 119414 11898
rect 118794 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 119414 -2576
rect 118794 -2896 119414 -2812
rect 118794 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 119414 -2896
rect 118794 -7964 119414 -3132
rect 123294 268954 123914 298000
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3536 123914 16398
rect 123294 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 123914 -3536
rect 123294 -3856 123914 -3772
rect 123294 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 123914 -3856
rect 123294 -7964 123914 -4092
rect 127794 273454 128414 298000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4496 128414 20898
rect 127794 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 128414 -4496
rect 127794 -4816 128414 -4732
rect 127794 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 128414 -4816
rect 127794 -7964 128414 -5052
rect 132294 277954 132914 298000
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5456 132914 25398
rect 132294 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 132914 -5456
rect 132294 -5776 132914 -5692
rect 132294 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 132914 -5776
rect 132294 -7964 132914 -6012
rect 136794 282454 137414 298000
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6416 137414 29898
rect 136794 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 137414 -6416
rect 136794 -6736 137414 -6652
rect 136794 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 137414 -6736
rect 136794 -7964 137414 -6972
rect 141294 286954 141914 298000
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7376 141914 34398
rect 141294 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 141914 -7376
rect 141294 -7696 141914 -7612
rect 141294 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 141914 -7696
rect 141294 -7964 141914 -7932
rect 145794 291454 146414 298000
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -656 146414 2898
rect 145794 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 146414 -656
rect 145794 -976 146414 -892
rect 145794 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 146414 -976
rect 145794 -7964 146414 -1212
rect 150294 295954 150914 298000
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1616 150914 7398
rect 150294 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 150914 -1616
rect 150294 -1936 150914 -1852
rect 150294 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 150914 -1936
rect 150294 -7964 150914 -2172
rect 154794 264454 155414 298000
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2576 155414 11898
rect 154794 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 155414 -2576
rect 154794 -2896 155414 -2812
rect 154794 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 155414 -2896
rect 154794 -7964 155414 -3132
rect 159294 268954 159914 298000
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3536 159914 16398
rect 159294 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 159914 -3536
rect 159294 -3856 159914 -3772
rect 159294 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 159914 -3856
rect 159294 -7964 159914 -4092
rect 163794 273454 164414 298000
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4496 164414 20898
rect 163794 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 164414 -4496
rect 163794 -4816 164414 -4732
rect 163794 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 164414 -4816
rect 163794 -7964 164414 -5052
rect 168294 277954 168914 298000
rect 169158 297941 169218 301139
rect 169342 299165 169402 308483
rect 169707 301612 169773 301613
rect 169707 301548 169708 301612
rect 169772 301548 169773 301612
rect 169707 301547 169773 301548
rect 169339 299164 169405 299165
rect 169339 299100 169340 299164
rect 169404 299100 169405 299164
rect 169339 299099 169405 299100
rect 169155 297940 169221 297941
rect 169155 297876 169156 297940
rect 169220 297876 169221 297940
rect 169155 297875 169221 297876
rect 169710 297805 169770 301547
rect 169707 297804 169773 297805
rect 169707 297740 169708 297804
rect 169772 297740 169773 297804
rect 169707 297739 169773 297740
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5456 168914 25398
rect 168294 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 168914 -5456
rect 168294 -5776 168914 -5692
rect 168294 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 168914 -5776
rect 168294 -7964 168914 -6012
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6416 173414 29898
rect 172794 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 173414 -6416
rect 172794 -6736 173414 -6652
rect 172794 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 173414 -6736
rect 172794 -7964 173414 -6972
rect 177294 711868 177914 711900
rect 177294 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 177914 711868
rect 177294 711548 177914 711632
rect 177294 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 177914 711548
rect 177294 682954 177914 711312
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7376 177914 34398
rect 177294 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 177914 -7376
rect 177294 -7696 177914 -7612
rect 177294 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 177914 -7696
rect 177294 -7964 177914 -7932
rect 181794 705148 182414 711900
rect 181794 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 182414 705148
rect 181794 704828 182414 704912
rect 181794 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 182414 704828
rect 181794 687454 182414 704592
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -656 182414 2898
rect 181794 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 182414 -656
rect 181794 -976 182414 -892
rect 181794 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 182414 -976
rect 181794 -7964 182414 -1212
rect 186294 706108 186914 711900
rect 186294 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 186914 706108
rect 186294 705788 186914 705872
rect 186294 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 186914 705788
rect 186294 691954 186914 705552
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1616 186914 7398
rect 186294 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 186914 -1616
rect 186294 -1936 186914 -1852
rect 186294 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 186914 -1936
rect 186294 -7964 186914 -2172
rect 190794 707068 191414 711900
rect 190794 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 191414 707068
rect 190794 706748 191414 706832
rect 190794 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 191414 706748
rect 190794 696454 191414 706512
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2576 191414 11898
rect 190794 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 191414 -2576
rect 190794 -2896 191414 -2812
rect 190794 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 191414 -2896
rect 190794 -7964 191414 -3132
rect 195294 708028 195914 711900
rect 195294 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 195914 708028
rect 195294 707708 195914 707792
rect 195294 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 195914 707708
rect 195294 700954 195914 707472
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3536 195914 16398
rect 195294 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 195914 -3536
rect 195294 -3856 195914 -3772
rect 195294 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 195914 -3856
rect 195294 -7964 195914 -4092
rect 199794 708988 200414 711900
rect 199794 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 200414 708988
rect 199794 708668 200414 708752
rect 199794 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 200414 708668
rect 199794 669454 200414 708432
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4496 200414 20898
rect 199794 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 200414 -4496
rect 199794 -4816 200414 -4732
rect 199794 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 200414 -4816
rect 199794 -7964 200414 -5052
rect 204294 709948 204914 711900
rect 204294 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 204914 709948
rect 204294 709628 204914 709712
rect 204294 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 204914 709628
rect 204294 673954 204914 709392
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5456 204914 25398
rect 204294 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 204914 -5456
rect 204294 -5776 204914 -5692
rect 204294 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 204914 -5776
rect 204294 -7964 204914 -6012
rect 208794 710908 209414 711900
rect 208794 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 209414 710908
rect 208794 710588 209414 710672
rect 208794 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 209414 710588
rect 208794 678454 209414 710352
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6416 209414 29898
rect 208794 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 209414 -6416
rect 208794 -6736 209414 -6652
rect 208794 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 209414 -6736
rect 208794 -7964 209414 -6972
rect 213294 711868 213914 711900
rect 213294 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 213914 711868
rect 213294 711548 213914 711632
rect 213294 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 213914 711548
rect 213294 682954 213914 711312
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 705148 218414 711900
rect 217794 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 218414 705148
rect 217794 704828 218414 704912
rect 217794 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 218414 704828
rect 217794 687454 218414 704592
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 706108 222914 711900
rect 222294 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 222914 706108
rect 222294 705788 222914 705872
rect 222294 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 222914 705788
rect 222294 691954 222914 705552
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 707068 227414 711900
rect 226794 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 227414 707068
rect 226794 706748 227414 706832
rect 226794 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 227414 706748
rect 226794 696454 227414 706512
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 708028 231914 711900
rect 231294 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 231914 708028
rect 231294 707708 231914 707792
rect 231294 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 231914 707708
rect 231294 700954 231914 707472
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708988 236414 711900
rect 235794 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 236414 708988
rect 235794 708668 236414 708752
rect 235794 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 236414 708668
rect 235794 669454 236414 708432
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709948 240914 711900
rect 240294 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 240914 709948
rect 240294 709628 240914 709712
rect 240294 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 240914 709628
rect 240294 673954 240914 709392
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710908 245414 711900
rect 244794 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 245414 710908
rect 244794 710588 245414 710672
rect 244794 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 245414 710588
rect 244794 678454 245414 710352
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711868 249914 711900
rect 249294 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 249914 711868
rect 249294 711548 249914 711632
rect 249294 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 249914 711548
rect 249294 682954 249914 711312
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 705148 254414 711900
rect 253794 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 254414 705148
rect 253794 704828 254414 704912
rect 253794 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 254414 704828
rect 253794 687454 254414 704592
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 706108 258914 711900
rect 258294 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 258914 706108
rect 258294 705788 258914 705872
rect 258294 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 258914 705788
rect 258294 691954 258914 705552
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 707068 263414 711900
rect 262794 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 263414 707068
rect 262794 706748 263414 706832
rect 262794 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 263414 706748
rect 262794 696454 263414 706512
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 708028 267914 711900
rect 267294 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 267914 708028
rect 267294 707708 267914 707792
rect 267294 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 267914 707708
rect 267294 700954 267914 707472
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708988 272414 711900
rect 271794 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 272414 708988
rect 271794 708668 272414 708752
rect 271794 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 272414 708668
rect 271794 669454 272414 708432
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709948 276914 711900
rect 276294 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 276914 709948
rect 276294 709628 276914 709712
rect 276294 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 276914 709628
rect 276294 673954 276914 709392
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710908 281414 711900
rect 280794 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 281414 710908
rect 280794 710588 281414 710672
rect 280794 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 281414 710588
rect 280794 678454 281414 710352
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711868 285914 711900
rect 285294 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 285914 711868
rect 285294 711548 285914 711632
rect 285294 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 285914 711548
rect 285294 682954 285914 711312
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 705148 290414 711900
rect 289794 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 290414 705148
rect 289794 704828 290414 704912
rect 289794 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 290414 704828
rect 289794 687454 290414 704592
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 706108 294914 711900
rect 294294 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 294914 706108
rect 294294 705788 294914 705872
rect 294294 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 294914 705788
rect 294294 691954 294914 705552
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 707068 299414 711900
rect 298794 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 299414 707068
rect 298794 706748 299414 706832
rect 298794 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 299414 706748
rect 298794 696454 299414 706512
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 708028 303914 711900
rect 303294 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 303914 708028
rect 303294 707708 303914 707792
rect 303294 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 303914 707708
rect 303294 700954 303914 707472
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708988 308414 711900
rect 307794 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 308414 708988
rect 307794 708668 308414 708752
rect 307794 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 308414 708668
rect 307794 669454 308414 708432
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709948 312914 711900
rect 312294 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 312914 709948
rect 312294 709628 312914 709712
rect 312294 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 312914 709628
rect 312294 673954 312914 709392
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710908 317414 711900
rect 316794 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 317414 710908
rect 316794 710588 317414 710672
rect 316794 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 317414 710588
rect 316794 678454 317414 710352
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711868 321914 711900
rect 321294 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 321914 711868
rect 321294 711548 321914 711632
rect 321294 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 321914 711548
rect 321294 682954 321914 711312
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 705148 326414 711900
rect 325794 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 326414 705148
rect 325794 704828 326414 704912
rect 325794 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 326414 704828
rect 325794 687454 326414 704592
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 706108 330914 711900
rect 330294 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 330914 706108
rect 330294 705788 330914 705872
rect 330294 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 330914 705788
rect 330294 691954 330914 705552
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 707068 335414 711900
rect 334794 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 335414 707068
rect 334794 706748 335414 706832
rect 334794 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 335414 706748
rect 334794 696454 335414 706512
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 708028 339914 711900
rect 339294 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 339914 708028
rect 339294 707708 339914 707792
rect 339294 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 339914 707708
rect 339294 700954 339914 707472
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708988 344414 711900
rect 343794 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 344414 708988
rect 343794 708668 344414 708752
rect 343794 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 344414 708668
rect 343794 669454 344414 708432
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709948 348914 711900
rect 348294 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 348914 709948
rect 348294 709628 348914 709712
rect 348294 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 348914 709628
rect 348294 673954 348914 709392
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710908 353414 711900
rect 352794 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 353414 710908
rect 352794 710588 353414 710672
rect 352794 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 353414 710588
rect 352794 678454 353414 710352
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711868 357914 711900
rect 357294 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 357914 711868
rect 357294 711548 357914 711632
rect 357294 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 357914 711548
rect 357294 682954 357914 711312
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 705148 362414 711900
rect 361794 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 362414 705148
rect 361794 704828 362414 704912
rect 361794 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 362414 704828
rect 361794 687454 362414 704592
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 236056 479710 236194 479770
rect 237144 479710 237298 479770
rect 238232 479710 238402 479770
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 214603 444820 214669 444821
rect 214603 444756 214604 444820
rect 214668 444756 214669 444820
rect 214603 444755 214669 444756
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 214419 284884 214485 284885
rect 214419 284820 214420 284884
rect 214484 284820 214485 284884
rect 214419 284819 214485 284820
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7376 213914 34398
rect 214422 3365 214482 284819
rect 214606 162893 214666 444755
rect 216075 441692 216141 441693
rect 216075 441628 216076 441692
rect 216140 441628 216141 441692
rect 216075 441627 216141 441628
rect 215155 303244 215221 303245
rect 215155 303180 215156 303244
rect 215220 303180 215221 303244
rect 215155 303179 215221 303180
rect 214603 162892 214669 162893
rect 214603 162828 214604 162892
rect 214668 162828 214669 162892
rect 214603 162827 214669 162828
rect 215158 3501 215218 303179
rect 215891 269788 215957 269789
rect 215891 269724 215892 269788
rect 215956 269724 215957 269788
rect 215891 269723 215957 269724
rect 215894 3637 215954 269723
rect 216078 187781 216138 441627
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217179 305828 217245 305829
rect 217179 305764 217180 305828
rect 217244 305764 217245 305828
rect 217179 305763 217245 305764
rect 216259 303108 216325 303109
rect 216259 303044 216260 303108
rect 216324 303044 216325 303108
rect 216259 303043 216325 303044
rect 216075 187780 216141 187781
rect 216075 187716 216076 187780
rect 216140 187716 216141 187780
rect 216075 187715 216141 187716
rect 216262 158405 216322 303043
rect 216995 301476 217061 301477
rect 216995 301412 216996 301476
rect 217060 301412 217061 301476
rect 216995 301411 217061 301412
rect 216443 254556 216509 254557
rect 216443 254492 216444 254556
rect 216508 254492 216509 254556
rect 216443 254491 216509 254492
rect 216259 158404 216325 158405
rect 216259 158340 216260 158404
rect 216324 158340 216325 158404
rect 216259 158339 216325 158340
rect 215891 3636 215957 3637
rect 215891 3572 215892 3636
rect 215956 3572 215957 3636
rect 215891 3571 215957 3572
rect 216446 3501 216506 254491
rect 216998 155549 217058 301411
rect 217182 158133 217242 305763
rect 217363 305692 217429 305693
rect 217363 305628 217364 305692
rect 217428 305628 217429 305692
rect 217363 305627 217429 305628
rect 217179 158132 217245 158133
rect 217179 158068 217180 158132
rect 217244 158068 217245 158132
rect 217179 158067 217245 158068
rect 217366 157997 217426 305627
rect 217794 291454 218414 326898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 218835 306100 218901 306101
rect 218835 306036 218836 306100
rect 218900 306036 218901 306100
rect 218835 306035 218901 306036
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217547 250476 217613 250477
rect 217547 250412 217548 250476
rect 217612 250412 217613 250476
rect 217547 250411 217613 250412
rect 217363 157996 217429 157997
rect 217363 157932 217364 157996
rect 217428 157932 217429 157996
rect 217363 157931 217429 157932
rect 216995 155548 217061 155549
rect 216995 155484 216996 155548
rect 217060 155484 217061 155548
rect 216995 155483 217061 155484
rect 217550 3501 217610 250411
rect 217794 245308 218414 254898
rect 218651 243540 218717 243541
rect 218651 243476 218652 243540
rect 218716 243476 218717 243540
rect 218651 243475 218717 243476
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 215155 3500 215221 3501
rect 215155 3436 215156 3500
rect 215220 3436 215221 3500
rect 215155 3435 215221 3436
rect 216443 3500 216509 3501
rect 216443 3436 216444 3500
rect 216508 3436 216509 3500
rect 216443 3435 216509 3436
rect 217547 3500 217613 3501
rect 217547 3436 217548 3500
rect 217612 3436 217613 3500
rect 217547 3435 217613 3436
rect 217794 3454 218414 38898
rect 218654 3501 218714 243475
rect 218838 158677 218898 306035
rect 219019 305964 219085 305965
rect 219019 305900 219020 305964
rect 219084 305900 219085 305964
rect 219019 305899 219085 305900
rect 218835 158676 218901 158677
rect 218835 158612 218836 158676
rect 218900 158612 218901 158676
rect 218835 158611 218901 158612
rect 219022 158541 219082 305899
rect 219203 301748 219269 301749
rect 219203 301684 219204 301748
rect 219268 301684 219269 301748
rect 219203 301683 219269 301684
rect 219019 158540 219085 158541
rect 219019 158476 219020 158540
rect 219084 158476 219085 158540
rect 219019 158475 219085 158476
rect 219206 3637 219266 301683
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 236134 476781 236194 479710
rect 236131 476780 236197 476781
rect 236131 476716 236132 476780
rect 236196 476716 236197 476780
rect 236131 476715 236197 476716
rect 237238 476237 237298 479710
rect 238342 477325 238402 479710
rect 238339 477324 238405 477325
rect 238339 477260 238340 477324
rect 238404 477260 238405 477324
rect 238339 477259 238405 477260
rect 239630 476917 239690 479710
rect 240550 476917 240610 479710
rect 241838 477189 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 245440 479710 245578 479770
rect 246528 479710 246682 479770
rect 247616 479710 247786 479770
rect 241835 477188 241901 477189
rect 241835 477124 241836 477188
rect 241900 477124 241901 477188
rect 241835 477123 241901 477124
rect 239627 476916 239693 476917
rect 239627 476852 239628 476916
rect 239692 476852 239693 476916
rect 239627 476851 239693 476852
rect 240547 476916 240613 476917
rect 240547 476852 240548 476916
rect 240612 476852 240613 476916
rect 240547 476851 240613 476852
rect 243126 476237 243186 479710
rect 244230 476373 244290 479710
rect 244227 476372 244293 476373
rect 244227 476308 244228 476372
rect 244292 476308 244293 476372
rect 244227 476307 244293 476308
rect 245518 476237 245578 479710
rect 246622 476237 246682 479710
rect 247726 476373 247786 479710
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 250064 479710 250178 479770
rect 250744 479710 250914 479770
rect 251288 479710 251466 479770
rect 247723 476372 247789 476373
rect 247723 476308 247724 476372
rect 247788 476308 247789 476372
rect 247723 476307 247789 476308
rect 248278 476237 248338 479710
rect 248646 476237 248706 479710
rect 250118 476373 250178 479710
rect 250115 476372 250181 476373
rect 250115 476308 250116 476372
rect 250180 476308 250181 476372
rect 250115 476307 250181 476308
rect 250854 476237 250914 479710
rect 251406 476373 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 251403 476372 251469 476373
rect 251403 476308 251404 476372
rect 251468 476308 251469 476372
rect 251403 476307 251469 476308
rect 252326 476237 252386 479710
rect 253430 476509 253490 479710
rect 253427 476508 253493 476509
rect 253427 476444 253428 476508
rect 253492 476444 253493 476508
rect 253427 476443 253493 476444
rect 253614 476237 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 254534 476237 254594 479710
rect 255822 476237 255882 479710
rect 256190 477053 256250 479710
rect 256187 477052 256253 477053
rect 256187 476988 256188 477052
rect 256252 476988 256253 477052
rect 256187 476987 256253 476988
rect 257110 476237 257170 479710
rect 257846 479710 258148 479770
rect 258496 479770 258556 480080
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 258496 479710 258642 479770
rect 259448 479710 259562 479770
rect 257846 476778 257906 479710
rect 258027 476780 258093 476781
rect 258027 476778 258028 476780
rect 257846 476718 258028 476778
rect 258027 476716 258028 476718
rect 258092 476716 258093 476780
rect 258027 476715 258093 476716
rect 258582 476237 258642 479710
rect 259502 476373 259562 479710
rect 260606 479710 260732 479770
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 261080 479710 261218 479770
rect 259499 476372 259565 476373
rect 259499 476308 259500 476372
rect 259564 476308 259565 476372
rect 259499 476307 259565 476308
rect 260606 476237 260666 479710
rect 261158 476509 261218 479710
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 261155 476508 261221 476509
rect 261155 476444 261156 476508
rect 261220 476444 261221 476508
rect 261155 476443 261221 476444
rect 261710 476237 261770 479710
rect 262814 476237 262874 479710
rect 263550 476781 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476780 263613 476781
rect 263547 476716 263548 476780
rect 263612 476716 263613 476780
rect 263547 476715 263613 476716
rect 263918 476237 263978 479710
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 476645 266002 479710
rect 265939 476644 266005 476645
rect 265939 476580 265940 476644
rect 266004 476580 266005 476644
rect 265939 476579 266005 476580
rect 266494 476373 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 266491 476372 266557 476373
rect 266491 476308 266492 476372
rect 266556 476308 266557 476372
rect 266491 476307 266557 476308
rect 267598 476237 267658 479710
rect 268334 476373 268394 479710
rect 268331 476372 268397 476373
rect 268331 476308 268332 476372
rect 268396 476308 268397 476372
rect 268331 476307 268397 476308
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 271144 479710 271338 479770
rect 270910 476645 270970 479710
rect 270907 476644 270973 476645
rect 270907 476580 270908 476644
rect 270972 476580 270973 476644
rect 270907 476579 270973 476580
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 273592 479710 273730 479770
rect 272198 476237 272258 479710
rect 273302 476237 273362 479710
rect 273670 476373 273730 479710
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 274406 476509 274466 479710
rect 274403 476508 274469 476509
rect 274403 476444 274404 476508
rect 274468 476444 274469 476508
rect 274403 476443 274469 476444
rect 273667 476372 273733 476373
rect 273667 476308 273668 476372
rect 273732 476308 273733 476372
rect 273667 476307 273733 476308
rect 275878 476237 275938 479710
rect 276062 476373 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476372 276125 476373
rect 276059 476308 276060 476372
rect 276124 476308 276125 476372
rect 276059 476307 276125 476308
rect 276982 476237 277042 479710
rect 278086 476373 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 279168 479710 279250 479770
rect 280936 479710 281090 479770
rect 283520 479710 283666 479770
rect 285968 479710 286058 479770
rect 278083 476372 278149 476373
rect 278083 476308 278084 476372
rect 278148 476308 278149 476372
rect 278083 476307 278149 476308
rect 278454 476237 278514 479710
rect 279190 476237 279250 479710
rect 281030 476237 281090 479710
rect 283606 476237 283666 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293448 479770 293508 480080
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 293448 479710 293602 479770
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293542 476237 293602 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 305960 479710 306114 479770
rect 308544 479710 308690 479770
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476237 303538 479710
rect 306054 476237 306114 479710
rect 308630 476781 308690 479710
rect 308627 476780 308693 476781
rect 308627 476716 308628 476780
rect 308692 476716 308693 476780
rect 308627 476715 308693 476716
rect 311022 476373 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318472 479770 318532 480080
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 318472 479710 318626 479770
rect 320920 479710 321018 479770
rect 313414 476781 313474 479710
rect 313411 476780 313477 476781
rect 313411 476716 313412 476780
rect 313476 476716 313477 476780
rect 313411 476715 313477 476716
rect 311019 476372 311085 476373
rect 311019 476308 311020 476372
rect 311084 476308 311085 476372
rect 311019 476307 311085 476308
rect 315806 476237 315866 479710
rect 318566 476509 318626 479710
rect 318563 476508 318629 476509
rect 318563 476444 318564 476508
rect 318628 476444 318629 476508
rect 318563 476443 318629 476444
rect 320958 476237 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 476237 323410 479710
rect 325926 476509 325986 479710
rect 325923 476508 325989 476509
rect 325923 476444 325924 476508
rect 325988 476444 325989 476508
rect 325923 476443 325989 476444
rect 237235 476236 237301 476237
rect 237235 476172 237236 476236
rect 237300 476172 237301 476236
rect 237235 476171 237301 476172
rect 243123 476236 243189 476237
rect 243123 476172 243124 476236
rect 243188 476172 243189 476236
rect 243123 476171 243189 476172
rect 245515 476236 245581 476237
rect 245515 476172 245516 476236
rect 245580 476172 245581 476236
rect 245515 476171 245581 476172
rect 246619 476236 246685 476237
rect 246619 476172 246620 476236
rect 246684 476172 246685 476236
rect 246619 476171 246685 476172
rect 248275 476236 248341 476237
rect 248275 476172 248276 476236
rect 248340 476172 248341 476236
rect 248275 476171 248341 476172
rect 248643 476236 248709 476237
rect 248643 476172 248644 476236
rect 248708 476172 248709 476236
rect 248643 476171 248709 476172
rect 250851 476236 250917 476237
rect 250851 476172 250852 476236
rect 250916 476172 250917 476236
rect 250851 476171 250917 476172
rect 252323 476236 252389 476237
rect 252323 476172 252324 476236
rect 252388 476172 252389 476236
rect 252323 476171 252389 476172
rect 253611 476236 253677 476237
rect 253611 476172 253612 476236
rect 253676 476172 253677 476236
rect 253611 476171 253677 476172
rect 254531 476236 254597 476237
rect 254531 476172 254532 476236
rect 254596 476172 254597 476236
rect 254531 476171 254597 476172
rect 255819 476236 255885 476237
rect 255819 476172 255820 476236
rect 255884 476172 255885 476236
rect 255819 476171 255885 476172
rect 257107 476236 257173 476237
rect 257107 476172 257108 476236
rect 257172 476172 257173 476236
rect 257107 476171 257173 476172
rect 258579 476236 258645 476237
rect 258579 476172 258580 476236
rect 258644 476172 258645 476236
rect 258579 476171 258645 476172
rect 260603 476236 260669 476237
rect 260603 476172 260604 476236
rect 260668 476172 260669 476236
rect 260603 476171 260669 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 262811 476236 262877 476237
rect 262811 476172 262812 476236
rect 262876 476172 262877 476236
rect 262811 476171 262877 476172
rect 263915 476236 263981 476237
rect 263915 476172 263916 476236
rect 263980 476172 263981 476236
rect 263915 476171 263981 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 267595 476236 267661 476237
rect 267595 476172 267596 476236
rect 267660 476172 267661 476236
rect 267595 476171 267661 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 273299 476236 273365 476237
rect 273299 476172 273300 476236
rect 273364 476172 273365 476236
rect 273299 476171 273365 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278451 476236 278517 476237
rect 278451 476172 278452 476236
rect 278516 476172 278517 476236
rect 278451 476171 278517 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 281027 476236 281093 476237
rect 281027 476172 281028 476236
rect 281092 476172 281093 476236
rect 281027 476171 281093 476172
rect 283603 476236 283669 476237
rect 283603 476172 283604 476236
rect 283668 476172 283669 476236
rect 283603 476171 283669 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293539 476236 293605 476237
rect 293539 476172 293540 476236
rect 293604 476172 293605 476236
rect 293539 476171 293605 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 303475 476236 303541 476237
rect 303475 476172 303476 476236
rect 303540 476172 303541 476236
rect 303475 476171 303541 476172
rect 306051 476236 306117 476237
rect 306051 476172 306052 476236
rect 306116 476172 306117 476236
rect 306051 476171 306117 476172
rect 315803 476236 315869 476237
rect 315803 476172 315804 476236
rect 315868 476172 315869 476236
rect 315803 476171 315869 476172
rect 320955 476236 321021 476237
rect 320955 476172 320956 476236
rect 321020 476172 321021 476236
rect 320955 476171 321021 476172
rect 323347 476236 323413 476237
rect 323347 476172 323348 476236
rect 323412 476172 323413 476236
rect 323347 476171 323413 476172
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 443544 362414 470898
rect 366294 706108 366914 711900
rect 366294 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 366914 706108
rect 366294 705788 366914 705872
rect 366294 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 366914 705788
rect 366294 691954 366914 705552
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 365115 445772 365181 445773
rect 365115 445708 365116 445772
rect 365180 445708 365181 445772
rect 365115 445707 365181 445708
rect 364931 444684 364997 444685
rect 364931 444620 364932 444684
rect 364996 444620 364997 444684
rect 364931 444619 364997 444620
rect 236608 435454 236928 435486
rect 236608 435218 236650 435454
rect 236886 435218 236928 435454
rect 236608 435134 236928 435218
rect 236608 434898 236650 435134
rect 236886 434898 236928 435134
rect 236608 434866 236928 434898
rect 267328 435454 267648 435486
rect 267328 435218 267370 435454
rect 267606 435218 267648 435454
rect 267328 435134 267648 435218
rect 267328 434898 267370 435134
rect 267606 434898 267648 435134
rect 267328 434866 267648 434898
rect 298048 435454 298368 435486
rect 298048 435218 298090 435454
rect 298326 435218 298368 435454
rect 298048 435134 298368 435218
rect 298048 434898 298090 435134
rect 298326 434898 298368 435134
rect 298048 434866 298368 434898
rect 328768 435454 329088 435486
rect 328768 435218 328810 435454
rect 329046 435218 329088 435454
rect 328768 435134 329088 435218
rect 328768 434898 328810 435134
rect 329046 434898 329088 435134
rect 328768 434866 329088 434898
rect 359488 435454 359808 435486
rect 359488 435218 359530 435454
rect 359766 435218 359808 435454
rect 359488 435134 359808 435218
rect 359488 434898 359530 435134
rect 359766 434898 359808 435134
rect 359488 434866 359808 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 251968 403954 252288 403986
rect 251968 403718 252010 403954
rect 252246 403718 252288 403954
rect 251968 403634 252288 403718
rect 251968 403398 252010 403634
rect 252246 403398 252288 403634
rect 251968 403366 252288 403398
rect 282688 403954 283008 403986
rect 282688 403718 282730 403954
rect 282966 403718 283008 403954
rect 282688 403634 283008 403718
rect 282688 403398 282730 403634
rect 282966 403398 283008 403634
rect 282688 403366 283008 403398
rect 313408 403954 313728 403986
rect 313408 403718 313450 403954
rect 313686 403718 313728 403954
rect 313408 403634 313728 403718
rect 313408 403398 313450 403634
rect 313686 403398 313728 403634
rect 313408 403366 313728 403398
rect 344128 403954 344448 403986
rect 344128 403718 344170 403954
rect 344406 403718 344448 403954
rect 344128 403634 344448 403718
rect 344128 403398 344170 403634
rect 344406 403398 344448 403634
rect 344128 403366 344448 403398
rect 236608 399454 236928 399486
rect 236608 399218 236650 399454
rect 236886 399218 236928 399454
rect 236608 399134 236928 399218
rect 236608 398898 236650 399134
rect 236886 398898 236928 399134
rect 236608 398866 236928 398898
rect 267328 399454 267648 399486
rect 267328 399218 267370 399454
rect 267606 399218 267648 399454
rect 267328 399134 267648 399218
rect 267328 398898 267370 399134
rect 267606 398898 267648 399134
rect 267328 398866 267648 398898
rect 298048 399454 298368 399486
rect 298048 399218 298090 399454
rect 298326 399218 298368 399454
rect 298048 399134 298368 399218
rect 298048 398898 298090 399134
rect 298326 398898 298368 399134
rect 298048 398866 298368 398898
rect 328768 399454 329088 399486
rect 328768 399218 328810 399454
rect 329046 399218 329088 399454
rect 328768 399134 329088 399218
rect 328768 398898 328810 399134
rect 329046 398898 329088 399134
rect 328768 398866 329088 398898
rect 359488 399454 359808 399486
rect 359488 399218 359530 399454
rect 359766 399218 359808 399454
rect 359488 399134 359808 399218
rect 359488 398898 359530 399134
rect 359766 398898 359808 399134
rect 359488 398866 359808 398898
rect 232083 374100 232149 374101
rect 232083 374036 232084 374100
rect 232148 374036 232149 374100
rect 232083 374035 232149 374036
rect 232086 373010 232146 374035
rect 232086 372950 232698 373010
rect 232083 372740 232149 372741
rect 232083 372676 232084 372740
rect 232148 372676 232149 372740
rect 232083 372675 232149 372676
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 232086 364350 232146 372675
rect 232086 364290 232514 364350
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 232454 308685 232514 364290
rect 232638 309773 232698 372950
rect 251968 367954 252288 367986
rect 251968 367718 252010 367954
rect 252246 367718 252288 367954
rect 251968 367634 252288 367718
rect 251968 367398 252010 367634
rect 252246 367398 252288 367634
rect 251968 367366 252288 367398
rect 282688 367954 283008 367986
rect 282688 367718 282730 367954
rect 282966 367718 283008 367954
rect 282688 367634 283008 367718
rect 282688 367398 282730 367634
rect 282966 367398 283008 367634
rect 282688 367366 283008 367398
rect 313408 367954 313728 367986
rect 313408 367718 313450 367954
rect 313686 367718 313728 367954
rect 313408 367634 313728 367718
rect 313408 367398 313450 367634
rect 313686 367398 313728 367634
rect 313408 367366 313728 367398
rect 344128 367954 344448 367986
rect 344128 367718 344170 367954
rect 344406 367718 344448 367954
rect 344128 367634 344448 367718
rect 344128 367398 344170 367634
rect 344406 367398 344448 367634
rect 344128 367366 344448 367398
rect 236608 363454 236928 363486
rect 236608 363218 236650 363454
rect 236886 363218 236928 363454
rect 236608 363134 236928 363218
rect 236608 362898 236650 363134
rect 236886 362898 236928 363134
rect 236608 362866 236928 362898
rect 267328 363454 267648 363486
rect 267328 363218 267370 363454
rect 267606 363218 267648 363454
rect 267328 363134 267648 363218
rect 267328 362898 267370 363134
rect 267606 362898 267648 363134
rect 267328 362866 267648 362898
rect 298048 363454 298368 363486
rect 298048 363218 298090 363454
rect 298326 363218 298368 363454
rect 298048 363134 298368 363218
rect 298048 362898 298090 363134
rect 298326 362898 298368 363134
rect 298048 362866 298368 362898
rect 328768 363454 329088 363486
rect 328768 363218 328810 363454
rect 329046 363218 329088 363454
rect 328768 363134 329088 363218
rect 328768 362898 328810 363134
rect 329046 362898 329088 363134
rect 328768 362866 329088 362898
rect 359488 363454 359808 363486
rect 359488 363218 359530 363454
rect 359766 363218 359808 363454
rect 359488 363134 359808 363218
rect 359488 362898 359530 363134
rect 359766 362898 359808 363134
rect 359488 362866 359808 362898
rect 251968 331954 252288 331986
rect 251968 331718 252010 331954
rect 252246 331718 252288 331954
rect 251968 331634 252288 331718
rect 251968 331398 252010 331634
rect 252246 331398 252288 331634
rect 251968 331366 252288 331398
rect 282688 331954 283008 331986
rect 282688 331718 282730 331954
rect 282966 331718 283008 331954
rect 282688 331634 283008 331718
rect 282688 331398 282730 331634
rect 282966 331398 283008 331634
rect 282688 331366 283008 331398
rect 313408 331954 313728 331986
rect 313408 331718 313450 331954
rect 313686 331718 313728 331954
rect 313408 331634 313728 331718
rect 313408 331398 313450 331634
rect 313686 331398 313728 331634
rect 313408 331366 313728 331398
rect 344128 331954 344448 331986
rect 344128 331718 344170 331954
rect 344406 331718 344448 331954
rect 344128 331634 344448 331718
rect 344128 331398 344170 331634
rect 344406 331398 344448 331634
rect 344128 331366 344448 331398
rect 236608 327454 236928 327486
rect 236608 327218 236650 327454
rect 236886 327218 236928 327454
rect 236608 327134 236928 327218
rect 236608 326898 236650 327134
rect 236886 326898 236928 327134
rect 236608 326866 236928 326898
rect 267328 327454 267648 327486
rect 267328 327218 267370 327454
rect 267606 327218 267648 327454
rect 267328 327134 267648 327218
rect 267328 326898 267370 327134
rect 267606 326898 267648 327134
rect 267328 326866 267648 326898
rect 298048 327454 298368 327486
rect 298048 327218 298090 327454
rect 298326 327218 298368 327454
rect 298048 327134 298368 327218
rect 298048 326898 298090 327134
rect 298326 326898 298368 327134
rect 298048 326866 298368 326898
rect 328768 327454 329088 327486
rect 328768 327218 328810 327454
rect 329046 327218 329088 327454
rect 328768 327134 329088 327218
rect 328768 326898 328810 327134
rect 329046 326898 329088 327134
rect 328768 326866 329088 326898
rect 359488 327454 359808 327486
rect 359488 327218 359530 327454
rect 359766 327218 359808 327454
rect 359488 327134 359808 327218
rect 359488 326898 359530 327134
rect 359766 326898 359808 327134
rect 359488 326866 359808 326898
rect 232819 310724 232885 310725
rect 232819 310660 232820 310724
rect 232884 310660 232885 310724
rect 232819 310659 232885 310660
rect 232822 310453 232882 310659
rect 232819 310452 232885 310453
rect 232819 310388 232820 310452
rect 232884 310388 232885 310452
rect 232819 310387 232885 310388
rect 232635 309772 232701 309773
rect 232635 309708 232636 309772
rect 232700 309708 232701 309772
rect 232635 309707 232701 309708
rect 232451 308684 232517 308685
rect 232451 308620 232452 308684
rect 232516 308620 232517 308684
rect 232451 308619 232517 308620
rect 359963 308548 360029 308549
rect 359963 308484 359964 308548
rect 360028 308484 360029 308548
rect 359963 308483 360029 308484
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 245308 245414 245898
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 245308 249914 250398
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 245308 254414 254898
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 245308 258914 259398
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 245308 263414 263898
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 245308 267914 268398
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 245308 281414 245898
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 245308 285914 250398
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 245308 290414 254898
rect 294294 295954 294914 308400
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 245308 294914 259398
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 358123 306508 358189 306509
rect 358123 306444 358124 306508
rect 358188 306444 358189 306508
rect 358123 306443 358189 306444
rect 358126 304333 358186 306443
rect 358123 304332 358189 304333
rect 358123 304268 358124 304332
rect 358188 304268 358189 304332
rect 358123 304267 358189 304268
rect 359966 302250 360026 308483
rect 359966 302190 360210 302250
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 358859 251020 358925 251021
rect 358859 250956 358860 251020
rect 358924 250956 358925 251020
rect 358859 250955 358925 250956
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 358307 250612 358373 250613
rect 358307 250548 358308 250612
rect 358372 250548 358373 250612
rect 358307 250547 358373 250548
rect 357294 245308 357914 250398
rect 358123 248028 358189 248029
rect 358123 247964 358124 248028
rect 358188 247964 358189 248028
rect 358123 247963 358189 247964
rect 357571 243540 357637 243541
rect 357571 243476 357572 243540
rect 357636 243476 357637 243540
rect 357571 243475 357637 243476
rect 220272 223954 220620 223986
rect 220272 223718 220328 223954
rect 220564 223718 220620 223954
rect 220272 223634 220620 223718
rect 220272 223398 220328 223634
rect 220564 223398 220620 223634
rect 220272 223366 220620 223398
rect 356000 223954 356348 223986
rect 356000 223718 356056 223954
rect 356292 223718 356348 223954
rect 356000 223634 356348 223718
rect 356000 223398 356056 223634
rect 356292 223398 356348 223634
rect 356000 223366 356348 223398
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 187954 220620 187986
rect 220272 187718 220328 187954
rect 220564 187718 220620 187954
rect 220272 187634 220620 187718
rect 220272 187398 220328 187634
rect 220564 187398 220620 187634
rect 220272 187366 220620 187398
rect 356000 187954 356348 187986
rect 356000 187718 356056 187954
rect 356292 187718 356348 187954
rect 356000 187634 356348 187718
rect 356000 187398 356056 187634
rect 356292 187398 356348 187634
rect 356000 187366 356348 187398
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 356835 160172 356901 160173
rect 356835 160108 356836 160172
rect 356900 160108 356901 160172
rect 356835 160107 356901 160108
rect 236056 159490 236116 160106
rect 237144 159490 237204 160106
rect 238232 159490 238292 160106
rect 236056 159430 236194 159490
rect 237144 159430 237298 159490
rect 236134 158949 236194 159430
rect 236131 158948 236197 158949
rect 236131 158884 236132 158948
rect 236196 158884 236197 158948
rect 236131 158883 236197 158884
rect 237238 158813 237298 159430
rect 238158 159430 238292 159490
rect 239592 159490 239652 160106
rect 240544 159490 240604 160106
rect 241768 159490 241828 160106
rect 243128 159490 243188 160106
rect 239592 159430 239690 159490
rect 240544 159430 240610 159490
rect 241768 159430 241898 159490
rect 237235 158812 237301 158813
rect 237235 158748 237236 158812
rect 237300 158748 237301 158812
rect 237235 158747 237301 158748
rect 238158 158677 238218 159430
rect 239630 158677 239690 159430
rect 240550 158677 240610 159430
rect 238155 158676 238221 158677
rect 238155 158612 238156 158676
rect 238220 158612 238221 158676
rect 238155 158611 238221 158612
rect 239627 158676 239693 158677
rect 239627 158612 239628 158676
rect 239692 158612 239693 158676
rect 239627 158611 239693 158612
rect 240547 158676 240613 158677
rect 240547 158612 240548 158676
rect 240612 158612 240613 158676
rect 240547 158611 240613 158612
rect 241838 158541 241898 159430
rect 243126 159430 243188 159490
rect 244216 159490 244276 160106
rect 245440 159490 245500 160106
rect 246528 159490 246588 160106
rect 247616 159490 247676 160106
rect 248296 159490 248356 160106
rect 248704 159490 248764 160106
rect 244216 159430 244290 159490
rect 245440 159430 245578 159490
rect 246528 159430 246682 159490
rect 247616 159430 247786 159490
rect 243126 159085 243186 159430
rect 243123 159084 243189 159085
rect 243123 159020 243124 159084
rect 243188 159020 243189 159084
rect 243123 159019 243189 159020
rect 241835 158540 241901 158541
rect 241835 158476 241836 158540
rect 241900 158476 241901 158540
rect 241835 158475 241901 158476
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 219203 3636 219269 3637
rect 219203 3572 219204 3636
rect 219268 3572 219269 3636
rect 219203 3571 219269 3572
rect 214419 3364 214485 3365
rect 214419 3300 214420 3364
rect 214484 3300 214485 3364
rect 214419 3299 214485 3300
rect 213294 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 213914 -7376
rect 213294 -7696 213914 -7612
rect 213294 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 213914 -7696
rect 213294 -7964 213914 -7932
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 218651 3500 218717 3501
rect 218651 3436 218652 3500
rect 218716 3436 218717 3500
rect 218651 3435 218717 3436
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -656 218414 2898
rect 217794 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 218414 -656
rect 217794 -976 218414 -892
rect 217794 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 218414 -976
rect 217794 -7964 218414 -1212
rect 222294 -1616 222914 7398
rect 222294 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 222914 -1616
rect 222294 -1936 222914 -1852
rect 222294 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 222914 -1936
rect 222294 -7964 222914 -2172
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2576 227414 11898
rect 226794 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 227414 -2576
rect 226794 -2896 227414 -2812
rect 226794 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 227414 -2896
rect 226794 -7964 227414 -3132
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3536 231914 16398
rect 231294 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 231914 -3536
rect 231294 -3856 231914 -3772
rect 231294 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 231914 -3856
rect 231294 -7964 231914 -4092
rect 235794 129454 236414 158000
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4496 236414 20898
rect 235794 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 236414 -4496
rect 235794 -4816 236414 -4732
rect 235794 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 236414 -4816
rect 235794 -7964 236414 -5052
rect 240294 133954 240914 158000
rect 244230 157453 244290 159430
rect 244227 157452 244293 157453
rect 244227 157388 244228 157452
rect 244292 157388 244293 157452
rect 244227 157387 244293 157388
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5456 240914 25398
rect 240294 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 240914 -5456
rect 240294 -5776 240914 -5692
rect 240294 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 240914 -5776
rect 240294 -7964 240914 -6012
rect 244794 138454 245414 158000
rect 245518 157453 245578 159430
rect 246622 158133 246682 159430
rect 246619 158132 246685 158133
rect 246619 158068 246620 158132
rect 246684 158068 246685 158132
rect 246619 158067 246685 158068
rect 245515 157452 245581 157453
rect 245515 157388 245516 157452
rect 245580 157388 245581 157452
rect 245515 157387 245581 157388
rect 247726 157045 247786 159430
rect 248278 159430 248356 159490
rect 248646 159430 248764 159490
rect 250064 159490 250124 160106
rect 250744 159490 250804 160106
rect 251288 159490 251348 160106
rect 252376 159490 252436 160106
rect 253464 159490 253524 160106
rect 250064 159430 250178 159490
rect 250744 159430 250914 159490
rect 251288 159430 251466 159490
rect 248278 158677 248338 159430
rect 248275 158676 248341 158677
rect 248275 158612 248276 158676
rect 248340 158612 248341 158676
rect 248275 158611 248341 158612
rect 248646 157997 248706 159430
rect 250118 158677 250178 159430
rect 250854 159221 250914 159430
rect 250851 159220 250917 159221
rect 250851 159156 250852 159220
rect 250916 159156 250917 159220
rect 250851 159155 250917 159156
rect 250115 158676 250181 158677
rect 250115 158612 250116 158676
rect 250180 158612 250181 158676
rect 250115 158611 250181 158612
rect 248643 157996 248709 157997
rect 248643 157932 248644 157996
rect 248708 157932 248709 157996
rect 248643 157931 248709 157932
rect 247723 157044 247789 157045
rect 247723 156980 247724 157044
rect 247788 156980 247789 157044
rect 247723 156979 247789 156980
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6416 245414 29898
rect 244794 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 245414 -6416
rect 244794 -6736 245414 -6652
rect 244794 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 245414 -6736
rect 244794 -7964 245414 -6972
rect 249294 142954 249914 158000
rect 251406 157997 251466 159430
rect 252326 159430 252436 159490
rect 253430 159430 253524 159490
rect 253600 159490 253660 160106
rect 254552 159490 254612 160106
rect 255912 159490 255972 160106
rect 253600 159430 253674 159490
rect 252326 158677 252386 159430
rect 252323 158676 252389 158677
rect 252323 158612 252324 158676
rect 252388 158612 252389 158676
rect 252323 158611 252389 158612
rect 253430 157997 253490 159430
rect 251403 157996 251469 157997
rect 251403 157932 251404 157996
rect 251468 157932 251469 157996
rect 251403 157931 251469 157932
rect 253427 157996 253493 157997
rect 253427 157932 253428 157996
rect 253492 157932 253493 157996
rect 253427 157931 253493 157932
rect 253614 157453 253674 159430
rect 254534 159430 254612 159490
rect 255822 159430 255972 159490
rect 256048 159490 256108 160106
rect 257000 159490 257060 160106
rect 258088 159490 258148 160106
rect 258496 159629 258556 160106
rect 258493 159628 258559 159629
rect 258493 159564 258494 159628
rect 258558 159564 258559 159628
rect 258493 159563 258559 159564
rect 259448 159490 259508 160106
rect 260672 159490 260732 160106
rect 256048 159430 256250 159490
rect 257000 159430 257170 159490
rect 258088 159430 258274 159490
rect 259448 159430 259562 159490
rect 254534 158677 254594 159430
rect 255822 158677 255882 159430
rect 254531 158676 254597 158677
rect 254531 158612 254532 158676
rect 254596 158612 254597 158676
rect 254531 158611 254597 158612
rect 255819 158676 255885 158677
rect 255819 158612 255820 158676
rect 255884 158612 255885 158676
rect 255819 158611 255885 158612
rect 253611 157452 253677 157453
rect 253611 157388 253612 157452
rect 253676 157388 253677 157452
rect 253611 157387 253677 157388
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7376 249914 34398
rect 249294 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 249914 -7376
rect 249294 -7696 249914 -7612
rect 249294 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 249914 -7696
rect 249294 -7964 249914 -7932
rect 253794 147454 254414 158000
rect 256190 157453 256250 159430
rect 257110 158677 257170 159430
rect 258214 158677 258274 159430
rect 259502 158677 259562 159430
rect 260606 159430 260732 159490
rect 261080 159490 261140 160106
rect 261760 159490 261820 160106
rect 262848 159490 262908 160106
rect 261080 159430 261218 159490
rect 257107 158676 257173 158677
rect 257107 158612 257108 158676
rect 257172 158612 257173 158676
rect 257107 158611 257173 158612
rect 258211 158676 258277 158677
rect 258211 158612 258212 158676
rect 258276 158612 258277 158676
rect 258211 158611 258277 158612
rect 259499 158676 259565 158677
rect 259499 158612 259500 158676
rect 259564 158612 259565 158676
rect 259499 158611 259565 158612
rect 256187 157452 256253 157453
rect 256187 157388 256188 157452
rect 256252 157388 256253 157452
rect 256187 157387 256253 157388
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -656 254414 2898
rect 253794 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 254414 -656
rect 253794 -976 254414 -892
rect 253794 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 254414 -976
rect 253794 -7964 254414 -1212
rect 258294 151954 258914 158000
rect 260606 157997 260666 159430
rect 261158 158677 261218 159430
rect 261710 159430 261820 159490
rect 262814 159430 262908 159490
rect 263528 159490 263588 160106
rect 263936 159490 263996 160106
rect 263528 159430 263610 159490
rect 261155 158676 261221 158677
rect 261155 158612 261156 158676
rect 261220 158612 261221 158676
rect 261155 158611 261221 158612
rect 260603 157996 260669 157997
rect 260603 157932 260604 157996
rect 260668 157932 260669 157996
rect 260603 157931 260669 157932
rect 261710 157861 261770 159430
rect 262814 158677 262874 159430
rect 263550 158677 263610 159430
rect 263918 159430 263996 159490
rect 265296 159490 265356 160106
rect 265976 159493 266036 160106
rect 265939 159492 266036 159493
rect 265296 159430 265450 159490
rect 262811 158676 262877 158677
rect 262811 158612 262812 158676
rect 262876 158612 262877 158676
rect 262811 158611 262877 158612
rect 263547 158676 263613 158677
rect 263547 158612 263548 158676
rect 263612 158612 263613 158676
rect 263547 158611 263613 158612
rect 261707 157860 261773 157861
rect 261707 157796 261708 157860
rect 261772 157796 261773 157860
rect 261707 157795 261773 157796
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1616 258914 7398
rect 258294 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 258914 -1616
rect 258294 -1936 258914 -1852
rect 258294 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 258914 -1936
rect 258294 -7964 258914 -2172
rect 262794 156454 263414 158000
rect 263918 157861 263978 159430
rect 263915 157860 263981 157861
rect 263915 157796 263916 157860
rect 263980 157796 263981 157860
rect 263915 157795 263981 157796
rect 265390 157725 265450 159430
rect 265939 159428 265940 159492
rect 266004 159430 266036 159492
rect 266384 159490 266444 160106
rect 267608 159490 267668 160106
rect 266384 159430 266554 159490
rect 266004 159428 266005 159430
rect 265939 159427 266005 159428
rect 266494 157861 266554 159430
rect 267598 159430 267668 159490
rect 268288 159490 268348 160106
rect 268696 159490 268756 160106
rect 269784 159490 269844 160106
rect 271008 159629 271068 160106
rect 271005 159628 271071 159629
rect 271005 159564 271006 159628
rect 271070 159564 271071 159628
rect 271005 159563 271071 159564
rect 271144 159490 271204 160106
rect 272232 159490 272292 160106
rect 273320 159490 273380 160106
rect 268288 159430 268394 159490
rect 268696 159430 268762 159490
rect 269784 159430 269866 159490
rect 267598 158269 267658 159430
rect 267595 158268 267661 158269
rect 267595 158204 267596 158268
rect 267660 158204 267661 158268
rect 267595 158203 267661 158204
rect 266491 157860 266557 157861
rect 266491 157796 266492 157860
rect 266556 157796 266557 157860
rect 266491 157795 266557 157796
rect 265387 157724 265453 157725
rect 265387 157660 265388 157724
rect 265452 157660 265453 157724
rect 265387 157659 265453 157660
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2576 263414 11898
rect 262794 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 263414 -2576
rect 262794 -2896 263414 -2812
rect 262794 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 263414 -2896
rect 262794 -7964 263414 -3132
rect 267294 124954 267914 158000
rect 268334 157861 268394 159430
rect 268702 158677 268762 159430
rect 269806 158677 269866 159430
rect 271094 159430 271204 159490
rect 272198 159430 272292 159490
rect 273302 159430 273380 159490
rect 273592 159490 273652 160106
rect 274408 159490 274468 160106
rect 275768 159629 275828 160106
rect 275765 159628 275831 159629
rect 275765 159564 275766 159628
rect 275830 159564 275831 159628
rect 275765 159563 275831 159564
rect 273592 159430 273730 159490
rect 271094 158677 271154 159430
rect 272198 158677 272258 159430
rect 268699 158676 268765 158677
rect 268699 158612 268700 158676
rect 268764 158612 268765 158676
rect 268699 158611 268765 158612
rect 269803 158676 269869 158677
rect 269803 158612 269804 158676
rect 269868 158612 269869 158676
rect 269803 158611 269869 158612
rect 271091 158676 271157 158677
rect 271091 158612 271092 158676
rect 271156 158612 271157 158676
rect 271091 158611 271157 158612
rect 272195 158676 272261 158677
rect 272195 158612 272196 158676
rect 272260 158612 272261 158676
rect 272195 158611 272261 158612
rect 273302 158405 273362 159430
rect 273299 158404 273365 158405
rect 273299 158340 273300 158404
rect 273364 158340 273365 158404
rect 273299 158339 273365 158340
rect 268331 157860 268397 157861
rect 268331 157796 268332 157860
rect 268396 157796 268397 157860
rect 268331 157795 268397 157796
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3536 267914 16398
rect 267294 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 267914 -3536
rect 267294 -3856 267914 -3772
rect 267294 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 267914 -3856
rect 267294 -7964 267914 -4092
rect 271794 129454 272414 158000
rect 273670 157725 273730 159430
rect 274406 159430 274468 159490
rect 276040 159490 276100 160106
rect 276992 159490 277052 160106
rect 278080 159901 278140 160106
rect 278077 159900 278143 159901
rect 278077 159836 278078 159900
rect 278142 159836 278143 159900
rect 278077 159835 278143 159836
rect 278488 159490 278548 160106
rect 279168 159629 279228 160106
rect 279165 159628 279231 159629
rect 279165 159564 279166 159628
rect 279230 159564 279231 159628
rect 279165 159563 279231 159564
rect 276040 159430 276122 159490
rect 274406 158677 274466 159430
rect 274403 158676 274469 158677
rect 274403 158612 274404 158676
rect 274468 158612 274469 158676
rect 274403 158611 274469 158612
rect 276062 158405 276122 159430
rect 276982 159430 277052 159490
rect 278454 159430 278548 159490
rect 280936 159490 280996 160106
rect 283520 159490 283580 160106
rect 285968 159490 286028 160106
rect 288280 159629 288340 160106
rect 288277 159628 288343 159629
rect 288277 159564 288278 159628
rect 288342 159564 288343 159628
rect 288277 159563 288343 159564
rect 291000 159490 291060 160106
rect 280936 159430 281090 159490
rect 283520 159430 283666 159490
rect 285968 159430 286058 159490
rect 276982 158677 277042 159430
rect 276979 158676 277045 158677
rect 276979 158612 276980 158676
rect 277044 158612 277045 158676
rect 276979 158611 277045 158612
rect 276059 158404 276125 158405
rect 276059 158340 276060 158404
rect 276124 158340 276125 158404
rect 276059 158339 276125 158340
rect 273667 157724 273733 157725
rect 273667 157660 273668 157724
rect 273732 157660 273733 157724
rect 273667 157659 273733 157660
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4496 272414 20898
rect 271794 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 272414 -4496
rect 271794 -4816 272414 -4732
rect 271794 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 272414 -4816
rect 271794 -7964 272414 -5052
rect 276294 133954 276914 158000
rect 278454 157725 278514 159430
rect 281030 158405 281090 159430
rect 281027 158404 281093 158405
rect 281027 158340 281028 158404
rect 281092 158340 281093 158404
rect 281027 158339 281093 158340
rect 278451 157724 278517 157725
rect 278451 157660 278452 157724
rect 278516 157660 278517 157724
rect 278451 157659 278517 157660
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5456 276914 25398
rect 276294 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 276914 -5456
rect 276294 -5776 276914 -5692
rect 276294 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 276914 -5776
rect 276294 -7964 276914 -6012
rect 280794 138454 281414 158000
rect 283606 157589 283666 159430
rect 285998 158405 286058 159430
rect 290966 159430 291060 159490
rect 293448 159490 293508 160106
rect 295896 159629 295956 160106
rect 295893 159628 295959 159629
rect 295893 159564 295894 159628
rect 295958 159564 295959 159628
rect 295893 159563 295959 159564
rect 298480 159490 298540 160106
rect 300928 159765 300988 160106
rect 300925 159764 300991 159765
rect 300925 159700 300926 159764
rect 300990 159700 300991 159764
rect 300925 159699 300991 159700
rect 303512 159490 303572 160106
rect 293448 159430 293602 159490
rect 298480 159430 298570 159490
rect 285995 158404 286061 158405
rect 285995 158340 285996 158404
rect 286060 158340 286061 158404
rect 285995 158339 286061 158340
rect 283603 157588 283669 157589
rect 283603 157524 283604 157588
rect 283668 157524 283669 157588
rect 283603 157523 283669 157524
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6416 281414 29898
rect 280794 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 281414 -6416
rect 280794 -6736 281414 -6652
rect 280794 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 281414 -6736
rect 280794 -7964 281414 -6972
rect 285294 142954 285914 158000
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7376 285914 34398
rect 285294 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 285914 -7376
rect 285294 -7696 285914 -7612
rect 285294 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 285914 -7696
rect 285294 -7964 285914 -7932
rect 289794 147454 290414 158000
rect 290966 157589 291026 159430
rect 293542 158405 293602 159430
rect 298510 158677 298570 159430
rect 303478 159430 303572 159490
rect 305960 159490 306020 160106
rect 308544 159490 308604 160106
rect 310992 159490 311052 160106
rect 313440 159490 313500 160106
rect 315888 159490 315948 160106
rect 305960 159430 306114 159490
rect 308544 159430 308690 159490
rect 310992 159430 311082 159490
rect 303478 158677 303538 159430
rect 306054 158677 306114 159430
rect 308630 158677 308690 159430
rect 298507 158676 298573 158677
rect 298507 158612 298508 158676
rect 298572 158612 298573 158676
rect 298507 158611 298573 158612
rect 303475 158676 303541 158677
rect 303475 158612 303476 158676
rect 303540 158612 303541 158676
rect 303475 158611 303541 158612
rect 306051 158676 306117 158677
rect 306051 158612 306052 158676
rect 306116 158612 306117 158676
rect 306051 158611 306117 158612
rect 308627 158676 308693 158677
rect 308627 158612 308628 158676
rect 308692 158612 308693 158676
rect 308627 158611 308693 158612
rect 293539 158404 293605 158405
rect 293539 158340 293540 158404
rect 293604 158340 293605 158404
rect 293539 158339 293605 158340
rect 311022 158269 311082 159430
rect 313414 159430 313500 159490
rect 315806 159430 315948 159490
rect 318472 159490 318532 160106
rect 320920 159490 320980 160106
rect 323368 159490 323428 160106
rect 325952 159490 326012 160106
rect 318472 159430 318626 159490
rect 320920 159430 321018 159490
rect 313414 158677 313474 159430
rect 315806 158677 315866 159430
rect 318566 158677 318626 159430
rect 320958 158677 321018 159430
rect 323350 159430 323428 159490
rect 325926 159430 326012 159490
rect 323350 158677 323410 159430
rect 325926 158677 325986 159430
rect 313411 158676 313477 158677
rect 313411 158612 313412 158676
rect 313476 158612 313477 158676
rect 313411 158611 313477 158612
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 318563 158676 318629 158677
rect 318563 158612 318564 158676
rect 318628 158612 318629 158676
rect 318563 158611 318629 158612
rect 320955 158676 321021 158677
rect 320955 158612 320956 158676
rect 321020 158612 321021 158676
rect 320955 158611 321021 158612
rect 323347 158676 323413 158677
rect 323347 158612 323348 158676
rect 323412 158612 323413 158676
rect 323347 158611 323413 158612
rect 325923 158676 325989 158677
rect 325923 158612 325924 158676
rect 325988 158612 325989 158676
rect 325923 158611 325989 158612
rect 311019 158268 311085 158269
rect 311019 158204 311020 158268
rect 311084 158204 311085 158268
rect 311019 158203 311085 158204
rect 290963 157588 291029 157589
rect 290963 157524 290964 157588
rect 291028 157524 291029 157588
rect 290963 157523 291029 157524
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -656 290414 2898
rect 289794 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 290414 -656
rect 289794 -976 290414 -892
rect 289794 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 290414 -976
rect 289794 -7964 290414 -1212
rect 294294 151954 294914 158000
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1616 294914 7398
rect 294294 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 294914 -1616
rect 294294 -1936 294914 -1852
rect 294294 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 294914 -1936
rect 294294 -7964 294914 -2172
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2576 299414 11898
rect 298794 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 299414 -2576
rect 298794 -2896 299414 -2812
rect 298794 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 299414 -2896
rect 298794 -7964 299414 -3132
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3536 303914 16398
rect 303294 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 303914 -3536
rect 303294 -3856 303914 -3772
rect 303294 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 303914 -3856
rect 303294 -7964 303914 -4092
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4496 308414 20898
rect 307794 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 308414 -4496
rect 307794 -4816 308414 -4732
rect 307794 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 308414 -4816
rect 307794 -7964 308414 -5052
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5456 312914 25398
rect 312294 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 312914 -5456
rect 312294 -5776 312914 -5692
rect 312294 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 312914 -5776
rect 312294 -7964 312914 -6012
rect 316794 138454 317414 158000
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6416 317414 29898
rect 316794 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 317414 -6416
rect 316794 -6736 317414 -6652
rect 316794 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 317414 -6736
rect 316794 -7964 317414 -6972
rect 321294 142954 321914 158000
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7376 321914 34398
rect 321294 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 321914 -7376
rect 321294 -7696 321914 -7612
rect 321294 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 321914 -7696
rect 321294 -7964 321914 -7932
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -656 326414 2898
rect 325794 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 326414 -656
rect 325794 -976 326414 -892
rect 325794 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 326414 -976
rect 325794 -7964 326414 -1212
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1616 330914 7398
rect 330294 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 330914 -1616
rect 330294 -1936 330914 -1852
rect 330294 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 330914 -1936
rect 330294 -7964 330914 -2172
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2576 335414 11898
rect 334794 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 335414 -2576
rect 334794 -2896 335414 -2812
rect 334794 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 335414 -2896
rect 334794 -7964 335414 -3132
rect 339294 124954 339914 158000
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3536 339914 16398
rect 339294 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 339914 -3536
rect 339294 -3856 339914 -3772
rect 339294 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 339914 -3856
rect 339294 -7964 339914 -4092
rect 343794 129454 344414 158000
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4496 344414 20898
rect 343794 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 344414 -4496
rect 343794 -4816 344414 -4732
rect 343794 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 344414 -4816
rect 343794 -7964 344414 -5052
rect 348294 133954 348914 158000
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5456 348914 25398
rect 348294 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 348914 -5456
rect 348294 -5776 348914 -5692
rect 348294 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 348914 -5776
rect 348294 -7964 348914 -6012
rect 352794 138454 353414 158000
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6416 353414 29898
rect 356838 3365 356898 160107
rect 357574 158949 357634 243475
rect 357571 158948 357637 158949
rect 357571 158884 357572 158948
rect 357636 158884 357637 158948
rect 357571 158883 357637 158884
rect 357294 142954 357914 158000
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 356835 3364 356901 3365
rect 356835 3300 356836 3364
rect 356900 3300 356901 3364
rect 356835 3299 356901 3300
rect 352794 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 353414 -6416
rect 352794 -6736 353414 -6652
rect 352794 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 353414 -6736
rect 352794 -7964 353414 -6972
rect 357294 -7376 357914 34398
rect 358126 3773 358186 247963
rect 358310 6357 358370 250547
rect 358491 244764 358557 244765
rect 358491 244700 358492 244764
rect 358556 244700 358557 244764
rect 358491 244699 358557 244700
rect 358307 6356 358373 6357
rect 358307 6292 358308 6356
rect 358372 6292 358373 6356
rect 358307 6291 358373 6292
rect 358123 3772 358189 3773
rect 358123 3708 358124 3772
rect 358188 3708 358189 3772
rect 358123 3707 358189 3708
rect 358494 3501 358554 244699
rect 358862 3501 358922 250955
rect 359043 250748 359109 250749
rect 359043 250684 359044 250748
rect 359108 250684 359109 250748
rect 359043 250683 359109 250684
rect 359046 6493 359106 250683
rect 359411 245444 359477 245445
rect 359411 245380 359412 245444
rect 359476 245380 359477 245444
rect 359411 245379 359477 245380
rect 359227 245172 359293 245173
rect 359227 245108 359228 245172
rect 359292 245108 359293 245172
rect 359227 245107 359293 245108
rect 359043 6492 359109 6493
rect 359043 6428 359044 6492
rect 359108 6428 359109 6492
rect 359043 6427 359109 6428
rect 358491 3500 358557 3501
rect 358491 3436 358492 3500
rect 358556 3436 358557 3500
rect 358491 3435 358557 3436
rect 358859 3500 358925 3501
rect 358859 3436 358860 3500
rect 358924 3436 358925 3500
rect 358859 3435 358925 3436
rect 359230 3365 359290 245107
rect 359414 4045 359474 245379
rect 359411 4044 359477 4045
rect 359411 3980 359412 4044
rect 359476 3980 359477 4044
rect 359411 3979 359477 3980
rect 360150 3909 360210 302190
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361619 260268 361685 260269
rect 361619 260204 361620 260268
rect 361684 260204 361685 260268
rect 361619 260203 361685 260204
rect 360331 248164 360397 248165
rect 360331 248100 360332 248164
rect 360396 248100 360397 248164
rect 360331 248099 360397 248100
rect 360147 3908 360213 3909
rect 360147 3844 360148 3908
rect 360212 3844 360213 3908
rect 360147 3843 360213 3844
rect 360334 3501 360394 248099
rect 360699 245580 360765 245581
rect 360699 245516 360700 245580
rect 360764 245516 360765 245580
rect 360699 245515 360765 245516
rect 360515 245036 360581 245037
rect 360515 244972 360516 245036
rect 360580 244972 360581 245036
rect 360515 244971 360581 244972
rect 360331 3500 360397 3501
rect 360331 3436 360332 3500
rect 360396 3436 360397 3500
rect 360331 3435 360397 3436
rect 359227 3364 359293 3365
rect 359227 3300 359228 3364
rect 359292 3300 359293 3364
rect 359227 3299 359293 3300
rect 360518 3229 360578 244971
rect 360702 3637 360762 245515
rect 360699 3636 360765 3637
rect 360699 3572 360700 3636
rect 360764 3572 360765 3636
rect 360699 3571 360765 3572
rect 361622 3501 361682 260203
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 364379 254556 364445 254557
rect 364379 254492 364380 254556
rect 364444 254492 364445 254556
rect 364379 254491 364445 254492
rect 362907 250884 362973 250885
rect 362907 250820 362908 250884
rect 362972 250820 362973 250884
rect 362907 250819 362973 250820
rect 362539 245308 362605 245309
rect 362539 245244 362540 245308
rect 362604 245244 362605 245308
rect 362539 245243 362605 245244
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 362542 158949 362602 245243
rect 362539 158948 362605 158949
rect 362539 158884 362540 158948
rect 362604 158884 362605 158948
rect 362539 158883 362605 158884
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361619 3500 361685 3501
rect 361619 3436 361620 3500
rect 361684 3436 361685 3500
rect 361619 3435 361685 3436
rect 361794 3454 362414 38898
rect 362910 3501 362970 250819
rect 363275 247892 363341 247893
rect 363275 247828 363276 247892
rect 363340 247828 363341 247892
rect 363275 247827 363341 247828
rect 363091 247620 363157 247621
rect 363091 247556 363092 247620
rect 363156 247556 363157 247620
rect 363091 247555 363157 247556
rect 360515 3228 360581 3229
rect 360515 3164 360516 3228
rect 360580 3164 360581 3228
rect 360515 3163 360581 3164
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 362907 3500 362973 3501
rect 362907 3436 362908 3500
rect 362972 3436 362973 3500
rect 362907 3435 362973 3436
rect 357294 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 357914 -7376
rect 357294 -7696 357914 -7612
rect 357294 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 357914 -7696
rect 357294 -7964 357914 -7932
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 363094 3093 363154 247555
rect 363278 157453 363338 247827
rect 363459 247756 363525 247757
rect 363459 247692 363460 247756
rect 363524 247692 363525 247756
rect 363459 247691 363525 247692
rect 363462 160173 363522 247691
rect 363459 160172 363525 160173
rect 363459 160108 363460 160172
rect 363524 160108 363525 160172
rect 363459 160107 363525 160108
rect 363275 157452 363341 157453
rect 363275 157388 363276 157452
rect 363340 157388 363341 157452
rect 363275 157387 363341 157388
rect 364382 3501 364442 254491
rect 364563 250476 364629 250477
rect 364563 250412 364564 250476
rect 364628 250412 364629 250476
rect 364563 250411 364629 250412
rect 364566 6629 364626 250411
rect 364934 45661 364994 444619
rect 365118 99517 365178 445707
rect 366294 439954 366914 475398
rect 370794 707068 371414 711900
rect 370794 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 371414 707068
rect 370794 706748 371414 706832
rect 370794 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 371414 706748
rect 370794 696454 371414 706512
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 367875 445908 367941 445909
rect 367875 445844 367876 445908
rect 367940 445844 367941 445908
rect 367875 445843 367941 445844
rect 367691 444412 367757 444413
rect 367691 444348 367692 444412
rect 367756 444348 367757 444412
rect 367691 444347 367757 444348
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 367139 306100 367205 306101
rect 367139 306036 367140 306100
rect 367204 306036 367205 306100
rect 367139 306035 367205 306036
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 365667 260132 365733 260133
rect 365667 260068 365668 260132
rect 365732 260068 365733 260132
rect 365667 260067 365733 260068
rect 365115 99516 365181 99517
rect 365115 99452 365116 99516
rect 365180 99452 365181 99516
rect 365115 99451 365181 99452
rect 364931 45660 364997 45661
rect 364931 45596 364932 45660
rect 364996 45596 364997 45660
rect 364931 45595 364997 45596
rect 364563 6628 364629 6629
rect 364563 6564 364564 6628
rect 364628 6564 364629 6628
rect 364563 6563 364629 6564
rect 365670 3501 365730 260067
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 365851 251836 365917 251837
rect 365851 251772 365852 251836
rect 365916 251772 365917 251836
rect 365851 251771 365917 251772
rect 365854 3637 365914 251771
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 365851 3636 365917 3637
rect 365851 3572 365852 3636
rect 365916 3572 365917 3636
rect 365851 3571 365917 3572
rect 364379 3500 364445 3501
rect 364379 3436 364380 3500
rect 364444 3436 364445 3500
rect 364379 3435 364445 3436
rect 365667 3500 365733 3501
rect 365667 3436 365668 3500
rect 365732 3436 365733 3500
rect 365667 3435 365733 3436
rect 363091 3092 363157 3093
rect 363091 3028 363092 3092
rect 363156 3028 363157 3092
rect 363091 3027 363157 3028
rect 361794 -656 362414 2898
rect 361794 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 362414 -656
rect 361794 -976 362414 -892
rect 361794 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 362414 -976
rect 361794 -7964 362414 -1212
rect 366294 -1616 366914 7398
rect 367142 3501 367202 306035
rect 367323 244900 367389 244901
rect 367323 244836 367324 244900
rect 367388 244836 367389 244900
rect 367323 244835 367389 244836
rect 367326 6221 367386 244835
rect 367694 85645 367754 444347
rect 367878 178125 367938 445843
rect 368979 444548 369045 444549
rect 368979 444484 368980 444548
rect 369044 444484 369045 444548
rect 368979 444483 369045 444484
rect 368611 300116 368677 300117
rect 368611 300052 368612 300116
rect 368676 300052 368677 300116
rect 368611 300051 368677 300052
rect 368427 280804 368493 280805
rect 368427 280740 368428 280804
rect 368492 280740 368493 280804
rect 368427 280739 368493 280740
rect 367875 178124 367941 178125
rect 367875 178060 367876 178124
rect 367940 178060 367941 178124
rect 367875 178059 367941 178060
rect 367691 85644 367757 85645
rect 367691 85580 367692 85644
rect 367756 85580 367757 85644
rect 367691 85579 367757 85580
rect 367323 6220 367389 6221
rect 367323 6156 367324 6220
rect 367388 6156 367389 6220
rect 367323 6155 367389 6156
rect 368430 3501 368490 280739
rect 368614 153781 368674 300051
rect 368611 153780 368677 153781
rect 368611 153716 368612 153780
rect 368676 153716 368677 153780
rect 368611 153715 368677 153716
rect 368982 125629 369042 444483
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 369899 303516 369965 303517
rect 369899 303452 369900 303516
rect 369964 303452 369965 303516
rect 369899 303451 369965 303452
rect 369163 265572 369229 265573
rect 369163 265508 369164 265572
rect 369228 265508 369229 265572
rect 369163 265507 369229 265508
rect 368979 125628 369045 125629
rect 368979 125564 368980 125628
rect 369044 125564 369045 125628
rect 368979 125563 369045 125564
rect 367139 3500 367205 3501
rect 367139 3436 367140 3500
rect 367204 3436 367205 3500
rect 367139 3435 367205 3436
rect 368427 3500 368493 3501
rect 368427 3436 368428 3500
rect 368492 3436 368493 3500
rect 368427 3435 368493 3436
rect 369166 3365 369226 265507
rect 369902 3501 369962 303451
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 369899 3500 369965 3501
rect 369899 3436 369900 3500
rect 369964 3436 369965 3500
rect 369899 3435 369965 3436
rect 369163 3364 369229 3365
rect 369163 3300 369164 3364
rect 369228 3300 369229 3364
rect 369163 3299 369229 3300
rect 366294 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 366914 -1616
rect 366294 -1936 366914 -1852
rect 366294 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 366914 -1936
rect 366294 -7964 366914 -2172
rect 370794 -2576 371414 11898
rect 370794 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 371414 -2576
rect 370794 -2896 371414 -2812
rect 370794 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 371414 -2896
rect 370794 -7964 371414 -3132
rect 375294 708028 375914 711900
rect 375294 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 375914 708028
rect 375294 707708 375914 707792
rect 375294 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 375914 707708
rect 375294 700954 375914 707472
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3536 375914 16398
rect 375294 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 375914 -3536
rect 375294 -3856 375914 -3772
rect 375294 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 375914 -3856
rect 375294 -7964 375914 -4092
rect 379794 708988 380414 711900
rect 379794 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 380414 708988
rect 379794 708668 380414 708752
rect 379794 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 380414 708668
rect 379794 669454 380414 708432
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4496 380414 20898
rect 379794 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 380414 -4496
rect 379794 -4816 380414 -4732
rect 379794 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 380414 -4816
rect 379794 -7964 380414 -5052
rect 384294 709948 384914 711900
rect 384294 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 384914 709948
rect 384294 709628 384914 709712
rect 384294 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 384914 709628
rect 384294 673954 384914 709392
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5456 384914 25398
rect 384294 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 384914 -5456
rect 384294 -5776 384914 -5692
rect 384294 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 384914 -5776
rect 384294 -7964 384914 -6012
rect 388794 710908 389414 711900
rect 388794 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 389414 710908
rect 388794 710588 389414 710672
rect 388794 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 389414 710588
rect 388794 678454 389414 710352
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6416 389414 29898
rect 388794 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 389414 -6416
rect 388794 -6736 389414 -6652
rect 388794 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 389414 -6736
rect 388794 -7964 389414 -6972
rect 393294 711868 393914 711900
rect 393294 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 393914 711868
rect 393294 711548 393914 711632
rect 393294 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 393914 711548
rect 393294 682954 393914 711312
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7376 393914 34398
rect 393294 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 393914 -7376
rect 393294 -7696 393914 -7612
rect 393294 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 393914 -7696
rect 393294 -7964 393914 -7932
rect 397794 705148 398414 711900
rect 397794 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 398414 705148
rect 397794 704828 398414 704912
rect 397794 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 398414 704828
rect 397794 687454 398414 704592
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -656 398414 2898
rect 397794 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 398414 -656
rect 397794 -976 398414 -892
rect 397794 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 398414 -976
rect 397794 -7964 398414 -1212
rect 402294 706108 402914 711900
rect 402294 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 402914 706108
rect 402294 705788 402914 705872
rect 402294 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 402914 705788
rect 402294 691954 402914 705552
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1616 402914 7398
rect 402294 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 402914 -1616
rect 402294 -1936 402914 -1852
rect 402294 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 402914 -1936
rect 402294 -7964 402914 -2172
rect 406794 707068 407414 711900
rect 406794 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 407414 707068
rect 406794 706748 407414 706832
rect 406794 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 407414 706748
rect 406794 696454 407414 706512
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2576 407414 11898
rect 406794 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 407414 -2576
rect 406794 -2896 407414 -2812
rect 406794 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 407414 -2896
rect 406794 -7964 407414 -3132
rect 411294 708028 411914 711900
rect 411294 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 411914 708028
rect 411294 707708 411914 707792
rect 411294 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 411914 707708
rect 411294 700954 411914 707472
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3536 411914 16398
rect 411294 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 411914 -3536
rect 411294 -3856 411914 -3772
rect 411294 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 411914 -3856
rect 411294 -7964 411914 -4092
rect 415794 708988 416414 711900
rect 415794 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 416414 708988
rect 415794 708668 416414 708752
rect 415794 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 416414 708668
rect 415794 669454 416414 708432
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4496 416414 20898
rect 415794 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 416414 -4496
rect 415794 -4816 416414 -4732
rect 415794 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 416414 -4816
rect 415794 -7964 416414 -5052
rect 420294 709948 420914 711900
rect 420294 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 420914 709948
rect 420294 709628 420914 709712
rect 420294 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 420914 709628
rect 420294 673954 420914 709392
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5456 420914 25398
rect 420294 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 420914 -5456
rect 420294 -5776 420914 -5692
rect 420294 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 420914 -5776
rect 420294 -7964 420914 -6012
rect 424794 710908 425414 711900
rect 424794 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 425414 710908
rect 424794 710588 425414 710672
rect 424794 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 425414 710588
rect 424794 678454 425414 710352
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6416 425414 29898
rect 424794 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 425414 -6416
rect 424794 -6736 425414 -6652
rect 424794 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 425414 -6736
rect 424794 -7964 425414 -6972
rect 429294 711868 429914 711900
rect 429294 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 429914 711868
rect 429294 711548 429914 711632
rect 429294 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 429914 711548
rect 429294 682954 429914 711312
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7376 429914 34398
rect 429294 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 429914 -7376
rect 429294 -7696 429914 -7612
rect 429294 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 429914 -7696
rect 429294 -7964 429914 -7932
rect 433794 705148 434414 711900
rect 433794 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 434414 705148
rect 433794 704828 434414 704912
rect 433794 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 434414 704828
rect 433794 687454 434414 704592
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -656 434414 2898
rect 433794 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 434414 -656
rect 433794 -976 434414 -892
rect 433794 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 434414 -976
rect 433794 -7964 434414 -1212
rect 438294 706108 438914 711900
rect 438294 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 438914 706108
rect 438294 705788 438914 705872
rect 438294 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 438914 705788
rect 438294 691954 438914 705552
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1616 438914 7398
rect 438294 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 438914 -1616
rect 438294 -1936 438914 -1852
rect 438294 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 438914 -1936
rect 438294 -7964 438914 -2172
rect 442794 707068 443414 711900
rect 442794 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 443414 707068
rect 442794 706748 443414 706832
rect 442794 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 443414 706748
rect 442794 696454 443414 706512
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2576 443414 11898
rect 442794 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 443414 -2576
rect 442794 -2896 443414 -2812
rect 442794 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 443414 -2896
rect 442794 -7964 443414 -3132
rect 447294 708028 447914 711900
rect 447294 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 447914 708028
rect 447294 707708 447914 707792
rect 447294 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 447914 707708
rect 447294 700954 447914 707472
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3536 447914 16398
rect 447294 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 447914 -3536
rect 447294 -3856 447914 -3772
rect 447294 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 447914 -3856
rect 447294 -7964 447914 -4092
rect 451794 708988 452414 711900
rect 451794 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 452414 708988
rect 451794 708668 452414 708752
rect 451794 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 452414 708668
rect 451794 669454 452414 708432
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4496 452414 20898
rect 451794 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 452414 -4496
rect 451794 -4816 452414 -4732
rect 451794 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 452414 -4816
rect 451794 -7964 452414 -5052
rect 456294 709948 456914 711900
rect 456294 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 456914 709948
rect 456294 709628 456914 709712
rect 456294 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 456914 709628
rect 456294 673954 456914 709392
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5456 456914 25398
rect 456294 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 456914 -5456
rect 456294 -5776 456914 -5692
rect 456294 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 456914 -5776
rect 456294 -7964 456914 -6012
rect 460794 710908 461414 711900
rect 460794 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 461414 710908
rect 460794 710588 461414 710672
rect 460794 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 461414 710588
rect 460794 678454 461414 710352
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6416 461414 29898
rect 460794 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 461414 -6416
rect 460794 -6736 461414 -6652
rect 460794 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 461414 -6736
rect 460794 -7964 461414 -6972
rect 465294 711868 465914 711900
rect 465294 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 465914 711868
rect 465294 711548 465914 711632
rect 465294 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 465914 711548
rect 465294 682954 465914 711312
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7376 465914 34398
rect 465294 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 465914 -7376
rect 465294 -7696 465914 -7612
rect 465294 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 465914 -7696
rect 465294 -7964 465914 -7932
rect 469794 705148 470414 711900
rect 469794 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 470414 705148
rect 469794 704828 470414 704912
rect 469794 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 470414 704828
rect 469794 687454 470414 704592
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -656 470414 2898
rect 469794 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 470414 -656
rect 469794 -976 470414 -892
rect 469794 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 470414 -976
rect 469794 -7964 470414 -1212
rect 474294 706108 474914 711900
rect 474294 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 474914 706108
rect 474294 705788 474914 705872
rect 474294 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 474914 705788
rect 474294 691954 474914 705552
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1616 474914 7398
rect 474294 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 474914 -1616
rect 474294 -1936 474914 -1852
rect 474294 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 474914 -1936
rect 474294 -7964 474914 -2172
rect 478794 707068 479414 711900
rect 478794 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 479414 707068
rect 478794 706748 479414 706832
rect 478794 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 479414 706748
rect 478794 696454 479414 706512
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2576 479414 11898
rect 478794 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 479414 -2576
rect 478794 -2896 479414 -2812
rect 478794 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 479414 -2896
rect 478794 -7964 479414 -3132
rect 483294 708028 483914 711900
rect 483294 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 483914 708028
rect 483294 707708 483914 707792
rect 483294 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 483914 707708
rect 483294 700954 483914 707472
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3536 483914 16398
rect 483294 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 483914 -3536
rect 483294 -3856 483914 -3772
rect 483294 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 483914 -3856
rect 483294 -7964 483914 -4092
rect 487794 708988 488414 711900
rect 487794 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 488414 708988
rect 487794 708668 488414 708752
rect 487794 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 488414 708668
rect 487794 669454 488414 708432
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4496 488414 20898
rect 487794 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 488414 -4496
rect 487794 -4816 488414 -4732
rect 487794 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 488414 -4816
rect 487794 -7964 488414 -5052
rect 492294 709948 492914 711900
rect 492294 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 492914 709948
rect 492294 709628 492914 709712
rect 492294 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 492914 709628
rect 492294 673954 492914 709392
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5456 492914 25398
rect 492294 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 492914 -5456
rect 492294 -5776 492914 -5692
rect 492294 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 492914 -5776
rect 492294 -7964 492914 -6012
rect 496794 710908 497414 711900
rect 496794 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 497414 710908
rect 496794 710588 497414 710672
rect 496794 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 497414 710588
rect 496794 678454 497414 710352
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6416 497414 29898
rect 496794 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 497414 -6416
rect 496794 -6736 497414 -6652
rect 496794 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 497414 -6736
rect 496794 -7964 497414 -6972
rect 501294 711868 501914 711900
rect 501294 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 501914 711868
rect 501294 711548 501914 711632
rect 501294 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 501914 711548
rect 501294 682954 501914 711312
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7376 501914 34398
rect 501294 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 501914 -7376
rect 501294 -7696 501914 -7612
rect 501294 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 501914 -7696
rect 501294 -7964 501914 -7932
rect 505794 705148 506414 711900
rect 505794 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 506414 705148
rect 505794 704828 506414 704912
rect 505794 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 506414 704828
rect 505794 687454 506414 704592
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -656 506414 2898
rect 505794 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 506414 -656
rect 505794 -976 506414 -892
rect 505794 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 506414 -976
rect 505794 -7964 506414 -1212
rect 510294 706108 510914 711900
rect 510294 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 510914 706108
rect 510294 705788 510914 705872
rect 510294 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 510914 705788
rect 510294 691954 510914 705552
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1616 510914 7398
rect 510294 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 510914 -1616
rect 510294 -1936 510914 -1852
rect 510294 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 510914 -1936
rect 510294 -7964 510914 -2172
rect 514794 707068 515414 711900
rect 514794 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 515414 707068
rect 514794 706748 515414 706832
rect 514794 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 515414 706748
rect 514794 696454 515414 706512
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2576 515414 11898
rect 514794 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 515414 -2576
rect 514794 -2896 515414 -2812
rect 514794 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 515414 -2896
rect 514794 -7964 515414 -3132
rect 519294 708028 519914 711900
rect 519294 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 519914 708028
rect 519294 707708 519914 707792
rect 519294 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 519914 707708
rect 519294 700954 519914 707472
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3536 519914 16398
rect 519294 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 519914 -3536
rect 519294 -3856 519914 -3772
rect 519294 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 519914 -3856
rect 519294 -7964 519914 -4092
rect 523794 708988 524414 711900
rect 523794 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 524414 708988
rect 523794 708668 524414 708752
rect 523794 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 524414 708668
rect 523794 669454 524414 708432
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4496 524414 20898
rect 523794 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 524414 -4496
rect 523794 -4816 524414 -4732
rect 523794 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 524414 -4816
rect 523794 -7964 524414 -5052
rect 528294 709948 528914 711900
rect 528294 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 528914 709948
rect 528294 709628 528914 709712
rect 528294 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 528914 709628
rect 528294 673954 528914 709392
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5456 528914 25398
rect 528294 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 528914 -5456
rect 528294 -5776 528914 -5692
rect 528294 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 528914 -5776
rect 528294 -7964 528914 -6012
rect 532794 710908 533414 711900
rect 532794 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 533414 710908
rect 532794 710588 533414 710672
rect 532794 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 533414 710588
rect 532794 678454 533414 710352
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6416 533414 29898
rect 532794 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 533414 -6416
rect 532794 -6736 533414 -6652
rect 532794 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 533414 -6736
rect 532794 -7964 533414 -6972
rect 537294 711868 537914 711900
rect 537294 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 537914 711868
rect 537294 711548 537914 711632
rect 537294 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 537914 711548
rect 537294 682954 537914 711312
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7376 537914 34398
rect 537294 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 537914 -7376
rect 537294 -7696 537914 -7612
rect 537294 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 537914 -7696
rect 537294 -7964 537914 -7932
rect 541794 705148 542414 711900
rect 541794 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 542414 705148
rect 541794 704828 542414 704912
rect 541794 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 542414 704828
rect 541794 687454 542414 704592
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -656 542414 2898
rect 541794 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 542414 -656
rect 541794 -976 542414 -892
rect 541794 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 542414 -976
rect 541794 -7964 542414 -1212
rect 546294 706108 546914 711900
rect 546294 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 546914 706108
rect 546294 705788 546914 705872
rect 546294 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 546914 705788
rect 546294 691954 546914 705552
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1616 546914 7398
rect 546294 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 546914 -1616
rect 546294 -1936 546914 -1852
rect 546294 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 546914 -1936
rect 546294 -7964 546914 -2172
rect 550794 707068 551414 711900
rect 550794 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 551414 707068
rect 550794 706748 551414 706832
rect 550794 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 551414 706748
rect 550794 696454 551414 706512
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2576 551414 11898
rect 550794 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 551414 -2576
rect 550794 -2896 551414 -2812
rect 550794 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 551414 -2896
rect 550794 -7964 551414 -3132
rect 555294 708028 555914 711900
rect 555294 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 555914 708028
rect 555294 707708 555914 707792
rect 555294 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 555914 707708
rect 555294 700954 555914 707472
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3536 555914 16398
rect 555294 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 555914 -3536
rect 555294 -3856 555914 -3772
rect 555294 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 555914 -3856
rect 555294 -7964 555914 -4092
rect 559794 708988 560414 711900
rect 559794 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 560414 708988
rect 559794 708668 560414 708752
rect 559794 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 560414 708668
rect 559794 669454 560414 708432
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4496 560414 20898
rect 559794 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 560414 -4496
rect 559794 -4816 560414 -4732
rect 559794 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 560414 -4816
rect 559794 -7964 560414 -5052
rect 564294 709948 564914 711900
rect 564294 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 564914 709948
rect 564294 709628 564914 709712
rect 564294 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 564914 709628
rect 564294 673954 564914 709392
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5456 564914 25398
rect 564294 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 564914 -5456
rect 564294 -5776 564914 -5692
rect 564294 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 564914 -5776
rect 564294 -7964 564914 -6012
rect 568794 710908 569414 711900
rect 568794 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 569414 710908
rect 568794 710588 569414 710672
rect 568794 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 569414 710588
rect 568794 678454 569414 710352
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6416 569414 29898
rect 568794 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 569414 -6416
rect 568794 -6736 569414 -6652
rect 568794 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 569414 -6736
rect 568794 -7964 569414 -6972
rect 573294 711868 573914 711900
rect 573294 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 573914 711868
rect 573294 711548 573914 711632
rect 573294 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 573914 711548
rect 573294 682954 573914 711312
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7376 573914 34398
rect 573294 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 573914 -7376
rect 573294 -7696 573914 -7612
rect 573294 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 573914 -7696
rect 573294 -7964 573914 -7932
rect 577794 705148 578414 711900
rect 577794 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 578414 705148
rect 577794 704828 578414 704912
rect 577794 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 578414 704828
rect 577794 687454 578414 704592
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -656 578414 2898
rect 577794 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 578414 -656
rect 577794 -976 578414 -892
rect 577794 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 578414 -976
rect 577794 -7964 578414 -1212
rect 582294 706108 582914 711900
rect 592340 711868 592960 711900
rect 592340 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect 592340 711548 592960 711632
rect 592340 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect 591380 710908 592000 710940
rect 591380 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect 591380 710588 592000 710672
rect 591380 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect 590420 709948 591040 709980
rect 590420 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect 590420 709628 591040 709712
rect 590420 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect 589460 708988 590080 709020
rect 589460 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect 589460 708668 590080 708752
rect 589460 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect 588500 708028 589120 708060
rect 588500 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect 588500 707708 589120 707792
rect 588500 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect 587540 707068 588160 707100
rect 587540 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect 587540 706748 588160 706832
rect 587540 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect 582294 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 582914 706108
rect 582294 705788 582914 705872
rect 582294 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 582914 705788
rect 582294 691954 582914 705552
rect 586580 706108 587200 706140
rect 586580 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect 586580 705788 587200 705872
rect 586580 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1616 582914 7398
rect 585620 705148 586240 705180
rect 585620 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect 585620 704828 586240 704912
rect 585620 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect 585620 687454 586240 704592
rect 585620 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 586240 687454
rect 585620 687134 586240 687218
rect 585620 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 586240 687134
rect 585620 651454 586240 686898
rect 585620 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 586240 651454
rect 585620 651134 586240 651218
rect 585620 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 586240 651134
rect 585620 615454 586240 650898
rect 585620 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 586240 615454
rect 585620 615134 586240 615218
rect 585620 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 586240 615134
rect 585620 579454 586240 614898
rect 585620 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 586240 579454
rect 585620 579134 586240 579218
rect 585620 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 586240 579134
rect 585620 543454 586240 578898
rect 585620 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 586240 543454
rect 585620 543134 586240 543218
rect 585620 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 586240 543134
rect 585620 507454 586240 542898
rect 585620 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 586240 507454
rect 585620 507134 586240 507218
rect 585620 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 586240 507134
rect 585620 471454 586240 506898
rect 585620 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 586240 471454
rect 585620 471134 586240 471218
rect 585620 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 586240 471134
rect 585620 435454 586240 470898
rect 585620 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 586240 435454
rect 585620 435134 586240 435218
rect 585620 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 586240 435134
rect 585620 399454 586240 434898
rect 585620 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 586240 399454
rect 585620 399134 586240 399218
rect 585620 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 586240 399134
rect 585620 363454 586240 398898
rect 585620 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 586240 363454
rect 585620 363134 586240 363218
rect 585620 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 586240 363134
rect 585620 327454 586240 362898
rect 585620 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 586240 327454
rect 585620 327134 586240 327218
rect 585620 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 586240 327134
rect 585620 291454 586240 326898
rect 585620 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 586240 291454
rect 585620 291134 586240 291218
rect 585620 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 586240 291134
rect 585620 255454 586240 290898
rect 585620 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 586240 255454
rect 585620 255134 586240 255218
rect 585620 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 586240 255134
rect 585620 219454 586240 254898
rect 585620 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 586240 219454
rect 585620 219134 586240 219218
rect 585620 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 586240 219134
rect 585620 183454 586240 218898
rect 585620 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 586240 183454
rect 585620 183134 586240 183218
rect 585620 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 586240 183134
rect 585620 147454 586240 182898
rect 585620 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 586240 147454
rect 585620 147134 586240 147218
rect 585620 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 586240 147134
rect 585620 111454 586240 146898
rect 585620 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 586240 111454
rect 585620 111134 586240 111218
rect 585620 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 586240 111134
rect 585620 75454 586240 110898
rect 585620 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 586240 75454
rect 585620 75134 586240 75218
rect 585620 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 586240 75134
rect 585620 39454 586240 74898
rect 585620 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 586240 39454
rect 585620 39134 586240 39218
rect 585620 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 586240 39134
rect 585620 3454 586240 38898
rect 585620 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 586240 3454
rect 585620 3134 586240 3218
rect 585620 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 586240 3134
rect 585620 -656 586240 2898
rect 585620 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect 585620 -976 586240 -892
rect 585620 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect 585620 -1244 586240 -1212
rect 586580 691954 587200 705552
rect 586580 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 587200 691954
rect 586580 691634 587200 691718
rect 586580 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 587200 691634
rect 586580 655954 587200 691398
rect 586580 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 587200 655954
rect 586580 655634 587200 655718
rect 586580 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 587200 655634
rect 586580 619954 587200 655398
rect 586580 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 587200 619954
rect 586580 619634 587200 619718
rect 586580 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 587200 619634
rect 586580 583954 587200 619398
rect 586580 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 587200 583954
rect 586580 583634 587200 583718
rect 586580 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 587200 583634
rect 586580 547954 587200 583398
rect 586580 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 587200 547954
rect 586580 547634 587200 547718
rect 586580 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 587200 547634
rect 586580 511954 587200 547398
rect 586580 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 587200 511954
rect 586580 511634 587200 511718
rect 586580 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 587200 511634
rect 586580 475954 587200 511398
rect 586580 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 587200 475954
rect 586580 475634 587200 475718
rect 586580 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 587200 475634
rect 586580 439954 587200 475398
rect 586580 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 587200 439954
rect 586580 439634 587200 439718
rect 586580 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 587200 439634
rect 586580 403954 587200 439398
rect 586580 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 587200 403954
rect 586580 403634 587200 403718
rect 586580 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 587200 403634
rect 586580 367954 587200 403398
rect 586580 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 587200 367954
rect 586580 367634 587200 367718
rect 586580 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 587200 367634
rect 586580 331954 587200 367398
rect 586580 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 587200 331954
rect 586580 331634 587200 331718
rect 586580 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 587200 331634
rect 586580 295954 587200 331398
rect 586580 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 587200 295954
rect 586580 295634 587200 295718
rect 586580 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 587200 295634
rect 586580 259954 587200 295398
rect 586580 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 587200 259954
rect 586580 259634 587200 259718
rect 586580 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 587200 259634
rect 586580 223954 587200 259398
rect 586580 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 587200 223954
rect 586580 223634 587200 223718
rect 586580 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 587200 223634
rect 586580 187954 587200 223398
rect 586580 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 587200 187954
rect 586580 187634 587200 187718
rect 586580 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 587200 187634
rect 586580 151954 587200 187398
rect 586580 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 587200 151954
rect 586580 151634 587200 151718
rect 586580 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 587200 151634
rect 586580 115954 587200 151398
rect 586580 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 587200 115954
rect 586580 115634 587200 115718
rect 586580 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 587200 115634
rect 586580 79954 587200 115398
rect 586580 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 587200 79954
rect 586580 79634 587200 79718
rect 586580 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 587200 79634
rect 586580 43954 587200 79398
rect 586580 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 587200 43954
rect 586580 43634 587200 43718
rect 586580 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 587200 43634
rect 586580 7954 587200 43398
rect 586580 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 587200 7954
rect 586580 7634 587200 7718
rect 586580 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 587200 7634
rect 582294 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 582914 -1616
rect 582294 -1936 582914 -1852
rect 582294 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 582914 -1936
rect 582294 -7964 582914 -2172
rect 586580 -1616 587200 7398
rect 586580 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect 586580 -1936 587200 -1852
rect 586580 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect 586580 -2204 587200 -2172
rect 587540 696454 588160 706512
rect 587540 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 588160 696454
rect 587540 696134 588160 696218
rect 587540 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 588160 696134
rect 587540 660454 588160 695898
rect 587540 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 588160 660454
rect 587540 660134 588160 660218
rect 587540 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 588160 660134
rect 587540 624454 588160 659898
rect 587540 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 588160 624454
rect 587540 624134 588160 624218
rect 587540 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 588160 624134
rect 587540 588454 588160 623898
rect 587540 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 588160 588454
rect 587540 588134 588160 588218
rect 587540 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 588160 588134
rect 587540 552454 588160 587898
rect 587540 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 588160 552454
rect 587540 552134 588160 552218
rect 587540 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 588160 552134
rect 587540 516454 588160 551898
rect 587540 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 588160 516454
rect 587540 516134 588160 516218
rect 587540 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 588160 516134
rect 587540 480454 588160 515898
rect 587540 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 588160 480454
rect 587540 480134 588160 480218
rect 587540 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 588160 480134
rect 587540 444454 588160 479898
rect 587540 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 588160 444454
rect 587540 444134 588160 444218
rect 587540 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 588160 444134
rect 587540 408454 588160 443898
rect 587540 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 588160 408454
rect 587540 408134 588160 408218
rect 587540 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 588160 408134
rect 587540 372454 588160 407898
rect 587540 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 588160 372454
rect 587540 372134 588160 372218
rect 587540 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 588160 372134
rect 587540 336454 588160 371898
rect 587540 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 588160 336454
rect 587540 336134 588160 336218
rect 587540 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 588160 336134
rect 587540 300454 588160 335898
rect 587540 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 588160 300454
rect 587540 300134 588160 300218
rect 587540 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 588160 300134
rect 587540 264454 588160 299898
rect 587540 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 588160 264454
rect 587540 264134 588160 264218
rect 587540 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 588160 264134
rect 587540 228454 588160 263898
rect 587540 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 588160 228454
rect 587540 228134 588160 228218
rect 587540 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 588160 228134
rect 587540 192454 588160 227898
rect 587540 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 588160 192454
rect 587540 192134 588160 192218
rect 587540 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 588160 192134
rect 587540 156454 588160 191898
rect 587540 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 588160 156454
rect 587540 156134 588160 156218
rect 587540 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 588160 156134
rect 587540 120454 588160 155898
rect 587540 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 588160 120454
rect 587540 120134 588160 120218
rect 587540 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 588160 120134
rect 587540 84454 588160 119898
rect 587540 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 588160 84454
rect 587540 84134 588160 84218
rect 587540 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 588160 84134
rect 587540 48454 588160 83898
rect 587540 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 588160 48454
rect 587540 48134 588160 48218
rect 587540 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 588160 48134
rect 587540 12454 588160 47898
rect 587540 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 588160 12454
rect 587540 12134 588160 12218
rect 587540 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 588160 12134
rect 587540 -2576 588160 11898
rect 587540 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect 587540 -2896 588160 -2812
rect 587540 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect 587540 -3164 588160 -3132
rect 588500 700954 589120 707472
rect 588500 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 589120 700954
rect 588500 700634 589120 700718
rect 588500 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 589120 700634
rect 588500 664954 589120 700398
rect 588500 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 589120 664954
rect 588500 664634 589120 664718
rect 588500 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 589120 664634
rect 588500 628954 589120 664398
rect 588500 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 589120 628954
rect 588500 628634 589120 628718
rect 588500 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 589120 628634
rect 588500 592954 589120 628398
rect 588500 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 589120 592954
rect 588500 592634 589120 592718
rect 588500 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 589120 592634
rect 588500 556954 589120 592398
rect 588500 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 589120 556954
rect 588500 556634 589120 556718
rect 588500 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 589120 556634
rect 588500 520954 589120 556398
rect 588500 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 589120 520954
rect 588500 520634 589120 520718
rect 588500 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 589120 520634
rect 588500 484954 589120 520398
rect 588500 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 589120 484954
rect 588500 484634 589120 484718
rect 588500 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 589120 484634
rect 588500 448954 589120 484398
rect 588500 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 589120 448954
rect 588500 448634 589120 448718
rect 588500 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 589120 448634
rect 588500 412954 589120 448398
rect 588500 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 589120 412954
rect 588500 412634 589120 412718
rect 588500 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 589120 412634
rect 588500 376954 589120 412398
rect 588500 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 589120 376954
rect 588500 376634 589120 376718
rect 588500 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 589120 376634
rect 588500 340954 589120 376398
rect 588500 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 589120 340954
rect 588500 340634 589120 340718
rect 588500 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 589120 340634
rect 588500 304954 589120 340398
rect 588500 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 589120 304954
rect 588500 304634 589120 304718
rect 588500 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 589120 304634
rect 588500 268954 589120 304398
rect 588500 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 589120 268954
rect 588500 268634 589120 268718
rect 588500 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 589120 268634
rect 588500 232954 589120 268398
rect 588500 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 589120 232954
rect 588500 232634 589120 232718
rect 588500 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 589120 232634
rect 588500 196954 589120 232398
rect 588500 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 589120 196954
rect 588500 196634 589120 196718
rect 588500 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 589120 196634
rect 588500 160954 589120 196398
rect 588500 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 589120 160954
rect 588500 160634 589120 160718
rect 588500 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 589120 160634
rect 588500 124954 589120 160398
rect 588500 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 589120 124954
rect 588500 124634 589120 124718
rect 588500 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 589120 124634
rect 588500 88954 589120 124398
rect 588500 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 589120 88954
rect 588500 88634 589120 88718
rect 588500 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 589120 88634
rect 588500 52954 589120 88398
rect 588500 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 589120 52954
rect 588500 52634 589120 52718
rect 588500 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 589120 52634
rect 588500 16954 589120 52398
rect 588500 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 589120 16954
rect 588500 16634 589120 16718
rect 588500 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 589120 16634
rect 588500 -3536 589120 16398
rect 588500 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect 588500 -3856 589120 -3772
rect 588500 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect 588500 -4124 589120 -4092
rect 589460 669454 590080 708432
rect 589460 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 590080 669454
rect 589460 669134 590080 669218
rect 589460 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 590080 669134
rect 589460 633454 590080 668898
rect 589460 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 590080 633454
rect 589460 633134 590080 633218
rect 589460 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 590080 633134
rect 589460 597454 590080 632898
rect 589460 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 590080 597454
rect 589460 597134 590080 597218
rect 589460 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 590080 597134
rect 589460 561454 590080 596898
rect 589460 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 590080 561454
rect 589460 561134 590080 561218
rect 589460 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 590080 561134
rect 589460 525454 590080 560898
rect 589460 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 590080 525454
rect 589460 525134 590080 525218
rect 589460 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 590080 525134
rect 589460 489454 590080 524898
rect 589460 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 590080 489454
rect 589460 489134 590080 489218
rect 589460 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 590080 489134
rect 589460 453454 590080 488898
rect 589460 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 590080 453454
rect 589460 453134 590080 453218
rect 589460 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 590080 453134
rect 589460 417454 590080 452898
rect 589460 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 590080 417454
rect 589460 417134 590080 417218
rect 589460 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 590080 417134
rect 589460 381454 590080 416898
rect 589460 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 590080 381454
rect 589460 381134 590080 381218
rect 589460 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 590080 381134
rect 589460 345454 590080 380898
rect 589460 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 590080 345454
rect 589460 345134 590080 345218
rect 589460 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 590080 345134
rect 589460 309454 590080 344898
rect 589460 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 590080 309454
rect 589460 309134 590080 309218
rect 589460 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 590080 309134
rect 589460 273454 590080 308898
rect 589460 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 590080 273454
rect 589460 273134 590080 273218
rect 589460 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 590080 273134
rect 589460 237454 590080 272898
rect 589460 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 590080 237454
rect 589460 237134 590080 237218
rect 589460 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 590080 237134
rect 589460 201454 590080 236898
rect 589460 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 590080 201454
rect 589460 201134 590080 201218
rect 589460 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 590080 201134
rect 589460 165454 590080 200898
rect 589460 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 590080 165454
rect 589460 165134 590080 165218
rect 589460 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 590080 165134
rect 589460 129454 590080 164898
rect 589460 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 590080 129454
rect 589460 129134 590080 129218
rect 589460 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 590080 129134
rect 589460 93454 590080 128898
rect 589460 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 590080 93454
rect 589460 93134 590080 93218
rect 589460 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 590080 93134
rect 589460 57454 590080 92898
rect 589460 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 590080 57454
rect 589460 57134 590080 57218
rect 589460 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 590080 57134
rect 589460 21454 590080 56898
rect 589460 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 590080 21454
rect 589460 21134 590080 21218
rect 589460 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 590080 21134
rect 589460 -4496 590080 20898
rect 589460 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect 589460 -4816 590080 -4732
rect 589460 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect 589460 -5084 590080 -5052
rect 590420 673954 591040 709392
rect 590420 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 591040 673954
rect 590420 673634 591040 673718
rect 590420 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 591040 673634
rect 590420 637954 591040 673398
rect 590420 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 591040 637954
rect 590420 637634 591040 637718
rect 590420 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 591040 637634
rect 590420 601954 591040 637398
rect 590420 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 591040 601954
rect 590420 601634 591040 601718
rect 590420 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 591040 601634
rect 590420 565954 591040 601398
rect 590420 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 591040 565954
rect 590420 565634 591040 565718
rect 590420 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 591040 565634
rect 590420 529954 591040 565398
rect 590420 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 591040 529954
rect 590420 529634 591040 529718
rect 590420 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 591040 529634
rect 590420 493954 591040 529398
rect 590420 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 591040 493954
rect 590420 493634 591040 493718
rect 590420 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 591040 493634
rect 590420 457954 591040 493398
rect 590420 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 591040 457954
rect 590420 457634 591040 457718
rect 590420 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 591040 457634
rect 590420 421954 591040 457398
rect 590420 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 591040 421954
rect 590420 421634 591040 421718
rect 590420 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 591040 421634
rect 590420 385954 591040 421398
rect 590420 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 591040 385954
rect 590420 385634 591040 385718
rect 590420 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 591040 385634
rect 590420 349954 591040 385398
rect 590420 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 591040 349954
rect 590420 349634 591040 349718
rect 590420 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 591040 349634
rect 590420 313954 591040 349398
rect 590420 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 591040 313954
rect 590420 313634 591040 313718
rect 590420 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 591040 313634
rect 590420 277954 591040 313398
rect 590420 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 591040 277954
rect 590420 277634 591040 277718
rect 590420 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 591040 277634
rect 590420 241954 591040 277398
rect 590420 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 591040 241954
rect 590420 241634 591040 241718
rect 590420 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 591040 241634
rect 590420 205954 591040 241398
rect 590420 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 591040 205954
rect 590420 205634 591040 205718
rect 590420 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 591040 205634
rect 590420 169954 591040 205398
rect 590420 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 591040 169954
rect 590420 169634 591040 169718
rect 590420 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 591040 169634
rect 590420 133954 591040 169398
rect 590420 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 591040 133954
rect 590420 133634 591040 133718
rect 590420 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 591040 133634
rect 590420 97954 591040 133398
rect 590420 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 591040 97954
rect 590420 97634 591040 97718
rect 590420 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 591040 97634
rect 590420 61954 591040 97398
rect 590420 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 591040 61954
rect 590420 61634 591040 61718
rect 590420 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 591040 61634
rect 590420 25954 591040 61398
rect 590420 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 591040 25954
rect 590420 25634 591040 25718
rect 590420 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 591040 25634
rect 590420 -5456 591040 25398
rect 590420 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect 590420 -5776 591040 -5692
rect 590420 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect 590420 -6044 591040 -6012
rect 591380 678454 592000 710352
rect 591380 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592000 678454
rect 591380 678134 592000 678218
rect 591380 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592000 678134
rect 591380 642454 592000 677898
rect 591380 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592000 642454
rect 591380 642134 592000 642218
rect 591380 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592000 642134
rect 591380 606454 592000 641898
rect 591380 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592000 606454
rect 591380 606134 592000 606218
rect 591380 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592000 606134
rect 591380 570454 592000 605898
rect 591380 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592000 570454
rect 591380 570134 592000 570218
rect 591380 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592000 570134
rect 591380 534454 592000 569898
rect 591380 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592000 534454
rect 591380 534134 592000 534218
rect 591380 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592000 534134
rect 591380 498454 592000 533898
rect 591380 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592000 498454
rect 591380 498134 592000 498218
rect 591380 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592000 498134
rect 591380 462454 592000 497898
rect 591380 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592000 462454
rect 591380 462134 592000 462218
rect 591380 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592000 462134
rect 591380 426454 592000 461898
rect 591380 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592000 426454
rect 591380 426134 592000 426218
rect 591380 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592000 426134
rect 591380 390454 592000 425898
rect 591380 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592000 390454
rect 591380 390134 592000 390218
rect 591380 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592000 390134
rect 591380 354454 592000 389898
rect 591380 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592000 354454
rect 591380 354134 592000 354218
rect 591380 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592000 354134
rect 591380 318454 592000 353898
rect 591380 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592000 318454
rect 591380 318134 592000 318218
rect 591380 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592000 318134
rect 591380 282454 592000 317898
rect 591380 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592000 282454
rect 591380 282134 592000 282218
rect 591380 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592000 282134
rect 591380 246454 592000 281898
rect 591380 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592000 246454
rect 591380 246134 592000 246218
rect 591380 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592000 246134
rect 591380 210454 592000 245898
rect 591380 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592000 210454
rect 591380 210134 592000 210218
rect 591380 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592000 210134
rect 591380 174454 592000 209898
rect 591380 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592000 174454
rect 591380 174134 592000 174218
rect 591380 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592000 174134
rect 591380 138454 592000 173898
rect 591380 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592000 138454
rect 591380 138134 592000 138218
rect 591380 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592000 138134
rect 591380 102454 592000 137898
rect 591380 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592000 102454
rect 591380 102134 592000 102218
rect 591380 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592000 102134
rect 591380 66454 592000 101898
rect 591380 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592000 66454
rect 591380 66134 592000 66218
rect 591380 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592000 66134
rect 591380 30454 592000 65898
rect 591380 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592000 30454
rect 591380 30134 592000 30218
rect 591380 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592000 30134
rect 591380 -6416 592000 29898
rect 591380 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect 591380 -6736 592000 -6652
rect 591380 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect 591380 -7004 592000 -6972
rect 592340 682954 592960 711312
rect 592340 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect 592340 682634 592960 682718
rect 592340 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect 592340 646954 592960 682398
rect 592340 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect 592340 646634 592960 646718
rect 592340 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect 592340 610954 592960 646398
rect 592340 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect 592340 610634 592960 610718
rect 592340 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect 592340 574954 592960 610398
rect 592340 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect 592340 574634 592960 574718
rect 592340 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect 592340 538954 592960 574398
rect 592340 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect 592340 538634 592960 538718
rect 592340 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect 592340 502954 592960 538398
rect 592340 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect 592340 502634 592960 502718
rect 592340 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect 592340 466954 592960 502398
rect 592340 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect 592340 466634 592960 466718
rect 592340 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect 592340 430954 592960 466398
rect 592340 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect 592340 430634 592960 430718
rect 592340 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect 592340 394954 592960 430398
rect 592340 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect 592340 394634 592960 394718
rect 592340 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect 592340 358954 592960 394398
rect 592340 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect 592340 358634 592960 358718
rect 592340 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect 592340 322954 592960 358398
rect 592340 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect 592340 322634 592960 322718
rect 592340 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect 592340 286954 592960 322398
rect 592340 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect 592340 286634 592960 286718
rect 592340 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect 592340 250954 592960 286398
rect 592340 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect 592340 250634 592960 250718
rect 592340 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect 592340 214954 592960 250398
rect 592340 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect 592340 214634 592960 214718
rect 592340 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect 592340 178954 592960 214398
rect 592340 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect 592340 178634 592960 178718
rect 592340 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect 592340 142954 592960 178398
rect 592340 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect 592340 142634 592960 142718
rect 592340 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect 592340 106954 592960 142398
rect 592340 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect 592340 106634 592960 106718
rect 592340 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect 592340 70954 592960 106398
rect 592340 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect 592340 70634 592960 70718
rect 592340 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect 592340 34954 592960 70398
rect 592340 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect 592340 34634 592960 34718
rect 592340 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect 592340 -7376 592960 34398
rect 592340 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect 592340 -7696 592960 -7612
rect 592340 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect 592340 -7964 592960 -7932
<< via4 >>
rect -9004 711632 -8768 711868
rect -8684 711632 -8448 711868
rect -9004 711312 -8768 711548
rect -8684 711312 -8448 711548
rect -9004 682718 -8768 682954
rect -8684 682718 -8448 682954
rect -9004 682398 -8768 682634
rect -8684 682398 -8448 682634
rect -9004 646718 -8768 646954
rect -8684 646718 -8448 646954
rect -9004 646398 -8768 646634
rect -8684 646398 -8448 646634
rect -9004 610718 -8768 610954
rect -8684 610718 -8448 610954
rect -9004 610398 -8768 610634
rect -8684 610398 -8448 610634
rect -9004 574718 -8768 574954
rect -8684 574718 -8448 574954
rect -9004 574398 -8768 574634
rect -8684 574398 -8448 574634
rect -9004 538718 -8768 538954
rect -8684 538718 -8448 538954
rect -9004 538398 -8768 538634
rect -8684 538398 -8448 538634
rect -9004 502718 -8768 502954
rect -8684 502718 -8448 502954
rect -9004 502398 -8768 502634
rect -8684 502398 -8448 502634
rect -9004 466718 -8768 466954
rect -8684 466718 -8448 466954
rect -9004 466398 -8768 466634
rect -8684 466398 -8448 466634
rect -9004 430718 -8768 430954
rect -8684 430718 -8448 430954
rect -9004 430398 -8768 430634
rect -8684 430398 -8448 430634
rect -9004 394718 -8768 394954
rect -8684 394718 -8448 394954
rect -9004 394398 -8768 394634
rect -8684 394398 -8448 394634
rect -9004 358718 -8768 358954
rect -8684 358718 -8448 358954
rect -9004 358398 -8768 358634
rect -8684 358398 -8448 358634
rect -9004 322718 -8768 322954
rect -8684 322718 -8448 322954
rect -9004 322398 -8768 322634
rect -8684 322398 -8448 322634
rect -9004 286718 -8768 286954
rect -8684 286718 -8448 286954
rect -9004 286398 -8768 286634
rect -8684 286398 -8448 286634
rect -9004 250718 -8768 250954
rect -8684 250718 -8448 250954
rect -9004 250398 -8768 250634
rect -8684 250398 -8448 250634
rect -9004 214718 -8768 214954
rect -8684 214718 -8448 214954
rect -9004 214398 -8768 214634
rect -8684 214398 -8448 214634
rect -9004 178718 -8768 178954
rect -8684 178718 -8448 178954
rect -9004 178398 -8768 178634
rect -8684 178398 -8448 178634
rect -9004 142718 -8768 142954
rect -8684 142718 -8448 142954
rect -9004 142398 -8768 142634
rect -8684 142398 -8448 142634
rect -9004 106718 -8768 106954
rect -8684 106718 -8448 106954
rect -9004 106398 -8768 106634
rect -8684 106398 -8448 106634
rect -9004 70718 -8768 70954
rect -8684 70718 -8448 70954
rect -9004 70398 -8768 70634
rect -8684 70398 -8448 70634
rect -9004 34718 -8768 34954
rect -8684 34718 -8448 34954
rect -9004 34398 -8768 34634
rect -8684 34398 -8448 34634
rect -8044 710672 -7808 710908
rect -7724 710672 -7488 710908
rect -8044 710352 -7808 710588
rect -7724 710352 -7488 710588
rect -8044 678218 -7808 678454
rect -7724 678218 -7488 678454
rect -8044 677898 -7808 678134
rect -7724 677898 -7488 678134
rect -8044 642218 -7808 642454
rect -7724 642218 -7488 642454
rect -8044 641898 -7808 642134
rect -7724 641898 -7488 642134
rect -8044 606218 -7808 606454
rect -7724 606218 -7488 606454
rect -8044 605898 -7808 606134
rect -7724 605898 -7488 606134
rect -8044 570218 -7808 570454
rect -7724 570218 -7488 570454
rect -8044 569898 -7808 570134
rect -7724 569898 -7488 570134
rect -8044 534218 -7808 534454
rect -7724 534218 -7488 534454
rect -8044 533898 -7808 534134
rect -7724 533898 -7488 534134
rect -8044 498218 -7808 498454
rect -7724 498218 -7488 498454
rect -8044 497898 -7808 498134
rect -7724 497898 -7488 498134
rect -8044 462218 -7808 462454
rect -7724 462218 -7488 462454
rect -8044 461898 -7808 462134
rect -7724 461898 -7488 462134
rect -8044 426218 -7808 426454
rect -7724 426218 -7488 426454
rect -8044 425898 -7808 426134
rect -7724 425898 -7488 426134
rect -8044 390218 -7808 390454
rect -7724 390218 -7488 390454
rect -8044 389898 -7808 390134
rect -7724 389898 -7488 390134
rect -8044 354218 -7808 354454
rect -7724 354218 -7488 354454
rect -8044 353898 -7808 354134
rect -7724 353898 -7488 354134
rect -8044 318218 -7808 318454
rect -7724 318218 -7488 318454
rect -8044 317898 -7808 318134
rect -7724 317898 -7488 318134
rect -8044 282218 -7808 282454
rect -7724 282218 -7488 282454
rect -8044 281898 -7808 282134
rect -7724 281898 -7488 282134
rect -8044 246218 -7808 246454
rect -7724 246218 -7488 246454
rect -8044 245898 -7808 246134
rect -7724 245898 -7488 246134
rect -8044 210218 -7808 210454
rect -7724 210218 -7488 210454
rect -8044 209898 -7808 210134
rect -7724 209898 -7488 210134
rect -8044 174218 -7808 174454
rect -7724 174218 -7488 174454
rect -8044 173898 -7808 174134
rect -7724 173898 -7488 174134
rect -8044 138218 -7808 138454
rect -7724 138218 -7488 138454
rect -8044 137898 -7808 138134
rect -7724 137898 -7488 138134
rect -8044 102218 -7808 102454
rect -7724 102218 -7488 102454
rect -8044 101898 -7808 102134
rect -7724 101898 -7488 102134
rect -8044 66218 -7808 66454
rect -7724 66218 -7488 66454
rect -8044 65898 -7808 66134
rect -7724 65898 -7488 66134
rect -8044 30218 -7808 30454
rect -7724 30218 -7488 30454
rect -8044 29898 -7808 30134
rect -7724 29898 -7488 30134
rect -7084 709712 -6848 709948
rect -6764 709712 -6528 709948
rect -7084 709392 -6848 709628
rect -6764 709392 -6528 709628
rect -7084 673718 -6848 673954
rect -6764 673718 -6528 673954
rect -7084 673398 -6848 673634
rect -6764 673398 -6528 673634
rect -7084 637718 -6848 637954
rect -6764 637718 -6528 637954
rect -7084 637398 -6848 637634
rect -6764 637398 -6528 637634
rect -7084 601718 -6848 601954
rect -6764 601718 -6528 601954
rect -7084 601398 -6848 601634
rect -6764 601398 -6528 601634
rect -7084 565718 -6848 565954
rect -6764 565718 -6528 565954
rect -7084 565398 -6848 565634
rect -6764 565398 -6528 565634
rect -7084 529718 -6848 529954
rect -6764 529718 -6528 529954
rect -7084 529398 -6848 529634
rect -6764 529398 -6528 529634
rect -7084 493718 -6848 493954
rect -6764 493718 -6528 493954
rect -7084 493398 -6848 493634
rect -6764 493398 -6528 493634
rect -7084 457718 -6848 457954
rect -6764 457718 -6528 457954
rect -7084 457398 -6848 457634
rect -6764 457398 -6528 457634
rect -7084 421718 -6848 421954
rect -6764 421718 -6528 421954
rect -7084 421398 -6848 421634
rect -6764 421398 -6528 421634
rect -7084 385718 -6848 385954
rect -6764 385718 -6528 385954
rect -7084 385398 -6848 385634
rect -6764 385398 -6528 385634
rect -7084 349718 -6848 349954
rect -6764 349718 -6528 349954
rect -7084 349398 -6848 349634
rect -6764 349398 -6528 349634
rect -7084 313718 -6848 313954
rect -6764 313718 -6528 313954
rect -7084 313398 -6848 313634
rect -6764 313398 -6528 313634
rect -7084 277718 -6848 277954
rect -6764 277718 -6528 277954
rect -7084 277398 -6848 277634
rect -6764 277398 -6528 277634
rect -7084 241718 -6848 241954
rect -6764 241718 -6528 241954
rect -7084 241398 -6848 241634
rect -6764 241398 -6528 241634
rect -7084 205718 -6848 205954
rect -6764 205718 -6528 205954
rect -7084 205398 -6848 205634
rect -6764 205398 -6528 205634
rect -7084 169718 -6848 169954
rect -6764 169718 -6528 169954
rect -7084 169398 -6848 169634
rect -6764 169398 -6528 169634
rect -7084 133718 -6848 133954
rect -6764 133718 -6528 133954
rect -7084 133398 -6848 133634
rect -6764 133398 -6528 133634
rect -7084 97718 -6848 97954
rect -6764 97718 -6528 97954
rect -7084 97398 -6848 97634
rect -6764 97398 -6528 97634
rect -7084 61718 -6848 61954
rect -6764 61718 -6528 61954
rect -7084 61398 -6848 61634
rect -6764 61398 -6528 61634
rect -7084 25718 -6848 25954
rect -6764 25718 -6528 25954
rect -7084 25398 -6848 25634
rect -6764 25398 -6528 25634
rect -6124 708752 -5888 708988
rect -5804 708752 -5568 708988
rect -6124 708432 -5888 708668
rect -5804 708432 -5568 708668
rect -6124 669218 -5888 669454
rect -5804 669218 -5568 669454
rect -6124 668898 -5888 669134
rect -5804 668898 -5568 669134
rect -6124 633218 -5888 633454
rect -5804 633218 -5568 633454
rect -6124 632898 -5888 633134
rect -5804 632898 -5568 633134
rect -6124 597218 -5888 597454
rect -5804 597218 -5568 597454
rect -6124 596898 -5888 597134
rect -5804 596898 -5568 597134
rect -6124 561218 -5888 561454
rect -5804 561218 -5568 561454
rect -6124 560898 -5888 561134
rect -5804 560898 -5568 561134
rect -6124 525218 -5888 525454
rect -5804 525218 -5568 525454
rect -6124 524898 -5888 525134
rect -5804 524898 -5568 525134
rect -6124 489218 -5888 489454
rect -5804 489218 -5568 489454
rect -6124 488898 -5888 489134
rect -5804 488898 -5568 489134
rect -6124 453218 -5888 453454
rect -5804 453218 -5568 453454
rect -6124 452898 -5888 453134
rect -5804 452898 -5568 453134
rect -6124 417218 -5888 417454
rect -5804 417218 -5568 417454
rect -6124 416898 -5888 417134
rect -5804 416898 -5568 417134
rect -6124 381218 -5888 381454
rect -5804 381218 -5568 381454
rect -6124 380898 -5888 381134
rect -5804 380898 -5568 381134
rect -6124 345218 -5888 345454
rect -5804 345218 -5568 345454
rect -6124 344898 -5888 345134
rect -5804 344898 -5568 345134
rect -6124 309218 -5888 309454
rect -5804 309218 -5568 309454
rect -6124 308898 -5888 309134
rect -5804 308898 -5568 309134
rect -6124 273218 -5888 273454
rect -5804 273218 -5568 273454
rect -6124 272898 -5888 273134
rect -5804 272898 -5568 273134
rect -6124 237218 -5888 237454
rect -5804 237218 -5568 237454
rect -6124 236898 -5888 237134
rect -5804 236898 -5568 237134
rect -6124 201218 -5888 201454
rect -5804 201218 -5568 201454
rect -6124 200898 -5888 201134
rect -5804 200898 -5568 201134
rect -6124 165218 -5888 165454
rect -5804 165218 -5568 165454
rect -6124 164898 -5888 165134
rect -5804 164898 -5568 165134
rect -6124 129218 -5888 129454
rect -5804 129218 -5568 129454
rect -6124 128898 -5888 129134
rect -5804 128898 -5568 129134
rect -6124 93218 -5888 93454
rect -5804 93218 -5568 93454
rect -6124 92898 -5888 93134
rect -5804 92898 -5568 93134
rect -6124 57218 -5888 57454
rect -5804 57218 -5568 57454
rect -6124 56898 -5888 57134
rect -5804 56898 -5568 57134
rect -6124 21218 -5888 21454
rect -5804 21218 -5568 21454
rect -6124 20898 -5888 21134
rect -5804 20898 -5568 21134
rect -5164 707792 -4928 708028
rect -4844 707792 -4608 708028
rect -5164 707472 -4928 707708
rect -4844 707472 -4608 707708
rect -5164 700718 -4928 700954
rect -4844 700718 -4608 700954
rect -5164 700398 -4928 700634
rect -4844 700398 -4608 700634
rect -5164 664718 -4928 664954
rect -4844 664718 -4608 664954
rect -5164 664398 -4928 664634
rect -4844 664398 -4608 664634
rect -5164 628718 -4928 628954
rect -4844 628718 -4608 628954
rect -5164 628398 -4928 628634
rect -4844 628398 -4608 628634
rect -5164 592718 -4928 592954
rect -4844 592718 -4608 592954
rect -5164 592398 -4928 592634
rect -4844 592398 -4608 592634
rect -5164 556718 -4928 556954
rect -4844 556718 -4608 556954
rect -5164 556398 -4928 556634
rect -4844 556398 -4608 556634
rect -5164 520718 -4928 520954
rect -4844 520718 -4608 520954
rect -5164 520398 -4928 520634
rect -4844 520398 -4608 520634
rect -5164 484718 -4928 484954
rect -4844 484718 -4608 484954
rect -5164 484398 -4928 484634
rect -4844 484398 -4608 484634
rect -5164 448718 -4928 448954
rect -4844 448718 -4608 448954
rect -5164 448398 -4928 448634
rect -4844 448398 -4608 448634
rect -5164 412718 -4928 412954
rect -4844 412718 -4608 412954
rect -5164 412398 -4928 412634
rect -4844 412398 -4608 412634
rect -5164 376718 -4928 376954
rect -4844 376718 -4608 376954
rect -5164 376398 -4928 376634
rect -4844 376398 -4608 376634
rect -5164 340718 -4928 340954
rect -4844 340718 -4608 340954
rect -5164 340398 -4928 340634
rect -4844 340398 -4608 340634
rect -5164 304718 -4928 304954
rect -4844 304718 -4608 304954
rect -5164 304398 -4928 304634
rect -4844 304398 -4608 304634
rect -5164 268718 -4928 268954
rect -4844 268718 -4608 268954
rect -5164 268398 -4928 268634
rect -4844 268398 -4608 268634
rect -5164 232718 -4928 232954
rect -4844 232718 -4608 232954
rect -5164 232398 -4928 232634
rect -4844 232398 -4608 232634
rect -5164 196718 -4928 196954
rect -4844 196718 -4608 196954
rect -5164 196398 -4928 196634
rect -4844 196398 -4608 196634
rect -5164 160718 -4928 160954
rect -4844 160718 -4608 160954
rect -5164 160398 -4928 160634
rect -4844 160398 -4608 160634
rect -5164 124718 -4928 124954
rect -4844 124718 -4608 124954
rect -5164 124398 -4928 124634
rect -4844 124398 -4608 124634
rect -5164 88718 -4928 88954
rect -4844 88718 -4608 88954
rect -5164 88398 -4928 88634
rect -4844 88398 -4608 88634
rect -5164 52718 -4928 52954
rect -4844 52718 -4608 52954
rect -5164 52398 -4928 52634
rect -4844 52398 -4608 52634
rect -5164 16718 -4928 16954
rect -4844 16718 -4608 16954
rect -5164 16398 -4928 16634
rect -4844 16398 -4608 16634
rect -4204 706832 -3968 707068
rect -3884 706832 -3648 707068
rect -4204 706512 -3968 706748
rect -3884 706512 -3648 706748
rect -4204 696218 -3968 696454
rect -3884 696218 -3648 696454
rect -4204 695898 -3968 696134
rect -3884 695898 -3648 696134
rect -4204 660218 -3968 660454
rect -3884 660218 -3648 660454
rect -4204 659898 -3968 660134
rect -3884 659898 -3648 660134
rect -4204 624218 -3968 624454
rect -3884 624218 -3648 624454
rect -4204 623898 -3968 624134
rect -3884 623898 -3648 624134
rect -4204 588218 -3968 588454
rect -3884 588218 -3648 588454
rect -4204 587898 -3968 588134
rect -3884 587898 -3648 588134
rect -4204 552218 -3968 552454
rect -3884 552218 -3648 552454
rect -4204 551898 -3968 552134
rect -3884 551898 -3648 552134
rect -4204 516218 -3968 516454
rect -3884 516218 -3648 516454
rect -4204 515898 -3968 516134
rect -3884 515898 -3648 516134
rect -4204 480218 -3968 480454
rect -3884 480218 -3648 480454
rect -4204 479898 -3968 480134
rect -3884 479898 -3648 480134
rect -4204 444218 -3968 444454
rect -3884 444218 -3648 444454
rect -4204 443898 -3968 444134
rect -3884 443898 -3648 444134
rect -4204 408218 -3968 408454
rect -3884 408218 -3648 408454
rect -4204 407898 -3968 408134
rect -3884 407898 -3648 408134
rect -4204 372218 -3968 372454
rect -3884 372218 -3648 372454
rect -4204 371898 -3968 372134
rect -3884 371898 -3648 372134
rect -4204 336218 -3968 336454
rect -3884 336218 -3648 336454
rect -4204 335898 -3968 336134
rect -3884 335898 -3648 336134
rect -4204 300218 -3968 300454
rect -3884 300218 -3648 300454
rect -4204 299898 -3968 300134
rect -3884 299898 -3648 300134
rect -4204 264218 -3968 264454
rect -3884 264218 -3648 264454
rect -4204 263898 -3968 264134
rect -3884 263898 -3648 264134
rect -4204 228218 -3968 228454
rect -3884 228218 -3648 228454
rect -4204 227898 -3968 228134
rect -3884 227898 -3648 228134
rect -4204 192218 -3968 192454
rect -3884 192218 -3648 192454
rect -4204 191898 -3968 192134
rect -3884 191898 -3648 192134
rect -4204 156218 -3968 156454
rect -3884 156218 -3648 156454
rect -4204 155898 -3968 156134
rect -3884 155898 -3648 156134
rect -4204 120218 -3968 120454
rect -3884 120218 -3648 120454
rect -4204 119898 -3968 120134
rect -3884 119898 -3648 120134
rect -4204 84218 -3968 84454
rect -3884 84218 -3648 84454
rect -4204 83898 -3968 84134
rect -3884 83898 -3648 84134
rect -4204 48218 -3968 48454
rect -3884 48218 -3648 48454
rect -4204 47898 -3968 48134
rect -3884 47898 -3648 48134
rect -4204 12218 -3968 12454
rect -3884 12218 -3648 12454
rect -4204 11898 -3968 12134
rect -3884 11898 -3648 12134
rect -3244 705872 -3008 706108
rect -2924 705872 -2688 706108
rect -3244 705552 -3008 705788
rect -2924 705552 -2688 705788
rect -3244 691718 -3008 691954
rect -2924 691718 -2688 691954
rect -3244 691398 -3008 691634
rect -2924 691398 -2688 691634
rect -3244 655718 -3008 655954
rect -2924 655718 -2688 655954
rect -3244 655398 -3008 655634
rect -2924 655398 -2688 655634
rect -3244 619718 -3008 619954
rect -2924 619718 -2688 619954
rect -3244 619398 -3008 619634
rect -2924 619398 -2688 619634
rect -3244 583718 -3008 583954
rect -2924 583718 -2688 583954
rect -3244 583398 -3008 583634
rect -2924 583398 -2688 583634
rect -3244 547718 -3008 547954
rect -2924 547718 -2688 547954
rect -3244 547398 -3008 547634
rect -2924 547398 -2688 547634
rect -3244 511718 -3008 511954
rect -2924 511718 -2688 511954
rect -3244 511398 -3008 511634
rect -2924 511398 -2688 511634
rect -3244 475718 -3008 475954
rect -2924 475718 -2688 475954
rect -3244 475398 -3008 475634
rect -2924 475398 -2688 475634
rect -3244 439718 -3008 439954
rect -2924 439718 -2688 439954
rect -3244 439398 -3008 439634
rect -2924 439398 -2688 439634
rect -3244 403718 -3008 403954
rect -2924 403718 -2688 403954
rect -3244 403398 -3008 403634
rect -2924 403398 -2688 403634
rect -3244 367718 -3008 367954
rect -2924 367718 -2688 367954
rect -3244 367398 -3008 367634
rect -2924 367398 -2688 367634
rect -3244 331718 -3008 331954
rect -2924 331718 -2688 331954
rect -3244 331398 -3008 331634
rect -2924 331398 -2688 331634
rect -3244 295718 -3008 295954
rect -2924 295718 -2688 295954
rect -3244 295398 -3008 295634
rect -2924 295398 -2688 295634
rect -3244 259718 -3008 259954
rect -2924 259718 -2688 259954
rect -3244 259398 -3008 259634
rect -2924 259398 -2688 259634
rect -3244 223718 -3008 223954
rect -2924 223718 -2688 223954
rect -3244 223398 -3008 223634
rect -2924 223398 -2688 223634
rect -3244 187718 -3008 187954
rect -2924 187718 -2688 187954
rect -3244 187398 -3008 187634
rect -2924 187398 -2688 187634
rect -3244 151718 -3008 151954
rect -2924 151718 -2688 151954
rect -3244 151398 -3008 151634
rect -2924 151398 -2688 151634
rect -3244 115718 -3008 115954
rect -2924 115718 -2688 115954
rect -3244 115398 -3008 115634
rect -2924 115398 -2688 115634
rect -3244 79718 -3008 79954
rect -2924 79718 -2688 79954
rect -3244 79398 -3008 79634
rect -2924 79398 -2688 79634
rect -3244 43718 -3008 43954
rect -2924 43718 -2688 43954
rect -3244 43398 -3008 43634
rect -2924 43398 -2688 43634
rect -3244 7718 -3008 7954
rect -2924 7718 -2688 7954
rect -3244 7398 -3008 7634
rect -2924 7398 -2688 7634
rect -2284 704912 -2048 705148
rect -1964 704912 -1728 705148
rect -2284 704592 -2048 704828
rect -1964 704592 -1728 704828
rect -2284 687218 -2048 687454
rect -1964 687218 -1728 687454
rect -2284 686898 -2048 687134
rect -1964 686898 -1728 687134
rect -2284 651218 -2048 651454
rect -1964 651218 -1728 651454
rect -2284 650898 -2048 651134
rect -1964 650898 -1728 651134
rect -2284 615218 -2048 615454
rect -1964 615218 -1728 615454
rect -2284 614898 -2048 615134
rect -1964 614898 -1728 615134
rect -2284 579218 -2048 579454
rect -1964 579218 -1728 579454
rect -2284 578898 -2048 579134
rect -1964 578898 -1728 579134
rect -2284 543218 -2048 543454
rect -1964 543218 -1728 543454
rect -2284 542898 -2048 543134
rect -1964 542898 -1728 543134
rect -2284 507218 -2048 507454
rect -1964 507218 -1728 507454
rect -2284 506898 -2048 507134
rect -1964 506898 -1728 507134
rect -2284 471218 -2048 471454
rect -1964 471218 -1728 471454
rect -2284 470898 -2048 471134
rect -1964 470898 -1728 471134
rect -2284 435218 -2048 435454
rect -1964 435218 -1728 435454
rect -2284 434898 -2048 435134
rect -1964 434898 -1728 435134
rect -2284 399218 -2048 399454
rect -1964 399218 -1728 399454
rect -2284 398898 -2048 399134
rect -1964 398898 -1728 399134
rect -2284 363218 -2048 363454
rect -1964 363218 -1728 363454
rect -2284 362898 -2048 363134
rect -1964 362898 -1728 363134
rect -2284 327218 -2048 327454
rect -1964 327218 -1728 327454
rect -2284 326898 -2048 327134
rect -1964 326898 -1728 327134
rect -2284 291218 -2048 291454
rect -1964 291218 -1728 291454
rect -2284 290898 -2048 291134
rect -1964 290898 -1728 291134
rect -2284 255218 -2048 255454
rect -1964 255218 -1728 255454
rect -2284 254898 -2048 255134
rect -1964 254898 -1728 255134
rect -2284 219218 -2048 219454
rect -1964 219218 -1728 219454
rect -2284 218898 -2048 219134
rect -1964 218898 -1728 219134
rect -2284 183218 -2048 183454
rect -1964 183218 -1728 183454
rect -2284 182898 -2048 183134
rect -1964 182898 -1728 183134
rect -2284 147218 -2048 147454
rect -1964 147218 -1728 147454
rect -2284 146898 -2048 147134
rect -1964 146898 -1728 147134
rect -2284 111218 -2048 111454
rect -1964 111218 -1728 111454
rect -2284 110898 -2048 111134
rect -1964 110898 -1728 111134
rect -2284 75218 -2048 75454
rect -1964 75218 -1728 75454
rect -2284 74898 -2048 75134
rect -1964 74898 -1728 75134
rect -2284 39218 -2048 39454
rect -1964 39218 -1728 39454
rect -2284 38898 -2048 39134
rect -1964 38898 -1728 39134
rect -2284 3218 -2048 3454
rect -1964 3218 -1728 3454
rect -2284 2898 -2048 3134
rect -1964 2898 -1728 3134
rect -2284 -892 -2048 -656
rect -1964 -892 -1728 -656
rect -2284 -1212 -2048 -976
rect -1964 -1212 -1728 -976
rect 1826 704912 2062 705148
rect 2146 704912 2382 705148
rect 1826 704592 2062 704828
rect 2146 704592 2382 704828
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -892 2062 -656
rect 2146 -892 2382 -656
rect 1826 -1212 2062 -976
rect 2146 -1212 2382 -976
rect -3244 -1852 -3008 -1616
rect -2924 -1852 -2688 -1616
rect -3244 -2172 -3008 -1936
rect -2924 -2172 -2688 -1936
rect -4204 -2812 -3968 -2576
rect -3884 -2812 -3648 -2576
rect -4204 -3132 -3968 -2896
rect -3884 -3132 -3648 -2896
rect -5164 -3772 -4928 -3536
rect -4844 -3772 -4608 -3536
rect -5164 -4092 -4928 -3856
rect -4844 -4092 -4608 -3856
rect -6124 -4732 -5888 -4496
rect -5804 -4732 -5568 -4496
rect -6124 -5052 -5888 -4816
rect -5804 -5052 -5568 -4816
rect -7084 -5692 -6848 -5456
rect -6764 -5692 -6528 -5456
rect -7084 -6012 -6848 -5776
rect -6764 -6012 -6528 -5776
rect -8044 -6652 -7808 -6416
rect -7724 -6652 -7488 -6416
rect -8044 -6972 -7808 -6736
rect -7724 -6972 -7488 -6736
rect -9004 -7612 -8768 -7376
rect -8684 -7612 -8448 -7376
rect -9004 -7932 -8768 -7696
rect -8684 -7932 -8448 -7696
rect 6326 705872 6562 706108
rect 6646 705872 6882 706108
rect 6326 705552 6562 705788
rect 6646 705552 6882 705788
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1852 6562 -1616
rect 6646 -1852 6882 -1616
rect 6326 -2172 6562 -1936
rect 6646 -2172 6882 -1936
rect 10826 706832 11062 707068
rect 11146 706832 11382 707068
rect 10826 706512 11062 706748
rect 11146 706512 11382 706748
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2812 11062 -2576
rect 11146 -2812 11382 -2576
rect 10826 -3132 11062 -2896
rect 11146 -3132 11382 -2896
rect 15326 707792 15562 708028
rect 15646 707792 15882 708028
rect 15326 707472 15562 707708
rect 15646 707472 15882 707708
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3772 15562 -3536
rect 15646 -3772 15882 -3536
rect 15326 -4092 15562 -3856
rect 15646 -4092 15882 -3856
rect 19826 708752 20062 708988
rect 20146 708752 20382 708988
rect 19826 708432 20062 708668
rect 20146 708432 20382 708668
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4732 20062 -4496
rect 20146 -4732 20382 -4496
rect 19826 -5052 20062 -4816
rect 20146 -5052 20382 -4816
rect 24326 709712 24562 709948
rect 24646 709712 24882 709948
rect 24326 709392 24562 709628
rect 24646 709392 24882 709628
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5692 24562 -5456
rect 24646 -5692 24882 -5456
rect 24326 -6012 24562 -5776
rect 24646 -6012 24882 -5776
rect 28826 710672 29062 710908
rect 29146 710672 29382 710908
rect 28826 710352 29062 710588
rect 29146 710352 29382 710588
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6652 29062 -6416
rect 29146 -6652 29382 -6416
rect 28826 -6972 29062 -6736
rect 29146 -6972 29382 -6736
rect 33326 711632 33562 711868
rect 33646 711632 33882 711868
rect 33326 711312 33562 711548
rect 33646 711312 33882 711548
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7612 33562 -7376
rect 33646 -7612 33882 -7376
rect 33326 -7932 33562 -7696
rect 33646 -7932 33882 -7696
rect 37826 704912 38062 705148
rect 38146 704912 38382 705148
rect 37826 704592 38062 704828
rect 38146 704592 38382 704828
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -892 38062 -656
rect 38146 -892 38382 -656
rect 37826 -1212 38062 -976
rect 38146 -1212 38382 -976
rect 42326 705872 42562 706108
rect 42646 705872 42882 706108
rect 42326 705552 42562 705788
rect 42646 705552 42882 705788
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1852 42562 -1616
rect 42646 -1852 42882 -1616
rect 42326 -2172 42562 -1936
rect 42646 -2172 42882 -1936
rect 46826 706832 47062 707068
rect 47146 706832 47382 707068
rect 46826 706512 47062 706748
rect 47146 706512 47382 706748
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2812 47062 -2576
rect 47146 -2812 47382 -2576
rect 46826 -3132 47062 -2896
rect 47146 -3132 47382 -2896
rect 51326 707792 51562 708028
rect 51646 707792 51882 708028
rect 51326 707472 51562 707708
rect 51646 707472 51882 707708
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3772 51562 -3536
rect 51646 -3772 51882 -3536
rect 51326 -4092 51562 -3856
rect 51646 -4092 51882 -3856
rect 55826 708752 56062 708988
rect 56146 708752 56382 708988
rect 55826 708432 56062 708668
rect 56146 708432 56382 708668
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4732 56062 -4496
rect 56146 -4732 56382 -4496
rect 55826 -5052 56062 -4816
rect 56146 -5052 56382 -4816
rect 60326 709712 60562 709948
rect 60646 709712 60882 709948
rect 60326 709392 60562 709628
rect 60646 709392 60882 709628
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5692 60562 -5456
rect 60646 -5692 60882 -5456
rect 60326 -6012 60562 -5776
rect 60646 -6012 60882 -5776
rect 64826 710672 65062 710908
rect 65146 710672 65382 710908
rect 64826 710352 65062 710588
rect 65146 710352 65382 710588
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6652 65062 -6416
rect 65146 -6652 65382 -6416
rect 64826 -6972 65062 -6736
rect 65146 -6972 65382 -6736
rect 69326 711632 69562 711868
rect 69646 711632 69882 711868
rect 69326 711312 69562 711548
rect 69646 711312 69882 711548
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7612 69562 -7376
rect 69646 -7612 69882 -7376
rect 69326 -7932 69562 -7696
rect 69646 -7932 69882 -7696
rect 73826 704912 74062 705148
rect 74146 704912 74382 705148
rect 73826 704592 74062 704828
rect 74146 704592 74382 704828
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -892 74062 -656
rect 74146 -892 74382 -656
rect 73826 -1212 74062 -976
rect 74146 -1212 74382 -976
rect 78326 705872 78562 706108
rect 78646 705872 78882 706108
rect 78326 705552 78562 705788
rect 78646 705552 78882 705788
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1852 78562 -1616
rect 78646 -1852 78882 -1616
rect 78326 -2172 78562 -1936
rect 78646 -2172 78882 -1936
rect 82826 706832 83062 707068
rect 83146 706832 83382 707068
rect 82826 706512 83062 706748
rect 83146 706512 83382 706748
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2812 83062 -2576
rect 83146 -2812 83382 -2576
rect 82826 -3132 83062 -2896
rect 83146 -3132 83382 -2896
rect 87326 707792 87562 708028
rect 87646 707792 87882 708028
rect 87326 707472 87562 707708
rect 87646 707472 87882 707708
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3772 87562 -3536
rect 87646 -3772 87882 -3536
rect 87326 -4092 87562 -3856
rect 87646 -4092 87882 -3856
rect 91826 708752 92062 708988
rect 92146 708752 92382 708988
rect 91826 708432 92062 708668
rect 92146 708432 92382 708668
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4732 92062 -4496
rect 92146 -4732 92382 -4496
rect 91826 -5052 92062 -4816
rect 92146 -5052 92382 -4816
rect 96326 709712 96562 709948
rect 96646 709712 96882 709948
rect 96326 709392 96562 709628
rect 96646 709392 96882 709628
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 100826 710672 101062 710908
rect 101146 710672 101382 710908
rect 100826 710352 101062 710588
rect 101146 710352 101382 710588
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 105326 711632 105562 711868
rect 105646 711632 105882 711868
rect 105326 711312 105562 711548
rect 105646 711312 105882 711548
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 109826 704912 110062 705148
rect 110146 704912 110382 705148
rect 109826 704592 110062 704828
rect 110146 704592 110382 704828
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 114326 705872 114562 706108
rect 114646 705872 114882 706108
rect 114326 705552 114562 705788
rect 114646 705552 114882 705788
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 118826 706832 119062 707068
rect 119146 706832 119382 707068
rect 118826 706512 119062 706748
rect 119146 706512 119382 706748
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 123326 707792 123562 708028
rect 123646 707792 123882 708028
rect 123326 707472 123562 707708
rect 123646 707472 123882 707708
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 127826 708752 128062 708988
rect 128146 708752 128382 708988
rect 127826 708432 128062 708668
rect 128146 708432 128382 708668
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 132326 709712 132562 709948
rect 132646 709712 132882 709948
rect 132326 709392 132562 709628
rect 132646 709392 132882 709628
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 136826 710672 137062 710908
rect 137146 710672 137382 710908
rect 136826 710352 137062 710588
rect 137146 710352 137382 710588
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 141326 711632 141562 711868
rect 141646 711632 141882 711868
rect 141326 711312 141562 711548
rect 141646 711312 141882 711548
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 145826 704912 146062 705148
rect 146146 704912 146382 705148
rect 145826 704592 146062 704828
rect 146146 704592 146382 704828
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 150326 705872 150562 706108
rect 150646 705872 150882 706108
rect 150326 705552 150562 705788
rect 150646 705552 150882 705788
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 154826 706832 155062 707068
rect 155146 706832 155382 707068
rect 154826 706512 155062 706748
rect 155146 706512 155382 706748
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 159326 707792 159562 708028
rect 159646 707792 159882 708028
rect 159326 707472 159562 707708
rect 159646 707472 159882 707708
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 163826 708752 164062 708988
rect 164146 708752 164382 708988
rect 163826 708432 164062 708668
rect 164146 708432 164382 708668
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 168326 709712 168562 709948
rect 168646 709712 168882 709948
rect 168326 709392 168562 709628
rect 168646 709392 168882 709628
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 172826 710672 173062 710908
rect 173146 710672 173382 710908
rect 172826 710352 173062 710588
rect 173146 710352 173382 710588
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 119610 367718 119846 367954
rect 119610 367398 119846 367634
rect 150330 367718 150566 367954
rect 150330 367398 150566 367634
rect 104250 363218 104486 363454
rect 104250 362898 104486 363134
rect 134970 363218 135206 363454
rect 134970 362898 135206 363134
rect 165690 363218 165926 363454
rect 165690 362898 165926 363134
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 119610 331718 119846 331954
rect 119610 331398 119846 331634
rect 150330 331718 150566 331954
rect 150330 331398 150566 331634
rect 104250 327218 104486 327454
rect 104250 326898 104486 327134
rect 134970 327218 135206 327454
rect 134970 326898 135206 327134
rect 165690 327218 165926 327454
rect 165690 326898 165926 327134
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5692 96562 -5456
rect 96646 -5692 96882 -5456
rect 96326 -6012 96562 -5776
rect 96646 -6012 96882 -5776
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6652 101062 -6416
rect 101146 -6652 101382 -6416
rect 100826 -6972 101062 -6736
rect 101146 -6972 101382 -6736
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7612 105562 -7376
rect 105646 -7612 105882 -7376
rect 105326 -7932 105562 -7696
rect 105646 -7932 105882 -7696
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -892 110062 -656
rect 110146 -892 110382 -656
rect 109826 -1212 110062 -976
rect 110146 -1212 110382 -976
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1852 114562 -1616
rect 114646 -1852 114882 -1616
rect 114326 -2172 114562 -1936
rect 114646 -2172 114882 -1936
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2812 119062 -2576
rect 119146 -2812 119382 -2576
rect 118826 -3132 119062 -2896
rect 119146 -3132 119382 -2896
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3772 123562 -3536
rect 123646 -3772 123882 -3536
rect 123326 -4092 123562 -3856
rect 123646 -4092 123882 -3856
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4732 128062 -4496
rect 128146 -4732 128382 -4496
rect 127826 -5052 128062 -4816
rect 128146 -5052 128382 -4816
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5692 132562 -5456
rect 132646 -5692 132882 -5456
rect 132326 -6012 132562 -5776
rect 132646 -6012 132882 -5776
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6652 137062 -6416
rect 137146 -6652 137382 -6416
rect 136826 -6972 137062 -6736
rect 137146 -6972 137382 -6736
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7612 141562 -7376
rect 141646 -7612 141882 -7376
rect 141326 -7932 141562 -7696
rect 141646 -7932 141882 -7696
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -892 146062 -656
rect 146146 -892 146382 -656
rect 145826 -1212 146062 -976
rect 146146 -1212 146382 -976
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1852 150562 -1616
rect 150646 -1852 150882 -1616
rect 150326 -2172 150562 -1936
rect 150646 -2172 150882 -1936
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2812 155062 -2576
rect 155146 -2812 155382 -2576
rect 154826 -3132 155062 -2896
rect 155146 -3132 155382 -2896
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3772 159562 -3536
rect 159646 -3772 159882 -3536
rect 159326 -4092 159562 -3856
rect 159646 -4092 159882 -3856
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4732 164062 -4496
rect 164146 -4732 164382 -4496
rect 163826 -5052 164062 -4816
rect 164146 -5052 164382 -4816
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5692 168562 -5456
rect 168646 -5692 168882 -5456
rect 168326 -6012 168562 -5776
rect 168646 -6012 168882 -5776
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6652 173062 -6416
rect 173146 -6652 173382 -6416
rect 172826 -6972 173062 -6736
rect 173146 -6972 173382 -6736
rect 177326 711632 177562 711868
rect 177646 711632 177882 711868
rect 177326 711312 177562 711548
rect 177646 711312 177882 711548
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7612 177562 -7376
rect 177646 -7612 177882 -7376
rect 177326 -7932 177562 -7696
rect 177646 -7932 177882 -7696
rect 181826 704912 182062 705148
rect 182146 704912 182382 705148
rect 181826 704592 182062 704828
rect 182146 704592 182382 704828
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -892 182062 -656
rect 182146 -892 182382 -656
rect 181826 -1212 182062 -976
rect 182146 -1212 182382 -976
rect 186326 705872 186562 706108
rect 186646 705872 186882 706108
rect 186326 705552 186562 705788
rect 186646 705552 186882 705788
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1852 186562 -1616
rect 186646 -1852 186882 -1616
rect 186326 -2172 186562 -1936
rect 186646 -2172 186882 -1936
rect 190826 706832 191062 707068
rect 191146 706832 191382 707068
rect 190826 706512 191062 706748
rect 191146 706512 191382 706748
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2812 191062 -2576
rect 191146 -2812 191382 -2576
rect 190826 -3132 191062 -2896
rect 191146 -3132 191382 -2896
rect 195326 707792 195562 708028
rect 195646 707792 195882 708028
rect 195326 707472 195562 707708
rect 195646 707472 195882 707708
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3772 195562 -3536
rect 195646 -3772 195882 -3536
rect 195326 -4092 195562 -3856
rect 195646 -4092 195882 -3856
rect 199826 708752 200062 708988
rect 200146 708752 200382 708988
rect 199826 708432 200062 708668
rect 200146 708432 200382 708668
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4732 200062 -4496
rect 200146 -4732 200382 -4496
rect 199826 -5052 200062 -4816
rect 200146 -5052 200382 -4816
rect 204326 709712 204562 709948
rect 204646 709712 204882 709948
rect 204326 709392 204562 709628
rect 204646 709392 204882 709628
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5692 204562 -5456
rect 204646 -5692 204882 -5456
rect 204326 -6012 204562 -5776
rect 204646 -6012 204882 -5776
rect 208826 710672 209062 710908
rect 209146 710672 209382 710908
rect 208826 710352 209062 710588
rect 209146 710352 209382 710588
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6652 209062 -6416
rect 209146 -6652 209382 -6416
rect 208826 -6972 209062 -6736
rect 209146 -6972 209382 -6736
rect 213326 711632 213562 711868
rect 213646 711632 213882 711868
rect 213326 711312 213562 711548
rect 213646 711312 213882 711548
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704912 218062 705148
rect 218146 704912 218382 705148
rect 217826 704592 218062 704828
rect 218146 704592 218382 704828
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705872 222562 706108
rect 222646 705872 222882 706108
rect 222326 705552 222562 705788
rect 222646 705552 222882 705788
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706832 227062 707068
rect 227146 706832 227382 707068
rect 226826 706512 227062 706748
rect 227146 706512 227382 706748
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707792 231562 708028
rect 231646 707792 231882 708028
rect 231326 707472 231562 707708
rect 231646 707472 231882 707708
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708752 236062 708988
rect 236146 708752 236382 708988
rect 235826 708432 236062 708668
rect 236146 708432 236382 708668
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709712 240562 709948
rect 240646 709712 240882 709948
rect 240326 709392 240562 709628
rect 240646 709392 240882 709628
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710672 245062 710908
rect 245146 710672 245382 710908
rect 244826 710352 245062 710588
rect 245146 710352 245382 710588
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711632 249562 711868
rect 249646 711632 249882 711868
rect 249326 711312 249562 711548
rect 249646 711312 249882 711548
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704912 254062 705148
rect 254146 704912 254382 705148
rect 253826 704592 254062 704828
rect 254146 704592 254382 704828
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705872 258562 706108
rect 258646 705872 258882 706108
rect 258326 705552 258562 705788
rect 258646 705552 258882 705788
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706832 263062 707068
rect 263146 706832 263382 707068
rect 262826 706512 263062 706748
rect 263146 706512 263382 706748
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707792 267562 708028
rect 267646 707792 267882 708028
rect 267326 707472 267562 707708
rect 267646 707472 267882 707708
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708752 272062 708988
rect 272146 708752 272382 708988
rect 271826 708432 272062 708668
rect 272146 708432 272382 708668
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709712 276562 709948
rect 276646 709712 276882 709948
rect 276326 709392 276562 709628
rect 276646 709392 276882 709628
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710672 281062 710908
rect 281146 710672 281382 710908
rect 280826 710352 281062 710588
rect 281146 710352 281382 710588
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711632 285562 711868
rect 285646 711632 285882 711868
rect 285326 711312 285562 711548
rect 285646 711312 285882 711548
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704912 290062 705148
rect 290146 704912 290382 705148
rect 289826 704592 290062 704828
rect 290146 704592 290382 704828
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705872 294562 706108
rect 294646 705872 294882 706108
rect 294326 705552 294562 705788
rect 294646 705552 294882 705788
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706832 299062 707068
rect 299146 706832 299382 707068
rect 298826 706512 299062 706748
rect 299146 706512 299382 706748
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707792 303562 708028
rect 303646 707792 303882 708028
rect 303326 707472 303562 707708
rect 303646 707472 303882 707708
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708752 308062 708988
rect 308146 708752 308382 708988
rect 307826 708432 308062 708668
rect 308146 708432 308382 708668
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709712 312562 709948
rect 312646 709712 312882 709948
rect 312326 709392 312562 709628
rect 312646 709392 312882 709628
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710672 317062 710908
rect 317146 710672 317382 710908
rect 316826 710352 317062 710588
rect 317146 710352 317382 710588
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711632 321562 711868
rect 321646 711632 321882 711868
rect 321326 711312 321562 711548
rect 321646 711312 321882 711548
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704912 326062 705148
rect 326146 704912 326382 705148
rect 325826 704592 326062 704828
rect 326146 704592 326382 704828
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705872 330562 706108
rect 330646 705872 330882 706108
rect 330326 705552 330562 705788
rect 330646 705552 330882 705788
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706832 335062 707068
rect 335146 706832 335382 707068
rect 334826 706512 335062 706748
rect 335146 706512 335382 706748
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707792 339562 708028
rect 339646 707792 339882 708028
rect 339326 707472 339562 707708
rect 339646 707472 339882 707708
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708752 344062 708988
rect 344146 708752 344382 708988
rect 343826 708432 344062 708668
rect 344146 708432 344382 708668
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709712 348562 709948
rect 348646 709712 348882 709948
rect 348326 709392 348562 709628
rect 348646 709392 348882 709628
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710672 353062 710908
rect 353146 710672 353382 710908
rect 352826 710352 353062 710588
rect 353146 710352 353382 710588
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711632 357562 711868
rect 357646 711632 357882 711868
rect 357326 711312 357562 711548
rect 357646 711312 357882 711548
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704912 362062 705148
rect 362146 704912 362382 705148
rect 361826 704592 362062 704828
rect 362146 704592 362382 704828
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705872 366562 706108
rect 366646 705872 366882 706108
rect 366326 705552 366562 705788
rect 366646 705552 366882 705788
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 236650 435218 236886 435454
rect 236650 434898 236886 435134
rect 267370 435218 267606 435454
rect 267370 434898 267606 435134
rect 298090 435218 298326 435454
rect 298090 434898 298326 435134
rect 328810 435218 329046 435454
rect 328810 434898 329046 435134
rect 359530 435218 359766 435454
rect 359530 434898 359766 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 252010 403718 252246 403954
rect 252010 403398 252246 403634
rect 282730 403718 282966 403954
rect 282730 403398 282966 403634
rect 313450 403718 313686 403954
rect 313450 403398 313686 403634
rect 344170 403718 344406 403954
rect 344170 403398 344406 403634
rect 236650 399218 236886 399454
rect 236650 398898 236886 399134
rect 267370 399218 267606 399454
rect 267370 398898 267606 399134
rect 298090 399218 298326 399454
rect 298090 398898 298326 399134
rect 328810 399218 329046 399454
rect 328810 398898 329046 399134
rect 359530 399218 359766 399454
rect 359530 398898 359766 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 252010 367718 252246 367954
rect 252010 367398 252246 367634
rect 282730 367718 282966 367954
rect 282730 367398 282966 367634
rect 313450 367718 313686 367954
rect 313450 367398 313686 367634
rect 344170 367718 344406 367954
rect 344170 367398 344406 367634
rect 236650 363218 236886 363454
rect 236650 362898 236886 363134
rect 267370 363218 267606 363454
rect 267370 362898 267606 363134
rect 298090 363218 298326 363454
rect 298090 362898 298326 363134
rect 328810 363218 329046 363454
rect 328810 362898 329046 363134
rect 359530 363218 359766 363454
rect 359530 362898 359766 363134
rect 252010 331718 252246 331954
rect 252010 331398 252246 331634
rect 282730 331718 282966 331954
rect 282730 331398 282966 331634
rect 313450 331718 313686 331954
rect 313450 331398 313686 331634
rect 344170 331718 344406 331954
rect 344170 331398 344406 331634
rect 236650 327218 236886 327454
rect 236650 326898 236886 327134
rect 267370 327218 267606 327454
rect 267370 326898 267606 327134
rect 298090 327218 298326 327454
rect 298090 326898 298326 327134
rect 328810 327218 329046 327454
rect 328810 326898 329046 327134
rect 359530 327218 359766 327454
rect 359530 326898 359766 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 220328 223718 220564 223954
rect 220328 223398 220564 223634
rect 356056 223718 356292 223954
rect 356056 223398 356292 223634
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 187718 220564 187954
rect 220328 187398 220564 187634
rect 356056 187718 356292 187954
rect 356056 187398 356292 187634
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 213326 -7612 213562 -7376
rect 213646 -7612 213882 -7376
rect 213326 -7932 213562 -7696
rect 213646 -7932 213882 -7696
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -892 218062 -656
rect 218146 -892 218382 -656
rect 217826 -1212 218062 -976
rect 218146 -1212 218382 -976
rect 222326 -1852 222562 -1616
rect 222646 -1852 222882 -1616
rect 222326 -2172 222562 -1936
rect 222646 -2172 222882 -1936
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2812 227062 -2576
rect 227146 -2812 227382 -2576
rect 226826 -3132 227062 -2896
rect 227146 -3132 227382 -2896
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3772 231562 -3536
rect 231646 -3772 231882 -3536
rect 231326 -4092 231562 -3856
rect 231646 -4092 231882 -3856
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4732 236062 -4496
rect 236146 -4732 236382 -4496
rect 235826 -5052 236062 -4816
rect 236146 -5052 236382 -4816
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5692 240562 -5456
rect 240646 -5692 240882 -5456
rect 240326 -6012 240562 -5776
rect 240646 -6012 240882 -5776
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6652 245062 -6416
rect 245146 -6652 245382 -6416
rect 244826 -6972 245062 -6736
rect 245146 -6972 245382 -6736
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7612 249562 -7376
rect 249646 -7612 249882 -7376
rect 249326 -7932 249562 -7696
rect 249646 -7932 249882 -7696
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -892 254062 -656
rect 254146 -892 254382 -656
rect 253826 -1212 254062 -976
rect 254146 -1212 254382 -976
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1852 258562 -1616
rect 258646 -1852 258882 -1616
rect 258326 -2172 258562 -1936
rect 258646 -2172 258882 -1936
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2812 263062 -2576
rect 263146 -2812 263382 -2576
rect 262826 -3132 263062 -2896
rect 263146 -3132 263382 -2896
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3772 267562 -3536
rect 267646 -3772 267882 -3536
rect 267326 -4092 267562 -3856
rect 267646 -4092 267882 -3856
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4732 272062 -4496
rect 272146 -4732 272382 -4496
rect 271826 -5052 272062 -4816
rect 272146 -5052 272382 -4816
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5692 276562 -5456
rect 276646 -5692 276882 -5456
rect 276326 -6012 276562 -5776
rect 276646 -6012 276882 -5776
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6652 281062 -6416
rect 281146 -6652 281382 -6416
rect 280826 -6972 281062 -6736
rect 281146 -6972 281382 -6736
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7612 285562 -7376
rect 285646 -7612 285882 -7376
rect 285326 -7932 285562 -7696
rect 285646 -7932 285882 -7696
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -892 290062 -656
rect 290146 -892 290382 -656
rect 289826 -1212 290062 -976
rect 290146 -1212 290382 -976
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1852 294562 -1616
rect 294646 -1852 294882 -1616
rect 294326 -2172 294562 -1936
rect 294646 -2172 294882 -1936
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2812 299062 -2576
rect 299146 -2812 299382 -2576
rect 298826 -3132 299062 -2896
rect 299146 -3132 299382 -2896
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3772 303562 -3536
rect 303646 -3772 303882 -3536
rect 303326 -4092 303562 -3856
rect 303646 -4092 303882 -3856
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4732 308062 -4496
rect 308146 -4732 308382 -4496
rect 307826 -5052 308062 -4816
rect 308146 -5052 308382 -4816
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5692 312562 -5456
rect 312646 -5692 312882 -5456
rect 312326 -6012 312562 -5776
rect 312646 -6012 312882 -5776
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6652 317062 -6416
rect 317146 -6652 317382 -6416
rect 316826 -6972 317062 -6736
rect 317146 -6972 317382 -6736
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7612 321562 -7376
rect 321646 -7612 321882 -7376
rect 321326 -7932 321562 -7696
rect 321646 -7932 321882 -7696
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -892 326062 -656
rect 326146 -892 326382 -656
rect 325826 -1212 326062 -976
rect 326146 -1212 326382 -976
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1852 330562 -1616
rect 330646 -1852 330882 -1616
rect 330326 -2172 330562 -1936
rect 330646 -2172 330882 -1936
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2812 335062 -2576
rect 335146 -2812 335382 -2576
rect 334826 -3132 335062 -2896
rect 335146 -3132 335382 -2896
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3772 339562 -3536
rect 339646 -3772 339882 -3536
rect 339326 -4092 339562 -3856
rect 339646 -4092 339882 -3856
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4732 344062 -4496
rect 344146 -4732 344382 -4496
rect 343826 -5052 344062 -4816
rect 344146 -5052 344382 -4816
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5692 348562 -5456
rect 348646 -5692 348882 -5456
rect 348326 -6012 348562 -5776
rect 348646 -6012 348882 -5776
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 352826 -6652 353062 -6416
rect 353146 -6652 353382 -6416
rect 352826 -6972 353062 -6736
rect 353146 -6972 353382 -6736
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 357326 -7612 357562 -7376
rect 357646 -7612 357882 -7376
rect 357326 -7932 357562 -7696
rect 357646 -7932 357882 -7696
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 370826 706832 371062 707068
rect 371146 706832 371382 707068
rect 370826 706512 371062 706748
rect 371146 706512 371382 706748
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 361826 -892 362062 -656
rect 362146 -892 362382 -656
rect 361826 -1212 362062 -976
rect 362146 -1212 362382 -976
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 366326 -1852 366562 -1616
rect 366646 -1852 366882 -1616
rect 366326 -2172 366562 -1936
rect 366646 -2172 366882 -1936
rect 370826 -2812 371062 -2576
rect 371146 -2812 371382 -2576
rect 370826 -3132 371062 -2896
rect 371146 -3132 371382 -2896
rect 375326 707792 375562 708028
rect 375646 707792 375882 708028
rect 375326 707472 375562 707708
rect 375646 707472 375882 707708
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3772 375562 -3536
rect 375646 -3772 375882 -3536
rect 375326 -4092 375562 -3856
rect 375646 -4092 375882 -3856
rect 379826 708752 380062 708988
rect 380146 708752 380382 708988
rect 379826 708432 380062 708668
rect 380146 708432 380382 708668
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4732 380062 -4496
rect 380146 -4732 380382 -4496
rect 379826 -5052 380062 -4816
rect 380146 -5052 380382 -4816
rect 384326 709712 384562 709948
rect 384646 709712 384882 709948
rect 384326 709392 384562 709628
rect 384646 709392 384882 709628
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5692 384562 -5456
rect 384646 -5692 384882 -5456
rect 384326 -6012 384562 -5776
rect 384646 -6012 384882 -5776
rect 388826 710672 389062 710908
rect 389146 710672 389382 710908
rect 388826 710352 389062 710588
rect 389146 710352 389382 710588
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6652 389062 -6416
rect 389146 -6652 389382 -6416
rect 388826 -6972 389062 -6736
rect 389146 -6972 389382 -6736
rect 393326 711632 393562 711868
rect 393646 711632 393882 711868
rect 393326 711312 393562 711548
rect 393646 711312 393882 711548
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7612 393562 -7376
rect 393646 -7612 393882 -7376
rect 393326 -7932 393562 -7696
rect 393646 -7932 393882 -7696
rect 397826 704912 398062 705148
rect 398146 704912 398382 705148
rect 397826 704592 398062 704828
rect 398146 704592 398382 704828
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -892 398062 -656
rect 398146 -892 398382 -656
rect 397826 -1212 398062 -976
rect 398146 -1212 398382 -976
rect 402326 705872 402562 706108
rect 402646 705872 402882 706108
rect 402326 705552 402562 705788
rect 402646 705552 402882 705788
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1852 402562 -1616
rect 402646 -1852 402882 -1616
rect 402326 -2172 402562 -1936
rect 402646 -2172 402882 -1936
rect 406826 706832 407062 707068
rect 407146 706832 407382 707068
rect 406826 706512 407062 706748
rect 407146 706512 407382 706748
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2812 407062 -2576
rect 407146 -2812 407382 -2576
rect 406826 -3132 407062 -2896
rect 407146 -3132 407382 -2896
rect 411326 707792 411562 708028
rect 411646 707792 411882 708028
rect 411326 707472 411562 707708
rect 411646 707472 411882 707708
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3772 411562 -3536
rect 411646 -3772 411882 -3536
rect 411326 -4092 411562 -3856
rect 411646 -4092 411882 -3856
rect 415826 708752 416062 708988
rect 416146 708752 416382 708988
rect 415826 708432 416062 708668
rect 416146 708432 416382 708668
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4732 416062 -4496
rect 416146 -4732 416382 -4496
rect 415826 -5052 416062 -4816
rect 416146 -5052 416382 -4816
rect 420326 709712 420562 709948
rect 420646 709712 420882 709948
rect 420326 709392 420562 709628
rect 420646 709392 420882 709628
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5692 420562 -5456
rect 420646 -5692 420882 -5456
rect 420326 -6012 420562 -5776
rect 420646 -6012 420882 -5776
rect 424826 710672 425062 710908
rect 425146 710672 425382 710908
rect 424826 710352 425062 710588
rect 425146 710352 425382 710588
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6652 425062 -6416
rect 425146 -6652 425382 -6416
rect 424826 -6972 425062 -6736
rect 425146 -6972 425382 -6736
rect 429326 711632 429562 711868
rect 429646 711632 429882 711868
rect 429326 711312 429562 711548
rect 429646 711312 429882 711548
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7612 429562 -7376
rect 429646 -7612 429882 -7376
rect 429326 -7932 429562 -7696
rect 429646 -7932 429882 -7696
rect 433826 704912 434062 705148
rect 434146 704912 434382 705148
rect 433826 704592 434062 704828
rect 434146 704592 434382 704828
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -892 434062 -656
rect 434146 -892 434382 -656
rect 433826 -1212 434062 -976
rect 434146 -1212 434382 -976
rect 438326 705872 438562 706108
rect 438646 705872 438882 706108
rect 438326 705552 438562 705788
rect 438646 705552 438882 705788
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1852 438562 -1616
rect 438646 -1852 438882 -1616
rect 438326 -2172 438562 -1936
rect 438646 -2172 438882 -1936
rect 442826 706832 443062 707068
rect 443146 706832 443382 707068
rect 442826 706512 443062 706748
rect 443146 706512 443382 706748
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2812 443062 -2576
rect 443146 -2812 443382 -2576
rect 442826 -3132 443062 -2896
rect 443146 -3132 443382 -2896
rect 447326 707792 447562 708028
rect 447646 707792 447882 708028
rect 447326 707472 447562 707708
rect 447646 707472 447882 707708
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3772 447562 -3536
rect 447646 -3772 447882 -3536
rect 447326 -4092 447562 -3856
rect 447646 -4092 447882 -3856
rect 451826 708752 452062 708988
rect 452146 708752 452382 708988
rect 451826 708432 452062 708668
rect 452146 708432 452382 708668
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4732 452062 -4496
rect 452146 -4732 452382 -4496
rect 451826 -5052 452062 -4816
rect 452146 -5052 452382 -4816
rect 456326 709712 456562 709948
rect 456646 709712 456882 709948
rect 456326 709392 456562 709628
rect 456646 709392 456882 709628
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5692 456562 -5456
rect 456646 -5692 456882 -5456
rect 456326 -6012 456562 -5776
rect 456646 -6012 456882 -5776
rect 460826 710672 461062 710908
rect 461146 710672 461382 710908
rect 460826 710352 461062 710588
rect 461146 710352 461382 710588
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6652 461062 -6416
rect 461146 -6652 461382 -6416
rect 460826 -6972 461062 -6736
rect 461146 -6972 461382 -6736
rect 465326 711632 465562 711868
rect 465646 711632 465882 711868
rect 465326 711312 465562 711548
rect 465646 711312 465882 711548
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7612 465562 -7376
rect 465646 -7612 465882 -7376
rect 465326 -7932 465562 -7696
rect 465646 -7932 465882 -7696
rect 469826 704912 470062 705148
rect 470146 704912 470382 705148
rect 469826 704592 470062 704828
rect 470146 704592 470382 704828
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -892 470062 -656
rect 470146 -892 470382 -656
rect 469826 -1212 470062 -976
rect 470146 -1212 470382 -976
rect 474326 705872 474562 706108
rect 474646 705872 474882 706108
rect 474326 705552 474562 705788
rect 474646 705552 474882 705788
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1852 474562 -1616
rect 474646 -1852 474882 -1616
rect 474326 -2172 474562 -1936
rect 474646 -2172 474882 -1936
rect 478826 706832 479062 707068
rect 479146 706832 479382 707068
rect 478826 706512 479062 706748
rect 479146 706512 479382 706748
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2812 479062 -2576
rect 479146 -2812 479382 -2576
rect 478826 -3132 479062 -2896
rect 479146 -3132 479382 -2896
rect 483326 707792 483562 708028
rect 483646 707792 483882 708028
rect 483326 707472 483562 707708
rect 483646 707472 483882 707708
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3772 483562 -3536
rect 483646 -3772 483882 -3536
rect 483326 -4092 483562 -3856
rect 483646 -4092 483882 -3856
rect 487826 708752 488062 708988
rect 488146 708752 488382 708988
rect 487826 708432 488062 708668
rect 488146 708432 488382 708668
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4732 488062 -4496
rect 488146 -4732 488382 -4496
rect 487826 -5052 488062 -4816
rect 488146 -5052 488382 -4816
rect 492326 709712 492562 709948
rect 492646 709712 492882 709948
rect 492326 709392 492562 709628
rect 492646 709392 492882 709628
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5692 492562 -5456
rect 492646 -5692 492882 -5456
rect 492326 -6012 492562 -5776
rect 492646 -6012 492882 -5776
rect 496826 710672 497062 710908
rect 497146 710672 497382 710908
rect 496826 710352 497062 710588
rect 497146 710352 497382 710588
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6652 497062 -6416
rect 497146 -6652 497382 -6416
rect 496826 -6972 497062 -6736
rect 497146 -6972 497382 -6736
rect 501326 711632 501562 711868
rect 501646 711632 501882 711868
rect 501326 711312 501562 711548
rect 501646 711312 501882 711548
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7612 501562 -7376
rect 501646 -7612 501882 -7376
rect 501326 -7932 501562 -7696
rect 501646 -7932 501882 -7696
rect 505826 704912 506062 705148
rect 506146 704912 506382 705148
rect 505826 704592 506062 704828
rect 506146 704592 506382 704828
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -892 506062 -656
rect 506146 -892 506382 -656
rect 505826 -1212 506062 -976
rect 506146 -1212 506382 -976
rect 510326 705872 510562 706108
rect 510646 705872 510882 706108
rect 510326 705552 510562 705788
rect 510646 705552 510882 705788
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1852 510562 -1616
rect 510646 -1852 510882 -1616
rect 510326 -2172 510562 -1936
rect 510646 -2172 510882 -1936
rect 514826 706832 515062 707068
rect 515146 706832 515382 707068
rect 514826 706512 515062 706748
rect 515146 706512 515382 706748
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2812 515062 -2576
rect 515146 -2812 515382 -2576
rect 514826 -3132 515062 -2896
rect 515146 -3132 515382 -2896
rect 519326 707792 519562 708028
rect 519646 707792 519882 708028
rect 519326 707472 519562 707708
rect 519646 707472 519882 707708
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3772 519562 -3536
rect 519646 -3772 519882 -3536
rect 519326 -4092 519562 -3856
rect 519646 -4092 519882 -3856
rect 523826 708752 524062 708988
rect 524146 708752 524382 708988
rect 523826 708432 524062 708668
rect 524146 708432 524382 708668
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4732 524062 -4496
rect 524146 -4732 524382 -4496
rect 523826 -5052 524062 -4816
rect 524146 -5052 524382 -4816
rect 528326 709712 528562 709948
rect 528646 709712 528882 709948
rect 528326 709392 528562 709628
rect 528646 709392 528882 709628
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5692 528562 -5456
rect 528646 -5692 528882 -5456
rect 528326 -6012 528562 -5776
rect 528646 -6012 528882 -5776
rect 532826 710672 533062 710908
rect 533146 710672 533382 710908
rect 532826 710352 533062 710588
rect 533146 710352 533382 710588
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6652 533062 -6416
rect 533146 -6652 533382 -6416
rect 532826 -6972 533062 -6736
rect 533146 -6972 533382 -6736
rect 537326 711632 537562 711868
rect 537646 711632 537882 711868
rect 537326 711312 537562 711548
rect 537646 711312 537882 711548
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7612 537562 -7376
rect 537646 -7612 537882 -7376
rect 537326 -7932 537562 -7696
rect 537646 -7932 537882 -7696
rect 541826 704912 542062 705148
rect 542146 704912 542382 705148
rect 541826 704592 542062 704828
rect 542146 704592 542382 704828
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -892 542062 -656
rect 542146 -892 542382 -656
rect 541826 -1212 542062 -976
rect 542146 -1212 542382 -976
rect 546326 705872 546562 706108
rect 546646 705872 546882 706108
rect 546326 705552 546562 705788
rect 546646 705552 546882 705788
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1852 546562 -1616
rect 546646 -1852 546882 -1616
rect 546326 -2172 546562 -1936
rect 546646 -2172 546882 -1936
rect 550826 706832 551062 707068
rect 551146 706832 551382 707068
rect 550826 706512 551062 706748
rect 551146 706512 551382 706748
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2812 551062 -2576
rect 551146 -2812 551382 -2576
rect 550826 -3132 551062 -2896
rect 551146 -3132 551382 -2896
rect 555326 707792 555562 708028
rect 555646 707792 555882 708028
rect 555326 707472 555562 707708
rect 555646 707472 555882 707708
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3772 555562 -3536
rect 555646 -3772 555882 -3536
rect 555326 -4092 555562 -3856
rect 555646 -4092 555882 -3856
rect 559826 708752 560062 708988
rect 560146 708752 560382 708988
rect 559826 708432 560062 708668
rect 560146 708432 560382 708668
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4732 560062 -4496
rect 560146 -4732 560382 -4496
rect 559826 -5052 560062 -4816
rect 560146 -5052 560382 -4816
rect 564326 709712 564562 709948
rect 564646 709712 564882 709948
rect 564326 709392 564562 709628
rect 564646 709392 564882 709628
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5692 564562 -5456
rect 564646 -5692 564882 -5456
rect 564326 -6012 564562 -5776
rect 564646 -6012 564882 -5776
rect 568826 710672 569062 710908
rect 569146 710672 569382 710908
rect 568826 710352 569062 710588
rect 569146 710352 569382 710588
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6652 569062 -6416
rect 569146 -6652 569382 -6416
rect 568826 -6972 569062 -6736
rect 569146 -6972 569382 -6736
rect 573326 711632 573562 711868
rect 573646 711632 573882 711868
rect 573326 711312 573562 711548
rect 573646 711312 573882 711548
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7612 573562 -7376
rect 573646 -7612 573882 -7376
rect 573326 -7932 573562 -7696
rect 573646 -7932 573882 -7696
rect 577826 704912 578062 705148
rect 578146 704912 578382 705148
rect 577826 704592 578062 704828
rect 578146 704592 578382 704828
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -892 578062 -656
rect 578146 -892 578382 -656
rect 577826 -1212 578062 -976
rect 578146 -1212 578382 -976
rect 592372 711632 592608 711868
rect 592692 711632 592928 711868
rect 592372 711312 592608 711548
rect 592692 711312 592928 711548
rect 591412 710672 591648 710908
rect 591732 710672 591968 710908
rect 591412 710352 591648 710588
rect 591732 710352 591968 710588
rect 590452 709712 590688 709948
rect 590772 709712 591008 709948
rect 590452 709392 590688 709628
rect 590772 709392 591008 709628
rect 589492 708752 589728 708988
rect 589812 708752 590048 708988
rect 589492 708432 589728 708668
rect 589812 708432 590048 708668
rect 588532 707792 588768 708028
rect 588852 707792 589088 708028
rect 588532 707472 588768 707708
rect 588852 707472 589088 707708
rect 587572 706832 587808 707068
rect 587892 706832 588128 707068
rect 587572 706512 587808 706748
rect 587892 706512 588128 706748
rect 582326 705872 582562 706108
rect 582646 705872 582882 706108
rect 582326 705552 582562 705788
rect 582646 705552 582882 705788
rect 586612 705872 586848 706108
rect 586932 705872 587168 706108
rect 586612 705552 586848 705788
rect 586932 705552 587168 705788
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585652 704912 585888 705148
rect 585972 704912 586208 705148
rect 585652 704592 585888 704828
rect 585972 704592 586208 704828
rect 585652 687218 585888 687454
rect 585972 687218 586208 687454
rect 585652 686898 585888 687134
rect 585972 686898 586208 687134
rect 585652 651218 585888 651454
rect 585972 651218 586208 651454
rect 585652 650898 585888 651134
rect 585972 650898 586208 651134
rect 585652 615218 585888 615454
rect 585972 615218 586208 615454
rect 585652 614898 585888 615134
rect 585972 614898 586208 615134
rect 585652 579218 585888 579454
rect 585972 579218 586208 579454
rect 585652 578898 585888 579134
rect 585972 578898 586208 579134
rect 585652 543218 585888 543454
rect 585972 543218 586208 543454
rect 585652 542898 585888 543134
rect 585972 542898 586208 543134
rect 585652 507218 585888 507454
rect 585972 507218 586208 507454
rect 585652 506898 585888 507134
rect 585972 506898 586208 507134
rect 585652 471218 585888 471454
rect 585972 471218 586208 471454
rect 585652 470898 585888 471134
rect 585972 470898 586208 471134
rect 585652 435218 585888 435454
rect 585972 435218 586208 435454
rect 585652 434898 585888 435134
rect 585972 434898 586208 435134
rect 585652 399218 585888 399454
rect 585972 399218 586208 399454
rect 585652 398898 585888 399134
rect 585972 398898 586208 399134
rect 585652 363218 585888 363454
rect 585972 363218 586208 363454
rect 585652 362898 585888 363134
rect 585972 362898 586208 363134
rect 585652 327218 585888 327454
rect 585972 327218 586208 327454
rect 585652 326898 585888 327134
rect 585972 326898 586208 327134
rect 585652 291218 585888 291454
rect 585972 291218 586208 291454
rect 585652 290898 585888 291134
rect 585972 290898 586208 291134
rect 585652 255218 585888 255454
rect 585972 255218 586208 255454
rect 585652 254898 585888 255134
rect 585972 254898 586208 255134
rect 585652 219218 585888 219454
rect 585972 219218 586208 219454
rect 585652 218898 585888 219134
rect 585972 218898 586208 219134
rect 585652 183218 585888 183454
rect 585972 183218 586208 183454
rect 585652 182898 585888 183134
rect 585972 182898 586208 183134
rect 585652 147218 585888 147454
rect 585972 147218 586208 147454
rect 585652 146898 585888 147134
rect 585972 146898 586208 147134
rect 585652 111218 585888 111454
rect 585972 111218 586208 111454
rect 585652 110898 585888 111134
rect 585972 110898 586208 111134
rect 585652 75218 585888 75454
rect 585972 75218 586208 75454
rect 585652 74898 585888 75134
rect 585972 74898 586208 75134
rect 585652 39218 585888 39454
rect 585972 39218 586208 39454
rect 585652 38898 585888 39134
rect 585972 38898 586208 39134
rect 585652 3218 585888 3454
rect 585972 3218 586208 3454
rect 585652 2898 585888 3134
rect 585972 2898 586208 3134
rect 585652 -892 585888 -656
rect 585972 -892 586208 -656
rect 585652 -1212 585888 -976
rect 585972 -1212 586208 -976
rect 586612 691718 586848 691954
rect 586932 691718 587168 691954
rect 586612 691398 586848 691634
rect 586932 691398 587168 691634
rect 586612 655718 586848 655954
rect 586932 655718 587168 655954
rect 586612 655398 586848 655634
rect 586932 655398 587168 655634
rect 586612 619718 586848 619954
rect 586932 619718 587168 619954
rect 586612 619398 586848 619634
rect 586932 619398 587168 619634
rect 586612 583718 586848 583954
rect 586932 583718 587168 583954
rect 586612 583398 586848 583634
rect 586932 583398 587168 583634
rect 586612 547718 586848 547954
rect 586932 547718 587168 547954
rect 586612 547398 586848 547634
rect 586932 547398 587168 547634
rect 586612 511718 586848 511954
rect 586932 511718 587168 511954
rect 586612 511398 586848 511634
rect 586932 511398 587168 511634
rect 586612 475718 586848 475954
rect 586932 475718 587168 475954
rect 586612 475398 586848 475634
rect 586932 475398 587168 475634
rect 586612 439718 586848 439954
rect 586932 439718 587168 439954
rect 586612 439398 586848 439634
rect 586932 439398 587168 439634
rect 586612 403718 586848 403954
rect 586932 403718 587168 403954
rect 586612 403398 586848 403634
rect 586932 403398 587168 403634
rect 586612 367718 586848 367954
rect 586932 367718 587168 367954
rect 586612 367398 586848 367634
rect 586932 367398 587168 367634
rect 586612 331718 586848 331954
rect 586932 331718 587168 331954
rect 586612 331398 586848 331634
rect 586932 331398 587168 331634
rect 586612 295718 586848 295954
rect 586932 295718 587168 295954
rect 586612 295398 586848 295634
rect 586932 295398 587168 295634
rect 586612 259718 586848 259954
rect 586932 259718 587168 259954
rect 586612 259398 586848 259634
rect 586932 259398 587168 259634
rect 586612 223718 586848 223954
rect 586932 223718 587168 223954
rect 586612 223398 586848 223634
rect 586932 223398 587168 223634
rect 586612 187718 586848 187954
rect 586932 187718 587168 187954
rect 586612 187398 586848 187634
rect 586932 187398 587168 187634
rect 586612 151718 586848 151954
rect 586932 151718 587168 151954
rect 586612 151398 586848 151634
rect 586932 151398 587168 151634
rect 586612 115718 586848 115954
rect 586932 115718 587168 115954
rect 586612 115398 586848 115634
rect 586932 115398 587168 115634
rect 586612 79718 586848 79954
rect 586932 79718 587168 79954
rect 586612 79398 586848 79634
rect 586932 79398 587168 79634
rect 586612 43718 586848 43954
rect 586932 43718 587168 43954
rect 586612 43398 586848 43634
rect 586932 43398 587168 43634
rect 586612 7718 586848 7954
rect 586932 7718 587168 7954
rect 586612 7398 586848 7634
rect 586932 7398 587168 7634
rect 582326 -1852 582562 -1616
rect 582646 -1852 582882 -1616
rect 582326 -2172 582562 -1936
rect 582646 -2172 582882 -1936
rect 586612 -1852 586848 -1616
rect 586932 -1852 587168 -1616
rect 586612 -2172 586848 -1936
rect 586932 -2172 587168 -1936
rect 587572 696218 587808 696454
rect 587892 696218 588128 696454
rect 587572 695898 587808 696134
rect 587892 695898 588128 696134
rect 587572 660218 587808 660454
rect 587892 660218 588128 660454
rect 587572 659898 587808 660134
rect 587892 659898 588128 660134
rect 587572 624218 587808 624454
rect 587892 624218 588128 624454
rect 587572 623898 587808 624134
rect 587892 623898 588128 624134
rect 587572 588218 587808 588454
rect 587892 588218 588128 588454
rect 587572 587898 587808 588134
rect 587892 587898 588128 588134
rect 587572 552218 587808 552454
rect 587892 552218 588128 552454
rect 587572 551898 587808 552134
rect 587892 551898 588128 552134
rect 587572 516218 587808 516454
rect 587892 516218 588128 516454
rect 587572 515898 587808 516134
rect 587892 515898 588128 516134
rect 587572 480218 587808 480454
rect 587892 480218 588128 480454
rect 587572 479898 587808 480134
rect 587892 479898 588128 480134
rect 587572 444218 587808 444454
rect 587892 444218 588128 444454
rect 587572 443898 587808 444134
rect 587892 443898 588128 444134
rect 587572 408218 587808 408454
rect 587892 408218 588128 408454
rect 587572 407898 587808 408134
rect 587892 407898 588128 408134
rect 587572 372218 587808 372454
rect 587892 372218 588128 372454
rect 587572 371898 587808 372134
rect 587892 371898 588128 372134
rect 587572 336218 587808 336454
rect 587892 336218 588128 336454
rect 587572 335898 587808 336134
rect 587892 335898 588128 336134
rect 587572 300218 587808 300454
rect 587892 300218 588128 300454
rect 587572 299898 587808 300134
rect 587892 299898 588128 300134
rect 587572 264218 587808 264454
rect 587892 264218 588128 264454
rect 587572 263898 587808 264134
rect 587892 263898 588128 264134
rect 587572 228218 587808 228454
rect 587892 228218 588128 228454
rect 587572 227898 587808 228134
rect 587892 227898 588128 228134
rect 587572 192218 587808 192454
rect 587892 192218 588128 192454
rect 587572 191898 587808 192134
rect 587892 191898 588128 192134
rect 587572 156218 587808 156454
rect 587892 156218 588128 156454
rect 587572 155898 587808 156134
rect 587892 155898 588128 156134
rect 587572 120218 587808 120454
rect 587892 120218 588128 120454
rect 587572 119898 587808 120134
rect 587892 119898 588128 120134
rect 587572 84218 587808 84454
rect 587892 84218 588128 84454
rect 587572 83898 587808 84134
rect 587892 83898 588128 84134
rect 587572 48218 587808 48454
rect 587892 48218 588128 48454
rect 587572 47898 587808 48134
rect 587892 47898 588128 48134
rect 587572 12218 587808 12454
rect 587892 12218 588128 12454
rect 587572 11898 587808 12134
rect 587892 11898 588128 12134
rect 587572 -2812 587808 -2576
rect 587892 -2812 588128 -2576
rect 587572 -3132 587808 -2896
rect 587892 -3132 588128 -2896
rect 588532 700718 588768 700954
rect 588852 700718 589088 700954
rect 588532 700398 588768 700634
rect 588852 700398 589088 700634
rect 588532 664718 588768 664954
rect 588852 664718 589088 664954
rect 588532 664398 588768 664634
rect 588852 664398 589088 664634
rect 588532 628718 588768 628954
rect 588852 628718 589088 628954
rect 588532 628398 588768 628634
rect 588852 628398 589088 628634
rect 588532 592718 588768 592954
rect 588852 592718 589088 592954
rect 588532 592398 588768 592634
rect 588852 592398 589088 592634
rect 588532 556718 588768 556954
rect 588852 556718 589088 556954
rect 588532 556398 588768 556634
rect 588852 556398 589088 556634
rect 588532 520718 588768 520954
rect 588852 520718 589088 520954
rect 588532 520398 588768 520634
rect 588852 520398 589088 520634
rect 588532 484718 588768 484954
rect 588852 484718 589088 484954
rect 588532 484398 588768 484634
rect 588852 484398 589088 484634
rect 588532 448718 588768 448954
rect 588852 448718 589088 448954
rect 588532 448398 588768 448634
rect 588852 448398 589088 448634
rect 588532 412718 588768 412954
rect 588852 412718 589088 412954
rect 588532 412398 588768 412634
rect 588852 412398 589088 412634
rect 588532 376718 588768 376954
rect 588852 376718 589088 376954
rect 588532 376398 588768 376634
rect 588852 376398 589088 376634
rect 588532 340718 588768 340954
rect 588852 340718 589088 340954
rect 588532 340398 588768 340634
rect 588852 340398 589088 340634
rect 588532 304718 588768 304954
rect 588852 304718 589088 304954
rect 588532 304398 588768 304634
rect 588852 304398 589088 304634
rect 588532 268718 588768 268954
rect 588852 268718 589088 268954
rect 588532 268398 588768 268634
rect 588852 268398 589088 268634
rect 588532 232718 588768 232954
rect 588852 232718 589088 232954
rect 588532 232398 588768 232634
rect 588852 232398 589088 232634
rect 588532 196718 588768 196954
rect 588852 196718 589088 196954
rect 588532 196398 588768 196634
rect 588852 196398 589088 196634
rect 588532 160718 588768 160954
rect 588852 160718 589088 160954
rect 588532 160398 588768 160634
rect 588852 160398 589088 160634
rect 588532 124718 588768 124954
rect 588852 124718 589088 124954
rect 588532 124398 588768 124634
rect 588852 124398 589088 124634
rect 588532 88718 588768 88954
rect 588852 88718 589088 88954
rect 588532 88398 588768 88634
rect 588852 88398 589088 88634
rect 588532 52718 588768 52954
rect 588852 52718 589088 52954
rect 588532 52398 588768 52634
rect 588852 52398 589088 52634
rect 588532 16718 588768 16954
rect 588852 16718 589088 16954
rect 588532 16398 588768 16634
rect 588852 16398 589088 16634
rect 588532 -3772 588768 -3536
rect 588852 -3772 589088 -3536
rect 588532 -4092 588768 -3856
rect 588852 -4092 589088 -3856
rect 589492 669218 589728 669454
rect 589812 669218 590048 669454
rect 589492 668898 589728 669134
rect 589812 668898 590048 669134
rect 589492 633218 589728 633454
rect 589812 633218 590048 633454
rect 589492 632898 589728 633134
rect 589812 632898 590048 633134
rect 589492 597218 589728 597454
rect 589812 597218 590048 597454
rect 589492 596898 589728 597134
rect 589812 596898 590048 597134
rect 589492 561218 589728 561454
rect 589812 561218 590048 561454
rect 589492 560898 589728 561134
rect 589812 560898 590048 561134
rect 589492 525218 589728 525454
rect 589812 525218 590048 525454
rect 589492 524898 589728 525134
rect 589812 524898 590048 525134
rect 589492 489218 589728 489454
rect 589812 489218 590048 489454
rect 589492 488898 589728 489134
rect 589812 488898 590048 489134
rect 589492 453218 589728 453454
rect 589812 453218 590048 453454
rect 589492 452898 589728 453134
rect 589812 452898 590048 453134
rect 589492 417218 589728 417454
rect 589812 417218 590048 417454
rect 589492 416898 589728 417134
rect 589812 416898 590048 417134
rect 589492 381218 589728 381454
rect 589812 381218 590048 381454
rect 589492 380898 589728 381134
rect 589812 380898 590048 381134
rect 589492 345218 589728 345454
rect 589812 345218 590048 345454
rect 589492 344898 589728 345134
rect 589812 344898 590048 345134
rect 589492 309218 589728 309454
rect 589812 309218 590048 309454
rect 589492 308898 589728 309134
rect 589812 308898 590048 309134
rect 589492 273218 589728 273454
rect 589812 273218 590048 273454
rect 589492 272898 589728 273134
rect 589812 272898 590048 273134
rect 589492 237218 589728 237454
rect 589812 237218 590048 237454
rect 589492 236898 589728 237134
rect 589812 236898 590048 237134
rect 589492 201218 589728 201454
rect 589812 201218 590048 201454
rect 589492 200898 589728 201134
rect 589812 200898 590048 201134
rect 589492 165218 589728 165454
rect 589812 165218 590048 165454
rect 589492 164898 589728 165134
rect 589812 164898 590048 165134
rect 589492 129218 589728 129454
rect 589812 129218 590048 129454
rect 589492 128898 589728 129134
rect 589812 128898 590048 129134
rect 589492 93218 589728 93454
rect 589812 93218 590048 93454
rect 589492 92898 589728 93134
rect 589812 92898 590048 93134
rect 589492 57218 589728 57454
rect 589812 57218 590048 57454
rect 589492 56898 589728 57134
rect 589812 56898 590048 57134
rect 589492 21218 589728 21454
rect 589812 21218 590048 21454
rect 589492 20898 589728 21134
rect 589812 20898 590048 21134
rect 589492 -4732 589728 -4496
rect 589812 -4732 590048 -4496
rect 589492 -5052 589728 -4816
rect 589812 -5052 590048 -4816
rect 590452 673718 590688 673954
rect 590772 673718 591008 673954
rect 590452 673398 590688 673634
rect 590772 673398 591008 673634
rect 590452 637718 590688 637954
rect 590772 637718 591008 637954
rect 590452 637398 590688 637634
rect 590772 637398 591008 637634
rect 590452 601718 590688 601954
rect 590772 601718 591008 601954
rect 590452 601398 590688 601634
rect 590772 601398 591008 601634
rect 590452 565718 590688 565954
rect 590772 565718 591008 565954
rect 590452 565398 590688 565634
rect 590772 565398 591008 565634
rect 590452 529718 590688 529954
rect 590772 529718 591008 529954
rect 590452 529398 590688 529634
rect 590772 529398 591008 529634
rect 590452 493718 590688 493954
rect 590772 493718 591008 493954
rect 590452 493398 590688 493634
rect 590772 493398 591008 493634
rect 590452 457718 590688 457954
rect 590772 457718 591008 457954
rect 590452 457398 590688 457634
rect 590772 457398 591008 457634
rect 590452 421718 590688 421954
rect 590772 421718 591008 421954
rect 590452 421398 590688 421634
rect 590772 421398 591008 421634
rect 590452 385718 590688 385954
rect 590772 385718 591008 385954
rect 590452 385398 590688 385634
rect 590772 385398 591008 385634
rect 590452 349718 590688 349954
rect 590772 349718 591008 349954
rect 590452 349398 590688 349634
rect 590772 349398 591008 349634
rect 590452 313718 590688 313954
rect 590772 313718 591008 313954
rect 590452 313398 590688 313634
rect 590772 313398 591008 313634
rect 590452 277718 590688 277954
rect 590772 277718 591008 277954
rect 590452 277398 590688 277634
rect 590772 277398 591008 277634
rect 590452 241718 590688 241954
rect 590772 241718 591008 241954
rect 590452 241398 590688 241634
rect 590772 241398 591008 241634
rect 590452 205718 590688 205954
rect 590772 205718 591008 205954
rect 590452 205398 590688 205634
rect 590772 205398 591008 205634
rect 590452 169718 590688 169954
rect 590772 169718 591008 169954
rect 590452 169398 590688 169634
rect 590772 169398 591008 169634
rect 590452 133718 590688 133954
rect 590772 133718 591008 133954
rect 590452 133398 590688 133634
rect 590772 133398 591008 133634
rect 590452 97718 590688 97954
rect 590772 97718 591008 97954
rect 590452 97398 590688 97634
rect 590772 97398 591008 97634
rect 590452 61718 590688 61954
rect 590772 61718 591008 61954
rect 590452 61398 590688 61634
rect 590772 61398 591008 61634
rect 590452 25718 590688 25954
rect 590772 25718 591008 25954
rect 590452 25398 590688 25634
rect 590772 25398 591008 25634
rect 590452 -5692 590688 -5456
rect 590772 -5692 591008 -5456
rect 590452 -6012 590688 -5776
rect 590772 -6012 591008 -5776
rect 591412 678218 591648 678454
rect 591732 678218 591968 678454
rect 591412 677898 591648 678134
rect 591732 677898 591968 678134
rect 591412 642218 591648 642454
rect 591732 642218 591968 642454
rect 591412 641898 591648 642134
rect 591732 641898 591968 642134
rect 591412 606218 591648 606454
rect 591732 606218 591968 606454
rect 591412 605898 591648 606134
rect 591732 605898 591968 606134
rect 591412 570218 591648 570454
rect 591732 570218 591968 570454
rect 591412 569898 591648 570134
rect 591732 569898 591968 570134
rect 591412 534218 591648 534454
rect 591732 534218 591968 534454
rect 591412 533898 591648 534134
rect 591732 533898 591968 534134
rect 591412 498218 591648 498454
rect 591732 498218 591968 498454
rect 591412 497898 591648 498134
rect 591732 497898 591968 498134
rect 591412 462218 591648 462454
rect 591732 462218 591968 462454
rect 591412 461898 591648 462134
rect 591732 461898 591968 462134
rect 591412 426218 591648 426454
rect 591732 426218 591968 426454
rect 591412 425898 591648 426134
rect 591732 425898 591968 426134
rect 591412 390218 591648 390454
rect 591732 390218 591968 390454
rect 591412 389898 591648 390134
rect 591732 389898 591968 390134
rect 591412 354218 591648 354454
rect 591732 354218 591968 354454
rect 591412 353898 591648 354134
rect 591732 353898 591968 354134
rect 591412 318218 591648 318454
rect 591732 318218 591968 318454
rect 591412 317898 591648 318134
rect 591732 317898 591968 318134
rect 591412 282218 591648 282454
rect 591732 282218 591968 282454
rect 591412 281898 591648 282134
rect 591732 281898 591968 282134
rect 591412 246218 591648 246454
rect 591732 246218 591968 246454
rect 591412 245898 591648 246134
rect 591732 245898 591968 246134
rect 591412 210218 591648 210454
rect 591732 210218 591968 210454
rect 591412 209898 591648 210134
rect 591732 209898 591968 210134
rect 591412 174218 591648 174454
rect 591732 174218 591968 174454
rect 591412 173898 591648 174134
rect 591732 173898 591968 174134
rect 591412 138218 591648 138454
rect 591732 138218 591968 138454
rect 591412 137898 591648 138134
rect 591732 137898 591968 138134
rect 591412 102218 591648 102454
rect 591732 102218 591968 102454
rect 591412 101898 591648 102134
rect 591732 101898 591968 102134
rect 591412 66218 591648 66454
rect 591732 66218 591968 66454
rect 591412 65898 591648 66134
rect 591732 65898 591968 66134
rect 591412 30218 591648 30454
rect 591732 30218 591968 30454
rect 591412 29898 591648 30134
rect 591732 29898 591968 30134
rect 591412 -6652 591648 -6416
rect 591732 -6652 591968 -6416
rect 591412 -6972 591648 -6736
rect 591732 -6972 591968 -6736
rect 592372 682718 592608 682954
rect 592692 682718 592928 682954
rect 592372 682398 592608 682634
rect 592692 682398 592928 682634
rect 592372 646718 592608 646954
rect 592692 646718 592928 646954
rect 592372 646398 592608 646634
rect 592692 646398 592928 646634
rect 592372 610718 592608 610954
rect 592692 610718 592928 610954
rect 592372 610398 592608 610634
rect 592692 610398 592928 610634
rect 592372 574718 592608 574954
rect 592692 574718 592928 574954
rect 592372 574398 592608 574634
rect 592692 574398 592928 574634
rect 592372 538718 592608 538954
rect 592692 538718 592928 538954
rect 592372 538398 592608 538634
rect 592692 538398 592928 538634
rect 592372 502718 592608 502954
rect 592692 502718 592928 502954
rect 592372 502398 592608 502634
rect 592692 502398 592928 502634
rect 592372 466718 592608 466954
rect 592692 466718 592928 466954
rect 592372 466398 592608 466634
rect 592692 466398 592928 466634
rect 592372 430718 592608 430954
rect 592692 430718 592928 430954
rect 592372 430398 592608 430634
rect 592692 430398 592928 430634
rect 592372 394718 592608 394954
rect 592692 394718 592928 394954
rect 592372 394398 592608 394634
rect 592692 394398 592928 394634
rect 592372 358718 592608 358954
rect 592692 358718 592928 358954
rect 592372 358398 592608 358634
rect 592692 358398 592928 358634
rect 592372 322718 592608 322954
rect 592692 322718 592928 322954
rect 592372 322398 592608 322634
rect 592692 322398 592928 322634
rect 592372 286718 592608 286954
rect 592692 286718 592928 286954
rect 592372 286398 592608 286634
rect 592692 286398 592928 286634
rect 592372 250718 592608 250954
rect 592692 250718 592928 250954
rect 592372 250398 592608 250634
rect 592692 250398 592928 250634
rect 592372 214718 592608 214954
rect 592692 214718 592928 214954
rect 592372 214398 592608 214634
rect 592692 214398 592928 214634
rect 592372 178718 592608 178954
rect 592692 178718 592928 178954
rect 592372 178398 592608 178634
rect 592692 178398 592928 178634
rect 592372 142718 592608 142954
rect 592692 142718 592928 142954
rect 592372 142398 592608 142634
rect 592692 142398 592928 142634
rect 592372 106718 592608 106954
rect 592692 106718 592928 106954
rect 592372 106398 592608 106634
rect 592692 106398 592928 106634
rect 592372 70718 592608 70954
rect 592692 70718 592928 70954
rect 592372 70398 592608 70634
rect 592692 70398 592928 70634
rect 592372 34718 592608 34954
rect 592692 34718 592928 34954
rect 592372 34398 592608 34634
rect 592692 34398 592928 34634
rect 592372 -7612 592608 -7376
rect 592692 -7612 592928 -7376
rect 592372 -7932 592608 -7696
rect 592692 -7932 592928 -7696
<< metal5 >>
rect -9036 711868 592960 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect -9036 711548 592960 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect -9036 711280 592960 711312
rect -8076 710908 592000 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect -8076 710588 592000 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect -8076 710320 592000 710352
rect -7116 709948 591040 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect -7116 709628 591040 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect -7116 709360 591040 709392
rect -6156 708988 590080 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect -6156 708668 590080 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect -6156 708400 590080 708432
rect -5196 708028 589120 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect -5196 707708 589120 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect -5196 707440 589120 707472
rect -4236 707068 588160 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect -4236 706748 588160 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect -4236 706480 588160 706512
rect -3276 706108 587200 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect -3276 705788 587200 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect -3276 705520 587200 705552
rect -2316 705148 586240 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect -2316 704828 586240 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect -2316 704560 586240 704592
rect -9036 700954 592960 700986
rect -9036 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 592960 700954
rect -9036 700634 592960 700718
rect -9036 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 592960 700634
rect -9036 700366 592960 700398
rect -9036 696454 592960 696486
rect -9036 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 592960 696454
rect -9036 696134 592960 696218
rect -9036 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 592960 696134
rect -9036 695866 592960 695898
rect -9036 691954 592960 691986
rect -9036 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 592960 691954
rect -9036 691634 592960 691718
rect -9036 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 592960 691634
rect -9036 691366 592960 691398
rect -9036 687454 592960 687486
rect -9036 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 592960 687454
rect -9036 687134 592960 687218
rect -9036 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 592960 687134
rect -9036 686866 592960 686898
rect -9036 682954 592960 682986
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect -9036 682634 592960 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect -9036 682366 592960 682398
rect -9036 678454 592960 678486
rect -9036 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592960 678454
rect -9036 678134 592960 678218
rect -9036 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592960 678134
rect -9036 677866 592960 677898
rect -9036 673954 592960 673986
rect -9036 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 592960 673954
rect -9036 673634 592960 673718
rect -9036 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 592960 673634
rect -9036 673366 592960 673398
rect -9036 669454 592960 669486
rect -9036 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 592960 669454
rect -9036 669134 592960 669218
rect -9036 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 592960 669134
rect -9036 668866 592960 668898
rect -9036 664954 592960 664986
rect -9036 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 592960 664954
rect -9036 664634 592960 664718
rect -9036 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 592960 664634
rect -9036 664366 592960 664398
rect -9036 660454 592960 660486
rect -9036 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 592960 660454
rect -9036 660134 592960 660218
rect -9036 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 592960 660134
rect -9036 659866 592960 659898
rect -9036 655954 592960 655986
rect -9036 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 592960 655954
rect -9036 655634 592960 655718
rect -9036 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 592960 655634
rect -9036 655366 592960 655398
rect -9036 651454 592960 651486
rect -9036 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 592960 651454
rect -9036 651134 592960 651218
rect -9036 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 592960 651134
rect -9036 650866 592960 650898
rect -9036 646954 592960 646986
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect -9036 646634 592960 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect -9036 646366 592960 646398
rect -9036 642454 592960 642486
rect -9036 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592960 642454
rect -9036 642134 592960 642218
rect -9036 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592960 642134
rect -9036 641866 592960 641898
rect -9036 637954 592960 637986
rect -9036 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 592960 637954
rect -9036 637634 592960 637718
rect -9036 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 592960 637634
rect -9036 637366 592960 637398
rect -9036 633454 592960 633486
rect -9036 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 592960 633454
rect -9036 633134 592960 633218
rect -9036 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 592960 633134
rect -9036 632866 592960 632898
rect -9036 628954 592960 628986
rect -9036 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 592960 628954
rect -9036 628634 592960 628718
rect -9036 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 592960 628634
rect -9036 628366 592960 628398
rect -9036 624454 592960 624486
rect -9036 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 592960 624454
rect -9036 624134 592960 624218
rect -9036 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 592960 624134
rect -9036 623866 592960 623898
rect -9036 619954 592960 619986
rect -9036 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 592960 619954
rect -9036 619634 592960 619718
rect -9036 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 592960 619634
rect -9036 619366 592960 619398
rect -9036 615454 592960 615486
rect -9036 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 592960 615454
rect -9036 615134 592960 615218
rect -9036 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 592960 615134
rect -9036 614866 592960 614898
rect -9036 610954 592960 610986
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect -9036 610634 592960 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect -9036 610366 592960 610398
rect -9036 606454 592960 606486
rect -9036 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592960 606454
rect -9036 606134 592960 606218
rect -9036 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592960 606134
rect -9036 605866 592960 605898
rect -9036 601954 592960 601986
rect -9036 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 592960 601954
rect -9036 601634 592960 601718
rect -9036 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 592960 601634
rect -9036 601366 592960 601398
rect -9036 597454 592960 597486
rect -9036 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 592960 597454
rect -9036 597134 592960 597218
rect -9036 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 592960 597134
rect -9036 596866 592960 596898
rect -9036 592954 592960 592986
rect -9036 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 592960 592954
rect -9036 592634 592960 592718
rect -9036 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 592960 592634
rect -9036 592366 592960 592398
rect -9036 588454 592960 588486
rect -9036 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 592960 588454
rect -9036 588134 592960 588218
rect -9036 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 592960 588134
rect -9036 587866 592960 587898
rect -9036 583954 592960 583986
rect -9036 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 592960 583954
rect -9036 583634 592960 583718
rect -9036 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 592960 583634
rect -9036 583366 592960 583398
rect -9036 579454 592960 579486
rect -9036 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 592960 579454
rect -9036 579134 592960 579218
rect -9036 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 592960 579134
rect -9036 578866 592960 578898
rect -9036 574954 592960 574986
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect -9036 574634 592960 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect -9036 574366 592960 574398
rect -9036 570454 592960 570486
rect -9036 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592960 570454
rect -9036 570134 592960 570218
rect -9036 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592960 570134
rect -9036 569866 592960 569898
rect -9036 565954 592960 565986
rect -9036 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 592960 565954
rect -9036 565634 592960 565718
rect -9036 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 592960 565634
rect -9036 565366 592960 565398
rect -9036 561454 592960 561486
rect -9036 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 592960 561454
rect -9036 561134 592960 561218
rect -9036 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 592960 561134
rect -9036 560866 592960 560898
rect -9036 556954 592960 556986
rect -9036 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 592960 556954
rect -9036 556634 592960 556718
rect -9036 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 592960 556634
rect -9036 556366 592960 556398
rect -9036 552454 592960 552486
rect -9036 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 592960 552454
rect -9036 552134 592960 552218
rect -9036 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 592960 552134
rect -9036 551866 592960 551898
rect -9036 547954 592960 547986
rect -9036 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 592960 547954
rect -9036 547634 592960 547718
rect -9036 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 592960 547634
rect -9036 547366 592960 547398
rect -9036 543454 592960 543486
rect -9036 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 592960 543454
rect -9036 543134 592960 543218
rect -9036 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 592960 543134
rect -9036 542866 592960 542898
rect -9036 538954 592960 538986
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect -9036 538634 592960 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect -9036 538366 592960 538398
rect -9036 534454 592960 534486
rect -9036 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592960 534454
rect -9036 534134 592960 534218
rect -9036 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592960 534134
rect -9036 533866 592960 533898
rect -9036 529954 592960 529986
rect -9036 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 592960 529954
rect -9036 529634 592960 529718
rect -9036 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 592960 529634
rect -9036 529366 592960 529398
rect -9036 525454 592960 525486
rect -9036 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 592960 525454
rect -9036 525134 592960 525218
rect -9036 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 592960 525134
rect -9036 524866 592960 524898
rect -9036 520954 592960 520986
rect -9036 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 592960 520954
rect -9036 520634 592960 520718
rect -9036 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 592960 520634
rect -9036 520366 592960 520398
rect -9036 516454 592960 516486
rect -9036 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 592960 516454
rect -9036 516134 592960 516218
rect -9036 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 592960 516134
rect -9036 515866 592960 515898
rect -9036 511954 592960 511986
rect -9036 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 592960 511954
rect -9036 511634 592960 511718
rect -9036 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 592960 511634
rect -9036 511366 592960 511398
rect -9036 507454 592960 507486
rect -9036 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 592960 507454
rect -9036 507134 592960 507218
rect -9036 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 592960 507134
rect -9036 506866 592960 506898
rect -9036 502954 592960 502986
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect -9036 502634 592960 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect -9036 502366 592960 502398
rect -9036 498454 592960 498486
rect -9036 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592960 498454
rect -9036 498134 592960 498218
rect -9036 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592960 498134
rect -9036 497866 592960 497898
rect -9036 493954 592960 493986
rect -9036 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 592960 493954
rect -9036 493634 592960 493718
rect -9036 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 592960 493634
rect -9036 493366 592960 493398
rect -9036 489454 592960 489486
rect -9036 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 592960 489454
rect -9036 489134 592960 489218
rect -9036 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 592960 489134
rect -9036 488866 592960 488898
rect -9036 484954 592960 484986
rect -9036 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 592960 484954
rect -9036 484634 592960 484718
rect -9036 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 592960 484634
rect -9036 484366 592960 484398
rect -9036 480454 592960 480486
rect -9036 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 592960 480454
rect -9036 480134 592960 480218
rect -9036 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 592960 480134
rect -9036 479866 592960 479898
rect -9036 475954 592960 475986
rect -9036 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 592960 475954
rect -9036 475634 592960 475718
rect -9036 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 592960 475634
rect -9036 475366 592960 475398
rect -9036 471454 592960 471486
rect -9036 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 592960 471454
rect -9036 471134 592960 471218
rect -9036 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 592960 471134
rect -9036 470866 592960 470898
rect -9036 466954 592960 466986
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect -9036 466634 592960 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect -9036 466366 592960 466398
rect -9036 462454 592960 462486
rect -9036 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592960 462454
rect -9036 462134 592960 462218
rect -9036 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592960 462134
rect -9036 461866 592960 461898
rect -9036 457954 592960 457986
rect -9036 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 592960 457954
rect -9036 457634 592960 457718
rect -9036 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 592960 457634
rect -9036 457366 592960 457398
rect -9036 453454 592960 453486
rect -9036 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 592960 453454
rect -9036 453134 592960 453218
rect -9036 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 592960 453134
rect -9036 452866 592960 452898
rect -9036 448954 592960 448986
rect -9036 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 592960 448954
rect -9036 448634 592960 448718
rect -9036 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 592960 448634
rect -9036 448366 592960 448398
rect -9036 444454 592960 444486
rect -9036 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 592960 444454
rect -9036 444134 592960 444218
rect -9036 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 592960 444134
rect -9036 443866 592960 443898
rect -9036 439954 592960 439986
rect -9036 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 592960 439954
rect -9036 439634 592960 439718
rect -9036 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 592960 439634
rect -9036 439366 592960 439398
rect -9036 435454 592960 435486
rect -9036 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 236650 435454
rect 236886 435218 267370 435454
rect 267606 435218 298090 435454
rect 298326 435218 328810 435454
rect 329046 435218 359530 435454
rect 359766 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 592960 435454
rect -9036 435134 592960 435218
rect -9036 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 236650 435134
rect 236886 434898 267370 435134
rect 267606 434898 298090 435134
rect 298326 434898 328810 435134
rect 329046 434898 359530 435134
rect 359766 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 592960 435134
rect -9036 434866 592960 434898
rect -9036 430954 592960 430986
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect -9036 430634 592960 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect -9036 430366 592960 430398
rect -9036 426454 592960 426486
rect -9036 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592960 426454
rect -9036 426134 592960 426218
rect -9036 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592960 426134
rect -9036 425866 592960 425898
rect -9036 421954 592960 421986
rect -9036 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 592960 421954
rect -9036 421634 592960 421718
rect -9036 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 592960 421634
rect -9036 421366 592960 421398
rect -9036 417454 592960 417486
rect -9036 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 592960 417454
rect -9036 417134 592960 417218
rect -9036 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 592960 417134
rect -9036 416866 592960 416898
rect -9036 412954 592960 412986
rect -9036 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 592960 412954
rect -9036 412634 592960 412718
rect -9036 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 592960 412634
rect -9036 412366 592960 412398
rect -9036 408454 592960 408486
rect -9036 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 592960 408454
rect -9036 408134 592960 408218
rect -9036 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 592960 408134
rect -9036 407866 592960 407898
rect -9036 403954 592960 403986
rect -9036 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 252010 403954
rect 252246 403718 282730 403954
rect 282966 403718 313450 403954
rect 313686 403718 344170 403954
rect 344406 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 592960 403954
rect -9036 403634 592960 403718
rect -9036 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 252010 403634
rect 252246 403398 282730 403634
rect 282966 403398 313450 403634
rect 313686 403398 344170 403634
rect 344406 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 592960 403634
rect -9036 403366 592960 403398
rect -9036 399454 592960 399486
rect -9036 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 236650 399454
rect 236886 399218 267370 399454
rect 267606 399218 298090 399454
rect 298326 399218 328810 399454
rect 329046 399218 359530 399454
rect 359766 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 592960 399454
rect -9036 399134 592960 399218
rect -9036 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 236650 399134
rect 236886 398898 267370 399134
rect 267606 398898 298090 399134
rect 298326 398898 328810 399134
rect 329046 398898 359530 399134
rect 359766 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 592960 399134
rect -9036 398866 592960 398898
rect -9036 394954 592960 394986
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect -9036 394634 592960 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect -9036 394366 592960 394398
rect -9036 390454 592960 390486
rect -9036 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592960 390454
rect -9036 390134 592960 390218
rect -9036 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592960 390134
rect -9036 389866 592960 389898
rect -9036 385954 592960 385986
rect -9036 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 592960 385954
rect -9036 385634 592960 385718
rect -9036 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 592960 385634
rect -9036 385366 592960 385398
rect -9036 381454 592960 381486
rect -9036 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 592960 381454
rect -9036 381134 592960 381218
rect -9036 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 592960 381134
rect -9036 380866 592960 380898
rect -9036 376954 592960 376986
rect -9036 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 592960 376954
rect -9036 376634 592960 376718
rect -9036 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 592960 376634
rect -9036 376366 592960 376398
rect -9036 372454 592960 372486
rect -9036 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 592960 372454
rect -9036 372134 592960 372218
rect -9036 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 592960 372134
rect -9036 371866 592960 371898
rect -9036 367954 592960 367986
rect -9036 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 119610 367954
rect 119846 367718 150330 367954
rect 150566 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 252010 367954
rect 252246 367718 282730 367954
rect 282966 367718 313450 367954
rect 313686 367718 344170 367954
rect 344406 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 592960 367954
rect -9036 367634 592960 367718
rect -9036 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 119610 367634
rect 119846 367398 150330 367634
rect 150566 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 252010 367634
rect 252246 367398 282730 367634
rect 282966 367398 313450 367634
rect 313686 367398 344170 367634
rect 344406 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 592960 367634
rect -9036 367366 592960 367398
rect -9036 363454 592960 363486
rect -9036 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 104250 363454
rect 104486 363218 134970 363454
rect 135206 363218 165690 363454
rect 165926 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 236650 363454
rect 236886 363218 267370 363454
rect 267606 363218 298090 363454
rect 298326 363218 328810 363454
rect 329046 363218 359530 363454
rect 359766 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 592960 363454
rect -9036 363134 592960 363218
rect -9036 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 104250 363134
rect 104486 362898 134970 363134
rect 135206 362898 165690 363134
rect 165926 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 236650 363134
rect 236886 362898 267370 363134
rect 267606 362898 298090 363134
rect 298326 362898 328810 363134
rect 329046 362898 359530 363134
rect 359766 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 592960 363134
rect -9036 362866 592960 362898
rect -9036 358954 592960 358986
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect -9036 358634 592960 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect -9036 358366 592960 358398
rect -9036 354454 592960 354486
rect -9036 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592960 354454
rect -9036 354134 592960 354218
rect -9036 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592960 354134
rect -9036 353866 592960 353898
rect -9036 349954 592960 349986
rect -9036 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 592960 349954
rect -9036 349634 592960 349718
rect -9036 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 592960 349634
rect -9036 349366 592960 349398
rect -9036 345454 592960 345486
rect -9036 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 592960 345454
rect -9036 345134 592960 345218
rect -9036 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 592960 345134
rect -9036 344866 592960 344898
rect -9036 340954 592960 340986
rect -9036 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 592960 340954
rect -9036 340634 592960 340718
rect -9036 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 592960 340634
rect -9036 340366 592960 340398
rect -9036 336454 592960 336486
rect -9036 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 592960 336454
rect -9036 336134 592960 336218
rect -9036 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 592960 336134
rect -9036 335866 592960 335898
rect -9036 331954 592960 331986
rect -9036 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 119610 331954
rect 119846 331718 150330 331954
rect 150566 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 252010 331954
rect 252246 331718 282730 331954
rect 282966 331718 313450 331954
rect 313686 331718 344170 331954
rect 344406 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 592960 331954
rect -9036 331634 592960 331718
rect -9036 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 119610 331634
rect 119846 331398 150330 331634
rect 150566 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 252010 331634
rect 252246 331398 282730 331634
rect 282966 331398 313450 331634
rect 313686 331398 344170 331634
rect 344406 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 592960 331634
rect -9036 331366 592960 331398
rect -9036 327454 592960 327486
rect -9036 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 104250 327454
rect 104486 327218 134970 327454
rect 135206 327218 165690 327454
rect 165926 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 236650 327454
rect 236886 327218 267370 327454
rect 267606 327218 298090 327454
rect 298326 327218 328810 327454
rect 329046 327218 359530 327454
rect 359766 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 592960 327454
rect -9036 327134 592960 327218
rect -9036 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 104250 327134
rect 104486 326898 134970 327134
rect 135206 326898 165690 327134
rect 165926 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 236650 327134
rect 236886 326898 267370 327134
rect 267606 326898 298090 327134
rect 298326 326898 328810 327134
rect 329046 326898 359530 327134
rect 359766 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 592960 327134
rect -9036 326866 592960 326898
rect -9036 322954 592960 322986
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect -9036 322634 592960 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect -9036 322366 592960 322398
rect -9036 318454 592960 318486
rect -9036 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592960 318454
rect -9036 318134 592960 318218
rect -9036 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592960 318134
rect -9036 317866 592960 317898
rect -9036 313954 592960 313986
rect -9036 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 592960 313954
rect -9036 313634 592960 313718
rect -9036 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 592960 313634
rect -9036 313366 592960 313398
rect -9036 309454 592960 309486
rect -9036 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 592960 309454
rect -9036 309134 592960 309218
rect -9036 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 592960 309134
rect -9036 308866 592960 308898
rect -9036 304954 592960 304986
rect -9036 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 592960 304954
rect -9036 304634 592960 304718
rect -9036 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 592960 304634
rect -9036 304366 592960 304398
rect -9036 300454 592960 300486
rect -9036 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 592960 300454
rect -9036 300134 592960 300218
rect -9036 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 592960 300134
rect -9036 299866 592960 299898
rect -9036 295954 592960 295986
rect -9036 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 592960 295954
rect -9036 295634 592960 295718
rect -9036 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 592960 295634
rect -9036 295366 592960 295398
rect -9036 291454 592960 291486
rect -9036 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 592960 291454
rect -9036 291134 592960 291218
rect -9036 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 592960 291134
rect -9036 290866 592960 290898
rect -9036 286954 592960 286986
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect -9036 286634 592960 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect -9036 286366 592960 286398
rect -9036 282454 592960 282486
rect -9036 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592960 282454
rect -9036 282134 592960 282218
rect -9036 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592960 282134
rect -9036 281866 592960 281898
rect -9036 277954 592960 277986
rect -9036 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 592960 277954
rect -9036 277634 592960 277718
rect -9036 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 592960 277634
rect -9036 277366 592960 277398
rect -9036 273454 592960 273486
rect -9036 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 592960 273454
rect -9036 273134 592960 273218
rect -9036 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 592960 273134
rect -9036 272866 592960 272898
rect -9036 268954 592960 268986
rect -9036 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 592960 268954
rect -9036 268634 592960 268718
rect -9036 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 592960 268634
rect -9036 268366 592960 268398
rect -9036 264454 592960 264486
rect -9036 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 592960 264454
rect -9036 264134 592960 264218
rect -9036 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 592960 264134
rect -9036 263866 592960 263898
rect -9036 259954 592960 259986
rect -9036 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 592960 259954
rect -9036 259634 592960 259718
rect -9036 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 592960 259634
rect -9036 259366 592960 259398
rect -9036 255454 592960 255486
rect -9036 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 592960 255454
rect -9036 255134 592960 255218
rect -9036 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 592960 255134
rect -9036 254866 592960 254898
rect -9036 250954 592960 250986
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect -9036 250634 592960 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect -9036 250366 592960 250398
rect -9036 246454 592960 246486
rect -9036 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592960 246454
rect -9036 246134 592960 246218
rect -9036 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592960 246134
rect -9036 245866 592960 245898
rect -9036 241954 592960 241986
rect -9036 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 592960 241954
rect -9036 241634 592960 241718
rect -9036 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 592960 241634
rect -9036 241366 592960 241398
rect -9036 237454 592960 237486
rect -9036 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 592960 237454
rect -9036 237134 592960 237218
rect -9036 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 592960 237134
rect -9036 236866 592960 236898
rect -9036 232954 592960 232986
rect -9036 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 592960 232954
rect -9036 232634 592960 232718
rect -9036 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 592960 232634
rect -9036 232366 592960 232398
rect -9036 228454 592960 228486
rect -9036 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 592960 228454
rect -9036 228134 592960 228218
rect -9036 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 592960 228134
rect -9036 227866 592960 227898
rect -9036 223954 592960 223986
rect -9036 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 220328 223954
rect 220564 223718 356056 223954
rect 356292 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 592960 223954
rect -9036 223634 592960 223718
rect -9036 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 220328 223634
rect 220564 223398 356056 223634
rect 356292 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 592960 223634
rect -9036 223366 592960 223398
rect -9036 219454 592960 219486
rect -9036 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 592960 219454
rect -9036 219134 592960 219218
rect -9036 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 592960 219134
rect -9036 218866 592960 218898
rect -9036 214954 592960 214986
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect -9036 214634 592960 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect -9036 214366 592960 214398
rect -9036 210454 592960 210486
rect -9036 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592960 210454
rect -9036 210134 592960 210218
rect -9036 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592960 210134
rect -9036 209866 592960 209898
rect -9036 205954 592960 205986
rect -9036 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 592960 205954
rect -9036 205634 592960 205718
rect -9036 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 592960 205634
rect -9036 205366 592960 205398
rect -9036 201454 592960 201486
rect -9036 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 592960 201454
rect -9036 201134 592960 201218
rect -9036 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 592960 201134
rect -9036 200866 592960 200898
rect -9036 196954 592960 196986
rect -9036 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 592960 196954
rect -9036 196634 592960 196718
rect -9036 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 592960 196634
rect -9036 196366 592960 196398
rect -9036 192454 592960 192486
rect -9036 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 592960 192454
rect -9036 192134 592960 192218
rect -9036 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 592960 192134
rect -9036 191866 592960 191898
rect -9036 187954 592960 187986
rect -9036 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 220328 187954
rect 220564 187718 356056 187954
rect 356292 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 592960 187954
rect -9036 187634 592960 187718
rect -9036 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 220328 187634
rect 220564 187398 356056 187634
rect 356292 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 592960 187634
rect -9036 187366 592960 187398
rect -9036 183454 592960 183486
rect -9036 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 592960 183454
rect -9036 183134 592960 183218
rect -9036 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 592960 183134
rect -9036 182866 592960 182898
rect -9036 178954 592960 178986
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect -9036 178634 592960 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect -9036 178366 592960 178398
rect -9036 174454 592960 174486
rect -9036 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592960 174454
rect -9036 174134 592960 174218
rect -9036 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592960 174134
rect -9036 173866 592960 173898
rect -9036 169954 592960 169986
rect -9036 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 592960 169954
rect -9036 169634 592960 169718
rect -9036 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 592960 169634
rect -9036 169366 592960 169398
rect -9036 165454 592960 165486
rect -9036 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 592960 165454
rect -9036 165134 592960 165218
rect -9036 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 592960 165134
rect -9036 164866 592960 164898
rect -9036 160954 592960 160986
rect -9036 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 592960 160954
rect -9036 160634 592960 160718
rect -9036 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 592960 160634
rect -9036 160366 592960 160398
rect -9036 156454 592960 156486
rect -9036 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 592960 156454
rect -9036 156134 592960 156218
rect -9036 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 592960 156134
rect -9036 155866 592960 155898
rect -9036 151954 592960 151986
rect -9036 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 592960 151954
rect -9036 151634 592960 151718
rect -9036 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 592960 151634
rect -9036 151366 592960 151398
rect -9036 147454 592960 147486
rect -9036 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 592960 147454
rect -9036 147134 592960 147218
rect -9036 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 592960 147134
rect -9036 146866 592960 146898
rect -9036 142954 592960 142986
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect -9036 142634 592960 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect -9036 142366 592960 142398
rect -9036 138454 592960 138486
rect -9036 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592960 138454
rect -9036 138134 592960 138218
rect -9036 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592960 138134
rect -9036 137866 592960 137898
rect -9036 133954 592960 133986
rect -9036 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 592960 133954
rect -9036 133634 592960 133718
rect -9036 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 592960 133634
rect -9036 133366 592960 133398
rect -9036 129454 592960 129486
rect -9036 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 592960 129454
rect -9036 129134 592960 129218
rect -9036 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 592960 129134
rect -9036 128866 592960 128898
rect -9036 124954 592960 124986
rect -9036 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 592960 124954
rect -9036 124634 592960 124718
rect -9036 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 592960 124634
rect -9036 124366 592960 124398
rect -9036 120454 592960 120486
rect -9036 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 592960 120454
rect -9036 120134 592960 120218
rect -9036 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 592960 120134
rect -9036 119866 592960 119898
rect -9036 115954 592960 115986
rect -9036 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 592960 115954
rect -9036 115634 592960 115718
rect -9036 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 592960 115634
rect -9036 115366 592960 115398
rect -9036 111454 592960 111486
rect -9036 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 592960 111454
rect -9036 111134 592960 111218
rect -9036 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 592960 111134
rect -9036 110866 592960 110898
rect -9036 106954 592960 106986
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect -9036 106634 592960 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect -9036 106366 592960 106398
rect -9036 102454 592960 102486
rect -9036 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592960 102454
rect -9036 102134 592960 102218
rect -9036 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592960 102134
rect -9036 101866 592960 101898
rect -9036 97954 592960 97986
rect -9036 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 592960 97954
rect -9036 97634 592960 97718
rect -9036 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 592960 97634
rect -9036 97366 592960 97398
rect -9036 93454 592960 93486
rect -9036 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 592960 93454
rect -9036 93134 592960 93218
rect -9036 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 592960 93134
rect -9036 92866 592960 92898
rect -9036 88954 592960 88986
rect -9036 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 592960 88954
rect -9036 88634 592960 88718
rect -9036 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 592960 88634
rect -9036 88366 592960 88398
rect -9036 84454 592960 84486
rect -9036 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 592960 84454
rect -9036 84134 592960 84218
rect -9036 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 592960 84134
rect -9036 83866 592960 83898
rect -9036 79954 592960 79986
rect -9036 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 592960 79954
rect -9036 79634 592960 79718
rect -9036 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 592960 79634
rect -9036 79366 592960 79398
rect -9036 75454 592960 75486
rect -9036 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 592960 75454
rect -9036 75134 592960 75218
rect -9036 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 592960 75134
rect -9036 74866 592960 74898
rect -9036 70954 592960 70986
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect -9036 70634 592960 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect -9036 70366 592960 70398
rect -9036 66454 592960 66486
rect -9036 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592960 66454
rect -9036 66134 592960 66218
rect -9036 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592960 66134
rect -9036 65866 592960 65898
rect -9036 61954 592960 61986
rect -9036 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 592960 61954
rect -9036 61634 592960 61718
rect -9036 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 592960 61634
rect -9036 61366 592960 61398
rect -9036 57454 592960 57486
rect -9036 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 592960 57454
rect -9036 57134 592960 57218
rect -9036 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 592960 57134
rect -9036 56866 592960 56898
rect -9036 52954 592960 52986
rect -9036 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 592960 52954
rect -9036 52634 592960 52718
rect -9036 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 592960 52634
rect -9036 52366 592960 52398
rect -9036 48454 592960 48486
rect -9036 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 592960 48454
rect -9036 48134 592960 48218
rect -9036 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 592960 48134
rect -9036 47866 592960 47898
rect -9036 43954 592960 43986
rect -9036 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 592960 43954
rect -9036 43634 592960 43718
rect -9036 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 592960 43634
rect -9036 43366 592960 43398
rect -9036 39454 592960 39486
rect -9036 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 592960 39454
rect -9036 39134 592960 39218
rect -9036 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 592960 39134
rect -9036 38866 592960 38898
rect -9036 34954 592960 34986
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect -9036 34634 592960 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect -9036 34366 592960 34398
rect -9036 30454 592960 30486
rect -9036 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592960 30454
rect -9036 30134 592960 30218
rect -9036 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592960 30134
rect -9036 29866 592960 29898
rect -9036 25954 592960 25986
rect -9036 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 592960 25954
rect -9036 25634 592960 25718
rect -9036 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 592960 25634
rect -9036 25366 592960 25398
rect -9036 21454 592960 21486
rect -9036 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 592960 21454
rect -9036 21134 592960 21218
rect -9036 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 592960 21134
rect -9036 20866 592960 20898
rect -9036 16954 592960 16986
rect -9036 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 592960 16954
rect -9036 16634 592960 16718
rect -9036 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 592960 16634
rect -9036 16366 592960 16398
rect -9036 12454 592960 12486
rect -9036 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 592960 12454
rect -9036 12134 592960 12218
rect -9036 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 592960 12134
rect -9036 11866 592960 11898
rect -9036 7954 592960 7986
rect -9036 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 592960 7954
rect -9036 7634 592960 7718
rect -9036 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 592960 7634
rect -9036 7366 592960 7398
rect -9036 3454 592960 3486
rect -9036 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 592960 3454
rect -9036 3134 592960 3218
rect -9036 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 592960 3134
rect -9036 2866 592960 2898
rect -2316 -656 586240 -624
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect -2316 -976 586240 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect -2316 -1244 586240 -1212
rect -3276 -1616 587200 -1584
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect -3276 -1936 587200 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect -3276 -2204 587200 -2172
rect -4236 -2576 588160 -2544
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect -4236 -2896 588160 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect -4236 -3164 588160 -3132
rect -5196 -3536 589120 -3504
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect -5196 -3856 589120 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect -5196 -4124 589120 -4092
rect -6156 -4496 590080 -4464
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect -6156 -4816 590080 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect -6156 -5084 590080 -5052
rect -7116 -5456 591040 -5424
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect -7116 -5776 591040 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect -7116 -6044 591040 -6012
rect -8076 -6416 592000 -6384
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect -8076 -6736 592000 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect -8076 -7004 592000 -6972
rect -9036 -7376 592960 -7344
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect -9036 -7696 592960 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect -9036 -7964 592960 -7932
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst
timestamp 0
transform 1 0 220000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 232400 0 1 310400
box 13 0 128970 131144
use wbuart_wrap  uart_inst
timestamp 0
transform 1 0 100000 0 1 300000
box 0 0 70020 72164
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2316 -1244 -1696 705180 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 -1244 586240 -624 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 704560 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585620 -1244 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7964 2414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7964 38414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7964 74414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7964 110414 298000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 374164 110414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7964 146414 298000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 374164 146414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7964 182414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7964 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7964 254414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 245308 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7964 290414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 245308 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7964 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7964 362414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 443544 362414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7964 398414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7964 434414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7964 470414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7964 506414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7964 542414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7964 578414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 2866 592960 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 38866 592960 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 74866 592960 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 110866 592960 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 146866 592960 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 182866 592960 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 218866 592960 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 254866 592960 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 290866 592960 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 326866 592960 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 362866 592960 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 398866 592960 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 434866 592960 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 470866 592960 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 506866 592960 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 542866 592960 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 578866 592960 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 614866 592960 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 650866 592960 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 686866 592960 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -4236 -3164 -3616 707100 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 -3164 588160 -2544 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 706480 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587540 -3164 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7964 11414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7964 47414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7964 83414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7964 119414 298000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 374164 119414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7964 155414 298000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 374164 155414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7964 191414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7964 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7964 263414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 245308 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7964 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7964 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7964 371414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7964 407414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7964 443414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7964 479414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7964 515414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7964 551414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 11866 592960 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 47866 592960 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 83866 592960 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 119866 592960 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 155866 592960 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 191866 592960 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 227866 592960 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 263866 592960 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 299866 592960 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 335866 592960 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 371866 592960 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 407866 592960 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 443866 592960 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 479866 592960 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 515866 592960 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 551866 592960 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 587866 592960 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 623866 592960 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 659866 592960 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 695866 592960 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5196 -4124 -4576 708060 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 -4124 589120 -3504 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 707440 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 588500 -4124 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 15294 -7964 15914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 51294 -7964 51914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 87294 -7964 87914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 -7964 123914 298000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 374164 123914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 -7964 159914 298000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 374164 159914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 195294 -7964 195914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 -7964 231914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 565308 231914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 -7964 267914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 245308 267914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 565308 267914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 -7964 303914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 565308 303914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 -7964 339914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 565308 339914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 375294 -7964 375914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 411294 -7964 411914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 447294 -7964 447914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 483294 -7964 483914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 519294 -7964 519914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 555294 -7964 555914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 16366 592960 16986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 52366 592960 52986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 88366 592960 88986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 124366 592960 124986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 160366 592960 160986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 196366 592960 196986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 232366 592960 232986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 268366 592960 268986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 304366 592960 304986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 340366 592960 340986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 376366 592960 376986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 412366 592960 412986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 448366 592960 448986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 484366 592960 484986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 520366 592960 520986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 556366 592960 556986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 592366 592960 592986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 628366 592960 628986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 664366 592960 664986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 700366 592960 700986 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -6156 -5084 -5536 709020 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 -5084 590080 -4464 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 708400 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 589460 -5084 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 19794 -7964 20414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 55794 -7964 56414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 91794 -7964 92414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 -7964 128414 298000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 374164 128414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 -7964 164414 298000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 374164 164414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 199794 -7964 200414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 -7964 236414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 -7964 272414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 -7964 308414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 -7964 344414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 379794 -7964 380414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 415794 -7964 416414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 451794 -7964 452414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 487794 -7964 488414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 523794 -7964 524414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 559794 -7964 560414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 20866 592960 21486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 56866 592960 57486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 92866 592960 93486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 128866 592960 129486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 164866 592960 165486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 200866 592960 201486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 236866 592960 237486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 272866 592960 273486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 308866 592960 309486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 344866 592960 345486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 380866 592960 381486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 416866 592960 417486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 452866 592960 453486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 488866 592960 489486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 524866 592960 525486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 560866 592960 561486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 596866 592960 597486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 632866 592960 633486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 668866 592960 669486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -8076 -7004 -7456 710940 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 -7004 592000 -6384 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 710320 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 591380 -7004 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 28794 -7964 29414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 64794 -7964 65414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 -7964 101414 298000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 374164 101414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 -7964 137414 298000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 374164 137414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 172794 -7964 173414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 208794 -7964 209414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 -7964 245414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 245308 245414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 565308 245414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 -7964 281414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 245308 281414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 565308 281414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 -7964 317414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 565308 317414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 -7964 353414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 565308 353414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 388794 -7964 389414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 424794 -7964 425414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 460794 -7964 461414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 496794 -7964 497414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 532794 -7964 533414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 568794 -7964 569414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 29866 592960 30486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 65866 592960 66486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 101866 592960 102486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 137866 592960 138486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 173866 592960 174486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 209866 592960 210486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 245866 592960 246486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 281866 592960 282486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 317866 592960 318486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 353866 592960 354486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 389866 592960 390486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 425866 592960 426486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 461866 592960 462486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 497866 592960 498486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 533866 592960 534486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 569866 592960 570486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 605866 592960 606486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 641866 592960 642486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 677866 592960 678486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -9036 -7964 -8416 711900 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 -7964 592960 -7344 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 711280 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592340 -7964 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7964 33914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7964 69914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7964 105914 298000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 374164 105914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7964 141914 298000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 374164 141914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7964 177914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7964 213914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7964 249914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 245308 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7964 285914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 245308 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7964 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7964 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7964 393914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7964 429914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7964 465914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7964 501914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7964 537914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7964 573914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 34366 592960 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 70366 592960 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 106366 592960 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 142366 592960 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 178366 592960 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 214366 592960 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 250366 592960 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 286366 592960 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 322366 592960 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 358366 592960 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 394366 592960 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 430366 592960 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 466366 592960 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 502366 592960 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 538366 592960 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 574366 592960 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 610366 592960 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 646366 592960 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 682366 592960 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -3276 -2204 -2656 706140 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 -2204 587200 -1584 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 705520 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586580 -2204 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7964 6914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7964 42914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7964 78914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7964 114914 298000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 374164 114914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7964 150914 298000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 374164 150914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7964 186914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7964 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7964 258914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 245308 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7964 294914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 245308 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7964 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7964 366914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7964 402914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7964 438914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7964 474914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7964 510914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7964 546914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7964 582914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 7366 592960 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 43366 592960 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 79366 592960 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 115366 592960 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 151366 592960 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 187366 592960 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 223366 592960 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 259366 592960 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 295366 592960 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 331366 592960 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 367366 592960 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 403366 592960 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 439366 592960 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 475366 592960 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 511366 592960 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 547366 592960 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 583366 592960 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 619366 592960 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 655366 592960 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 691366 592960 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -7116 -6044 -6496 709980 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 -6044 591040 -5424 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 709360 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 590420 -6044 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 24294 -7964 24914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 60294 -7964 60914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 96294 -7964 96914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 -7964 132914 298000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 374164 132914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 -7964 168914 298000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 374164 168914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 204294 -7964 204914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 -7964 240914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 -7964 276914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 -7964 312914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 -7964 348914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 384294 -7964 384914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 420294 -7964 420914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 456294 -7964 456914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 492294 -7964 492914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 528294 -7964 528914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 564294 -7964 564914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 25366 592960 25986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 61366 592960 61986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 97366 592960 97986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 133366 592960 133986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 169366 592960 169986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 205366 592960 205986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 241366 592960 241986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 277366 592960 277986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 313366 592960 313986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 349366 592960 349986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 385366 592960 385986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 421366 592960 421986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 457366 592960 457986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 493366 592960 493986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 529366 592960 529986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 565366 592960 565986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 601366 592960 601986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 637366 592960 637986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 673366 592960 673986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
