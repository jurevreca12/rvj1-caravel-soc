magic
tech sky130A
magscale 1 2
timestamp 1654606238
<< obsli1 >>
rect 1104 2159 130364 131121
<< obsm1 >>
rect 14 348 131362 131640
<< metal2 >>
rect 386 132826 442 133626
rect 1122 132826 1178 133626
rect 1858 132826 1914 133626
rect 2686 132826 2742 133626
rect 3422 132826 3478 133626
rect 4250 132826 4306 133626
rect 4986 132826 5042 133626
rect 5814 132826 5870 133626
rect 6550 132826 6606 133626
rect 7378 132826 7434 133626
rect 8114 132826 8170 133626
rect 8942 132826 8998 133626
rect 9678 132826 9734 133626
rect 10414 132826 10470 133626
rect 11242 132826 11298 133626
rect 11978 132826 12034 133626
rect 12806 132826 12862 133626
rect 13542 132826 13598 133626
rect 14370 132826 14426 133626
rect 15106 132826 15162 133626
rect 15934 132826 15990 133626
rect 16670 132826 16726 133626
rect 17498 132826 17554 133626
rect 18234 132826 18290 133626
rect 18970 132826 19026 133626
rect 19798 132826 19854 133626
rect 20534 132826 20590 133626
rect 21362 132826 21418 133626
rect 22098 132826 22154 133626
rect 22926 132826 22982 133626
rect 23662 132826 23718 133626
rect 24490 132826 24546 133626
rect 25226 132826 25282 133626
rect 26054 132826 26110 133626
rect 26790 132826 26846 133626
rect 27526 132826 27582 133626
rect 28354 132826 28410 133626
rect 29090 132826 29146 133626
rect 29918 132826 29974 133626
rect 30654 132826 30710 133626
rect 31482 132826 31538 133626
rect 32218 132826 32274 133626
rect 33046 132826 33102 133626
rect 33782 132826 33838 133626
rect 34610 132826 34666 133626
rect 35346 132826 35402 133626
rect 36082 132826 36138 133626
rect 36910 132826 36966 133626
rect 37646 132826 37702 133626
rect 38474 132826 38530 133626
rect 39210 132826 39266 133626
rect 40038 132826 40094 133626
rect 40774 132826 40830 133626
rect 41602 132826 41658 133626
rect 42338 132826 42394 133626
rect 43166 132826 43222 133626
rect 43902 132826 43958 133626
rect 44638 132826 44694 133626
rect 45466 132826 45522 133626
rect 46202 132826 46258 133626
rect 47030 132826 47086 133626
rect 47766 132826 47822 133626
rect 48594 132826 48650 133626
rect 49330 132826 49386 133626
rect 50158 132826 50214 133626
rect 50894 132826 50950 133626
rect 51722 132826 51778 133626
rect 52458 132826 52514 133626
rect 53194 132826 53250 133626
rect 54022 132826 54078 133626
rect 54758 132826 54814 133626
rect 55586 132826 55642 133626
rect 56322 132826 56378 133626
rect 57150 132826 57206 133626
rect 57886 132826 57942 133626
rect 58714 132826 58770 133626
rect 59450 132826 59506 133626
rect 60278 132826 60334 133626
rect 61014 132826 61070 133626
rect 61750 132826 61806 133626
rect 62578 132826 62634 133626
rect 63314 132826 63370 133626
rect 64142 132826 64198 133626
rect 64878 132826 64934 133626
rect 65706 132826 65762 133626
rect 66442 132826 66498 133626
rect 67270 132826 67326 133626
rect 68006 132826 68062 133626
rect 68834 132826 68890 133626
rect 69570 132826 69626 133626
rect 70398 132826 70454 133626
rect 71134 132826 71190 133626
rect 71870 132826 71926 133626
rect 72698 132826 72754 133626
rect 73434 132826 73490 133626
rect 74262 132826 74318 133626
rect 74998 132826 75054 133626
rect 75826 132826 75882 133626
rect 76562 132826 76618 133626
rect 77390 132826 77446 133626
rect 78126 132826 78182 133626
rect 78954 132826 79010 133626
rect 79690 132826 79746 133626
rect 80426 132826 80482 133626
rect 81254 132826 81310 133626
rect 81990 132826 82046 133626
rect 82818 132826 82874 133626
rect 83554 132826 83610 133626
rect 84382 132826 84438 133626
rect 85118 132826 85174 133626
rect 85946 132826 86002 133626
rect 86682 132826 86738 133626
rect 87510 132826 87566 133626
rect 88246 132826 88302 133626
rect 88982 132826 89038 133626
rect 89810 132826 89866 133626
rect 90546 132826 90602 133626
rect 91374 132826 91430 133626
rect 92110 132826 92166 133626
rect 92938 132826 92994 133626
rect 93674 132826 93730 133626
rect 94502 132826 94558 133626
rect 95238 132826 95294 133626
rect 96066 132826 96122 133626
rect 96802 132826 96858 133626
rect 97538 132826 97594 133626
rect 98366 132826 98422 133626
rect 99102 132826 99158 133626
rect 99930 132826 99986 133626
rect 100666 132826 100722 133626
rect 101494 132826 101550 133626
rect 102230 132826 102286 133626
rect 103058 132826 103114 133626
rect 103794 132826 103850 133626
rect 104622 132826 104678 133626
rect 105358 132826 105414 133626
rect 106094 132826 106150 133626
rect 106922 132826 106978 133626
rect 107658 132826 107714 133626
rect 108486 132826 108542 133626
rect 109222 132826 109278 133626
rect 110050 132826 110106 133626
rect 110786 132826 110842 133626
rect 111614 132826 111670 133626
rect 112350 132826 112406 133626
rect 113178 132826 113234 133626
rect 113914 132826 113970 133626
rect 114650 132826 114706 133626
rect 115478 132826 115534 133626
rect 116214 132826 116270 133626
rect 117042 132826 117098 133626
rect 117778 132826 117834 133626
rect 118606 132826 118662 133626
rect 119342 132826 119398 133626
rect 120170 132826 120226 133626
rect 120906 132826 120962 133626
rect 121734 132826 121790 133626
rect 122470 132826 122526 133626
rect 123206 132826 123262 133626
rect 124034 132826 124090 133626
rect 124770 132826 124826 133626
rect 125598 132826 125654 133626
rect 126334 132826 126390 133626
rect 127162 132826 127218 133626
rect 127898 132826 127954 133626
rect 128726 132826 128782 133626
rect 129462 132826 129518 133626
rect 130290 132826 130346 133626
rect 131026 132826 131082 133626
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65798 0 65854 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83554 0 83610 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89810 0 89866 800
rect 89994 0 90050 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91834 0 91890 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97354 0 97410 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98274 0 98330 800
rect 98550 0 98606 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 100850 0 100906 800
rect 101126 0 101182 800
rect 101310 0 101366 800
rect 101586 0 101642 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104070 0 104126 800
rect 104346 0 104402 800
rect 104530 0 104586 800
rect 104806 0 104862 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105450 0 105506 800
rect 105726 0 105782 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106370 0 106426 800
rect 106646 0 106702 800
rect 106830 0 106886 800
rect 107106 0 107162 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111430 0 111486 800
rect 111706 0 111762 800
rect 111890 0 111946 800
rect 112166 0 112222 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113270 0 113326 800
rect 113546 0 113602 800
rect 113730 0 113786 800
rect 114006 0 114062 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116766 0 116822 800
rect 117042 0 117098 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117686 0 117742 800
rect 117962 0 118018 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118606 0 118662 800
rect 118882 0 118938 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 119986 0 120042 800
rect 120262 0 120318 800
rect 120446 0 120502 800
rect 120722 0 120778 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122286 0 122342 800
rect 122562 0 122618 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123206 0 123262 800
rect 123482 0 123538 800
rect 123666 0 123722 800
rect 123942 0 123998 800
rect 124126 0 124182 800
rect 124402 0 124458 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 125966 0 126022 800
rect 126242 0 126298 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127346 0 127402 800
rect 127622 0 127678 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129186 0 129242 800
rect 129462 0 129518 800
rect 129646 0 129702 800
rect 129922 0 129978 800
rect 130106 0 130162 800
rect 130382 0 130438 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131026 0 131082 800
rect 131302 0 131358 800
<< obsm2 >>
rect 20 132770 330 132954
rect 498 132770 1066 132954
rect 1234 132770 1802 132954
rect 1970 132770 2630 132954
rect 2798 132770 3366 132954
rect 3534 132770 4194 132954
rect 4362 132770 4930 132954
rect 5098 132770 5758 132954
rect 5926 132770 6494 132954
rect 6662 132770 7322 132954
rect 7490 132770 8058 132954
rect 8226 132770 8886 132954
rect 9054 132770 9622 132954
rect 9790 132770 10358 132954
rect 10526 132770 11186 132954
rect 11354 132770 11922 132954
rect 12090 132770 12750 132954
rect 12918 132770 13486 132954
rect 13654 132770 14314 132954
rect 14482 132770 15050 132954
rect 15218 132770 15878 132954
rect 16046 132770 16614 132954
rect 16782 132770 17442 132954
rect 17610 132770 18178 132954
rect 18346 132770 18914 132954
rect 19082 132770 19742 132954
rect 19910 132770 20478 132954
rect 20646 132770 21306 132954
rect 21474 132770 22042 132954
rect 22210 132770 22870 132954
rect 23038 132770 23606 132954
rect 23774 132770 24434 132954
rect 24602 132770 25170 132954
rect 25338 132770 25998 132954
rect 26166 132770 26734 132954
rect 26902 132770 27470 132954
rect 27638 132770 28298 132954
rect 28466 132770 29034 132954
rect 29202 132770 29862 132954
rect 30030 132770 30598 132954
rect 30766 132770 31426 132954
rect 31594 132770 32162 132954
rect 32330 132770 32990 132954
rect 33158 132770 33726 132954
rect 33894 132770 34554 132954
rect 34722 132770 35290 132954
rect 35458 132770 36026 132954
rect 36194 132770 36854 132954
rect 37022 132770 37590 132954
rect 37758 132770 38418 132954
rect 38586 132770 39154 132954
rect 39322 132770 39982 132954
rect 40150 132770 40718 132954
rect 40886 132770 41546 132954
rect 41714 132770 42282 132954
rect 42450 132770 43110 132954
rect 43278 132770 43846 132954
rect 44014 132770 44582 132954
rect 44750 132770 45410 132954
rect 45578 132770 46146 132954
rect 46314 132770 46974 132954
rect 47142 132770 47710 132954
rect 47878 132770 48538 132954
rect 48706 132770 49274 132954
rect 49442 132770 50102 132954
rect 50270 132770 50838 132954
rect 51006 132770 51666 132954
rect 51834 132770 52402 132954
rect 52570 132770 53138 132954
rect 53306 132770 53966 132954
rect 54134 132770 54702 132954
rect 54870 132770 55530 132954
rect 55698 132770 56266 132954
rect 56434 132770 57094 132954
rect 57262 132770 57830 132954
rect 57998 132770 58658 132954
rect 58826 132770 59394 132954
rect 59562 132770 60222 132954
rect 60390 132770 60958 132954
rect 61126 132770 61694 132954
rect 61862 132770 62522 132954
rect 62690 132770 63258 132954
rect 63426 132770 64086 132954
rect 64254 132770 64822 132954
rect 64990 132770 65650 132954
rect 65818 132770 66386 132954
rect 66554 132770 67214 132954
rect 67382 132770 67950 132954
rect 68118 132770 68778 132954
rect 68946 132770 69514 132954
rect 69682 132770 70342 132954
rect 70510 132770 71078 132954
rect 71246 132770 71814 132954
rect 71982 132770 72642 132954
rect 72810 132770 73378 132954
rect 73546 132770 74206 132954
rect 74374 132770 74942 132954
rect 75110 132770 75770 132954
rect 75938 132770 76506 132954
rect 76674 132770 77334 132954
rect 77502 132770 78070 132954
rect 78238 132770 78898 132954
rect 79066 132770 79634 132954
rect 79802 132770 80370 132954
rect 80538 132770 81198 132954
rect 81366 132770 81934 132954
rect 82102 132770 82762 132954
rect 82930 132770 83498 132954
rect 83666 132770 84326 132954
rect 84494 132770 85062 132954
rect 85230 132770 85890 132954
rect 86058 132770 86626 132954
rect 86794 132770 87454 132954
rect 87622 132770 88190 132954
rect 88358 132770 88926 132954
rect 89094 132770 89754 132954
rect 89922 132770 90490 132954
rect 90658 132770 91318 132954
rect 91486 132770 92054 132954
rect 92222 132770 92882 132954
rect 93050 132770 93618 132954
rect 93786 132770 94446 132954
rect 94614 132770 95182 132954
rect 95350 132770 96010 132954
rect 96178 132770 96746 132954
rect 96914 132770 97482 132954
rect 97650 132770 98310 132954
rect 98478 132770 99046 132954
rect 99214 132770 99874 132954
rect 100042 132770 100610 132954
rect 100778 132770 101438 132954
rect 101606 132770 102174 132954
rect 102342 132770 103002 132954
rect 103170 132770 103738 132954
rect 103906 132770 104566 132954
rect 104734 132770 105302 132954
rect 105470 132770 106038 132954
rect 106206 132770 106866 132954
rect 107034 132770 107602 132954
rect 107770 132770 108430 132954
rect 108598 132770 109166 132954
rect 109334 132770 109994 132954
rect 110162 132770 110730 132954
rect 110898 132770 111558 132954
rect 111726 132770 112294 132954
rect 112462 132770 113122 132954
rect 113290 132770 113858 132954
rect 114026 132770 114594 132954
rect 114762 132770 115422 132954
rect 115590 132770 116158 132954
rect 116326 132770 116986 132954
rect 117154 132770 117722 132954
rect 117890 132770 118550 132954
rect 118718 132770 119286 132954
rect 119454 132770 120114 132954
rect 120282 132770 120850 132954
rect 121018 132770 121678 132954
rect 121846 132770 122414 132954
rect 122582 132770 123150 132954
rect 123318 132770 123978 132954
rect 124146 132770 124714 132954
rect 124882 132770 125542 132954
rect 125710 132770 126278 132954
rect 126446 132770 127106 132954
rect 127274 132770 127842 132954
rect 128010 132770 128670 132954
rect 128838 132770 129406 132954
rect 129574 132770 130234 132954
rect 130402 132770 130970 132954
rect 131138 132770 131356 132954
rect 20 856 131356 132770
rect 20 342 54 856
rect 222 342 238 856
rect 406 342 514 856
rect 682 342 698 856
rect 866 342 974 856
rect 1142 342 1158 856
rect 1326 342 1434 856
rect 1602 342 1618 856
rect 1786 342 1894 856
rect 2062 342 2078 856
rect 2246 342 2354 856
rect 2522 342 2538 856
rect 2706 342 2814 856
rect 2982 342 2998 856
rect 3166 342 3274 856
rect 3442 342 3458 856
rect 3626 342 3734 856
rect 3902 342 3918 856
rect 4086 342 4194 856
rect 4362 342 4378 856
rect 4546 342 4654 856
rect 4822 342 4838 856
rect 5006 342 5114 856
rect 5282 342 5298 856
rect 5466 342 5574 856
rect 5742 342 5758 856
rect 5926 342 6034 856
rect 6202 342 6218 856
rect 6386 342 6494 856
rect 6662 342 6678 856
rect 6846 342 6954 856
rect 7122 342 7138 856
rect 7306 342 7414 856
rect 7582 342 7598 856
rect 7766 342 7874 856
rect 8042 342 8058 856
rect 8226 342 8334 856
rect 8502 342 8518 856
rect 8686 342 8794 856
rect 8962 342 8978 856
rect 9146 342 9254 856
rect 9422 342 9438 856
rect 9606 342 9714 856
rect 9882 342 9898 856
rect 10066 342 10174 856
rect 10342 342 10358 856
rect 10526 342 10634 856
rect 10802 342 10818 856
rect 10986 342 11094 856
rect 11262 342 11278 856
rect 11446 342 11554 856
rect 11722 342 11738 856
rect 11906 342 12014 856
rect 12182 342 12198 856
rect 12366 342 12474 856
rect 12642 342 12658 856
rect 12826 342 12934 856
rect 13102 342 13118 856
rect 13286 342 13394 856
rect 13562 342 13578 856
rect 13746 342 13854 856
rect 14022 342 14038 856
rect 14206 342 14314 856
rect 14482 342 14498 856
rect 14666 342 14774 856
rect 14942 342 14958 856
rect 15126 342 15234 856
rect 15402 342 15418 856
rect 15586 342 15694 856
rect 15862 342 15878 856
rect 16046 342 16154 856
rect 16322 342 16338 856
rect 16506 342 16614 856
rect 16782 342 16890 856
rect 17058 342 17074 856
rect 17242 342 17350 856
rect 17518 342 17534 856
rect 17702 342 17810 856
rect 17978 342 17994 856
rect 18162 342 18270 856
rect 18438 342 18454 856
rect 18622 342 18730 856
rect 18898 342 18914 856
rect 19082 342 19190 856
rect 19358 342 19374 856
rect 19542 342 19650 856
rect 19818 342 19834 856
rect 20002 342 20110 856
rect 20278 342 20294 856
rect 20462 342 20570 856
rect 20738 342 20754 856
rect 20922 342 21030 856
rect 21198 342 21214 856
rect 21382 342 21490 856
rect 21658 342 21674 856
rect 21842 342 21950 856
rect 22118 342 22134 856
rect 22302 342 22410 856
rect 22578 342 22594 856
rect 22762 342 22870 856
rect 23038 342 23054 856
rect 23222 342 23330 856
rect 23498 342 23514 856
rect 23682 342 23790 856
rect 23958 342 23974 856
rect 24142 342 24250 856
rect 24418 342 24434 856
rect 24602 342 24710 856
rect 24878 342 24894 856
rect 25062 342 25170 856
rect 25338 342 25354 856
rect 25522 342 25630 856
rect 25798 342 25814 856
rect 25982 342 26090 856
rect 26258 342 26274 856
rect 26442 342 26550 856
rect 26718 342 26734 856
rect 26902 342 27010 856
rect 27178 342 27194 856
rect 27362 342 27470 856
rect 27638 342 27654 856
rect 27822 342 27930 856
rect 28098 342 28114 856
rect 28282 342 28390 856
rect 28558 342 28574 856
rect 28742 342 28850 856
rect 29018 342 29034 856
rect 29202 342 29310 856
rect 29478 342 29494 856
rect 29662 342 29770 856
rect 29938 342 29954 856
rect 30122 342 30230 856
rect 30398 342 30414 856
rect 30582 342 30690 856
rect 30858 342 30874 856
rect 31042 342 31150 856
rect 31318 342 31334 856
rect 31502 342 31610 856
rect 31778 342 31794 856
rect 31962 342 32070 856
rect 32238 342 32254 856
rect 32422 342 32530 856
rect 32698 342 32714 856
rect 32882 342 32990 856
rect 33158 342 33266 856
rect 33434 342 33450 856
rect 33618 342 33726 856
rect 33894 342 33910 856
rect 34078 342 34186 856
rect 34354 342 34370 856
rect 34538 342 34646 856
rect 34814 342 34830 856
rect 34998 342 35106 856
rect 35274 342 35290 856
rect 35458 342 35566 856
rect 35734 342 35750 856
rect 35918 342 36026 856
rect 36194 342 36210 856
rect 36378 342 36486 856
rect 36654 342 36670 856
rect 36838 342 36946 856
rect 37114 342 37130 856
rect 37298 342 37406 856
rect 37574 342 37590 856
rect 37758 342 37866 856
rect 38034 342 38050 856
rect 38218 342 38326 856
rect 38494 342 38510 856
rect 38678 342 38786 856
rect 38954 342 38970 856
rect 39138 342 39246 856
rect 39414 342 39430 856
rect 39598 342 39706 856
rect 39874 342 39890 856
rect 40058 342 40166 856
rect 40334 342 40350 856
rect 40518 342 40626 856
rect 40794 342 40810 856
rect 40978 342 41086 856
rect 41254 342 41270 856
rect 41438 342 41546 856
rect 41714 342 41730 856
rect 41898 342 42006 856
rect 42174 342 42190 856
rect 42358 342 42466 856
rect 42634 342 42650 856
rect 42818 342 42926 856
rect 43094 342 43110 856
rect 43278 342 43386 856
rect 43554 342 43570 856
rect 43738 342 43846 856
rect 44014 342 44030 856
rect 44198 342 44306 856
rect 44474 342 44490 856
rect 44658 342 44766 856
rect 44934 342 44950 856
rect 45118 342 45226 856
rect 45394 342 45410 856
rect 45578 342 45686 856
rect 45854 342 45870 856
rect 46038 342 46146 856
rect 46314 342 46330 856
rect 46498 342 46606 856
rect 46774 342 46790 856
rect 46958 342 47066 856
rect 47234 342 47250 856
rect 47418 342 47526 856
rect 47694 342 47710 856
rect 47878 342 47986 856
rect 48154 342 48170 856
rect 48338 342 48446 856
rect 48614 342 48630 856
rect 48798 342 48906 856
rect 49074 342 49090 856
rect 49258 342 49366 856
rect 49534 342 49642 856
rect 49810 342 49826 856
rect 49994 342 50102 856
rect 50270 342 50286 856
rect 50454 342 50562 856
rect 50730 342 50746 856
rect 50914 342 51022 856
rect 51190 342 51206 856
rect 51374 342 51482 856
rect 51650 342 51666 856
rect 51834 342 51942 856
rect 52110 342 52126 856
rect 52294 342 52402 856
rect 52570 342 52586 856
rect 52754 342 52862 856
rect 53030 342 53046 856
rect 53214 342 53322 856
rect 53490 342 53506 856
rect 53674 342 53782 856
rect 53950 342 53966 856
rect 54134 342 54242 856
rect 54410 342 54426 856
rect 54594 342 54702 856
rect 54870 342 54886 856
rect 55054 342 55162 856
rect 55330 342 55346 856
rect 55514 342 55622 856
rect 55790 342 55806 856
rect 55974 342 56082 856
rect 56250 342 56266 856
rect 56434 342 56542 856
rect 56710 342 56726 856
rect 56894 342 57002 856
rect 57170 342 57186 856
rect 57354 342 57462 856
rect 57630 342 57646 856
rect 57814 342 57922 856
rect 58090 342 58106 856
rect 58274 342 58382 856
rect 58550 342 58566 856
rect 58734 342 58842 856
rect 59010 342 59026 856
rect 59194 342 59302 856
rect 59470 342 59486 856
rect 59654 342 59762 856
rect 59930 342 59946 856
rect 60114 342 60222 856
rect 60390 342 60406 856
rect 60574 342 60682 856
rect 60850 342 60866 856
rect 61034 342 61142 856
rect 61310 342 61326 856
rect 61494 342 61602 856
rect 61770 342 61786 856
rect 61954 342 62062 856
rect 62230 342 62246 856
rect 62414 342 62522 856
rect 62690 342 62706 856
rect 62874 342 62982 856
rect 63150 342 63166 856
rect 63334 342 63442 856
rect 63610 342 63626 856
rect 63794 342 63902 856
rect 64070 342 64086 856
rect 64254 342 64362 856
rect 64530 342 64546 856
rect 64714 342 64822 856
rect 64990 342 65006 856
rect 65174 342 65282 856
rect 65450 342 65466 856
rect 65634 342 65742 856
rect 65910 342 66018 856
rect 66186 342 66202 856
rect 66370 342 66478 856
rect 66646 342 66662 856
rect 66830 342 66938 856
rect 67106 342 67122 856
rect 67290 342 67398 856
rect 67566 342 67582 856
rect 67750 342 67858 856
rect 68026 342 68042 856
rect 68210 342 68318 856
rect 68486 342 68502 856
rect 68670 342 68778 856
rect 68946 342 68962 856
rect 69130 342 69238 856
rect 69406 342 69422 856
rect 69590 342 69698 856
rect 69866 342 69882 856
rect 70050 342 70158 856
rect 70326 342 70342 856
rect 70510 342 70618 856
rect 70786 342 70802 856
rect 70970 342 71078 856
rect 71246 342 71262 856
rect 71430 342 71538 856
rect 71706 342 71722 856
rect 71890 342 71998 856
rect 72166 342 72182 856
rect 72350 342 72458 856
rect 72626 342 72642 856
rect 72810 342 72918 856
rect 73086 342 73102 856
rect 73270 342 73378 856
rect 73546 342 73562 856
rect 73730 342 73838 856
rect 74006 342 74022 856
rect 74190 342 74298 856
rect 74466 342 74482 856
rect 74650 342 74758 856
rect 74926 342 74942 856
rect 75110 342 75218 856
rect 75386 342 75402 856
rect 75570 342 75678 856
rect 75846 342 75862 856
rect 76030 342 76138 856
rect 76306 342 76322 856
rect 76490 342 76598 856
rect 76766 342 76782 856
rect 76950 342 77058 856
rect 77226 342 77242 856
rect 77410 342 77518 856
rect 77686 342 77702 856
rect 77870 342 77978 856
rect 78146 342 78162 856
rect 78330 342 78438 856
rect 78606 342 78622 856
rect 78790 342 78898 856
rect 79066 342 79082 856
rect 79250 342 79358 856
rect 79526 342 79542 856
rect 79710 342 79818 856
rect 79986 342 80002 856
rect 80170 342 80278 856
rect 80446 342 80462 856
rect 80630 342 80738 856
rect 80906 342 80922 856
rect 81090 342 81198 856
rect 81366 342 81382 856
rect 81550 342 81658 856
rect 81826 342 81842 856
rect 82010 342 82118 856
rect 82286 342 82394 856
rect 82562 342 82578 856
rect 82746 342 82854 856
rect 83022 342 83038 856
rect 83206 342 83314 856
rect 83482 342 83498 856
rect 83666 342 83774 856
rect 83942 342 83958 856
rect 84126 342 84234 856
rect 84402 342 84418 856
rect 84586 342 84694 856
rect 84862 342 84878 856
rect 85046 342 85154 856
rect 85322 342 85338 856
rect 85506 342 85614 856
rect 85782 342 85798 856
rect 85966 342 86074 856
rect 86242 342 86258 856
rect 86426 342 86534 856
rect 86702 342 86718 856
rect 86886 342 86994 856
rect 87162 342 87178 856
rect 87346 342 87454 856
rect 87622 342 87638 856
rect 87806 342 87914 856
rect 88082 342 88098 856
rect 88266 342 88374 856
rect 88542 342 88558 856
rect 88726 342 88834 856
rect 89002 342 89018 856
rect 89186 342 89294 856
rect 89462 342 89478 856
rect 89646 342 89754 856
rect 89922 342 89938 856
rect 90106 342 90214 856
rect 90382 342 90398 856
rect 90566 342 90674 856
rect 90842 342 90858 856
rect 91026 342 91134 856
rect 91302 342 91318 856
rect 91486 342 91594 856
rect 91762 342 91778 856
rect 91946 342 92054 856
rect 92222 342 92238 856
rect 92406 342 92514 856
rect 92682 342 92698 856
rect 92866 342 92974 856
rect 93142 342 93158 856
rect 93326 342 93434 856
rect 93602 342 93618 856
rect 93786 342 93894 856
rect 94062 342 94078 856
rect 94246 342 94354 856
rect 94522 342 94538 856
rect 94706 342 94814 856
rect 94982 342 94998 856
rect 95166 342 95274 856
rect 95442 342 95458 856
rect 95626 342 95734 856
rect 95902 342 95918 856
rect 96086 342 96194 856
rect 96362 342 96378 856
rect 96546 342 96654 856
rect 96822 342 96838 856
rect 97006 342 97114 856
rect 97282 342 97298 856
rect 97466 342 97574 856
rect 97742 342 97758 856
rect 97926 342 98034 856
rect 98202 342 98218 856
rect 98386 342 98494 856
rect 98662 342 98770 856
rect 98938 342 98954 856
rect 99122 342 99230 856
rect 99398 342 99414 856
rect 99582 342 99690 856
rect 99858 342 99874 856
rect 100042 342 100150 856
rect 100318 342 100334 856
rect 100502 342 100610 856
rect 100778 342 100794 856
rect 100962 342 101070 856
rect 101238 342 101254 856
rect 101422 342 101530 856
rect 101698 342 101714 856
rect 101882 342 101990 856
rect 102158 342 102174 856
rect 102342 342 102450 856
rect 102618 342 102634 856
rect 102802 342 102910 856
rect 103078 342 103094 856
rect 103262 342 103370 856
rect 103538 342 103554 856
rect 103722 342 103830 856
rect 103998 342 104014 856
rect 104182 342 104290 856
rect 104458 342 104474 856
rect 104642 342 104750 856
rect 104918 342 104934 856
rect 105102 342 105210 856
rect 105378 342 105394 856
rect 105562 342 105670 856
rect 105838 342 105854 856
rect 106022 342 106130 856
rect 106298 342 106314 856
rect 106482 342 106590 856
rect 106758 342 106774 856
rect 106942 342 107050 856
rect 107218 342 107234 856
rect 107402 342 107510 856
rect 107678 342 107694 856
rect 107862 342 107970 856
rect 108138 342 108154 856
rect 108322 342 108430 856
rect 108598 342 108614 856
rect 108782 342 108890 856
rect 109058 342 109074 856
rect 109242 342 109350 856
rect 109518 342 109534 856
rect 109702 342 109810 856
rect 109978 342 109994 856
rect 110162 342 110270 856
rect 110438 342 110454 856
rect 110622 342 110730 856
rect 110898 342 110914 856
rect 111082 342 111190 856
rect 111358 342 111374 856
rect 111542 342 111650 856
rect 111818 342 111834 856
rect 112002 342 112110 856
rect 112278 342 112294 856
rect 112462 342 112570 856
rect 112738 342 112754 856
rect 112922 342 113030 856
rect 113198 342 113214 856
rect 113382 342 113490 856
rect 113658 342 113674 856
rect 113842 342 113950 856
rect 114118 342 114134 856
rect 114302 342 114410 856
rect 114578 342 114594 856
rect 114762 342 114870 856
rect 115038 342 115146 856
rect 115314 342 115330 856
rect 115498 342 115606 856
rect 115774 342 115790 856
rect 115958 342 116066 856
rect 116234 342 116250 856
rect 116418 342 116526 856
rect 116694 342 116710 856
rect 116878 342 116986 856
rect 117154 342 117170 856
rect 117338 342 117446 856
rect 117614 342 117630 856
rect 117798 342 117906 856
rect 118074 342 118090 856
rect 118258 342 118366 856
rect 118534 342 118550 856
rect 118718 342 118826 856
rect 118994 342 119010 856
rect 119178 342 119286 856
rect 119454 342 119470 856
rect 119638 342 119746 856
rect 119914 342 119930 856
rect 120098 342 120206 856
rect 120374 342 120390 856
rect 120558 342 120666 856
rect 120834 342 120850 856
rect 121018 342 121126 856
rect 121294 342 121310 856
rect 121478 342 121586 856
rect 121754 342 121770 856
rect 121938 342 122046 856
rect 122214 342 122230 856
rect 122398 342 122506 856
rect 122674 342 122690 856
rect 122858 342 122966 856
rect 123134 342 123150 856
rect 123318 342 123426 856
rect 123594 342 123610 856
rect 123778 342 123886 856
rect 124054 342 124070 856
rect 124238 342 124346 856
rect 124514 342 124530 856
rect 124698 342 124806 856
rect 124974 342 124990 856
rect 125158 342 125266 856
rect 125434 342 125450 856
rect 125618 342 125726 856
rect 125894 342 125910 856
rect 126078 342 126186 856
rect 126354 342 126370 856
rect 126538 342 126646 856
rect 126814 342 126830 856
rect 126998 342 127106 856
rect 127274 342 127290 856
rect 127458 342 127566 856
rect 127734 342 127750 856
rect 127918 342 128026 856
rect 128194 342 128210 856
rect 128378 342 128486 856
rect 128654 342 128670 856
rect 128838 342 128946 856
rect 129114 342 129130 856
rect 129298 342 129406 856
rect 129574 342 129590 856
rect 129758 342 129866 856
rect 130034 342 130050 856
rect 130218 342 130326 856
rect 130494 342 130510 856
rect 130678 342 130786 856
rect 130954 342 130970 856
rect 131138 342 131246 856
<< obsm3 >>
rect 1761 444 129615 131137
<< metal4 >>
rect 4208 2128 4528 131152
rect 19568 2128 19888 131152
rect 34928 2128 35248 131152
rect 50288 2128 50608 131152
rect 65648 2128 65968 131152
rect 81008 2128 81328 131152
rect 96368 2128 96688 131152
rect 111728 2128 112048 131152
rect 127088 2128 127408 131152
<< obsm4 >>
rect 1899 2048 4128 130797
rect 4608 2048 19488 130797
rect 19968 2048 34848 130797
rect 35328 2048 50208 130797
rect 50688 2048 65568 130797
rect 66048 2048 80928 130797
rect 81408 2048 96288 130797
rect 96768 2048 111648 130797
rect 112128 2048 127008 130797
rect 127488 2048 128557 130797
rect 1899 443 128557 2048
<< labels >>
rlabel metal2 s 2686 132826 2742 133626 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 5814 132826 5870 133626 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 8942 132826 8998 133626 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 11978 132826 12034 133626 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 15106 132826 15162 133626 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 17498 132826 17554 133626 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 19798 132826 19854 133626 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 22098 132826 22154 133626 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 24490 132826 24546 133626 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 386 132826 442 133626 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 1122 132826 1178 133626 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 3422 132826 3478 133626 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 28354 132826 28410 133626 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 29918 132826 29974 133626 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 31482 132826 31538 133626 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 33046 132826 33102 133626 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 34610 132826 34666 133626 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 36082 132826 36138 133626 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 37646 132826 37702 133626 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 39210 132826 39266 133626 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 40774 132826 40830 133626 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 42338 132826 42394 133626 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 6550 132826 6606 133626 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 43902 132826 43958 133626 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 45466 132826 45522 133626 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 47030 132826 47086 133626 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 48594 132826 48650 133626 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 50158 132826 50214 133626 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 51722 132826 51778 133626 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 53194 132826 53250 133626 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 54758 132826 54814 133626 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 56322 132826 56378 133626 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 57886 132826 57942 133626 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 9678 132826 9734 133626 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 59450 132826 59506 133626 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 61014 132826 61070 133626 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 12806 132826 12862 133626 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 15934 132826 15990 133626 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 18234 132826 18290 133626 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 20534 132826 20590 133626 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 22926 132826 22982 133626 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 25226 132826 25282 133626 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 26790 132826 26846 133626 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 4250 132826 4306 133626 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 29090 132826 29146 133626 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 30654 132826 30710 133626 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 32218 132826 32274 133626 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 33782 132826 33838 133626 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 35346 132826 35402 133626 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 36910 132826 36966 133626 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 38474 132826 38530 133626 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 40038 132826 40094 133626 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 41602 132826 41658 133626 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 43166 132826 43222 133626 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 7378 132826 7434 133626 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 44638 132826 44694 133626 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 46202 132826 46258 133626 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 47766 132826 47822 133626 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 49330 132826 49386 133626 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 50894 132826 50950 133626 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 52458 132826 52514 133626 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 54022 132826 54078 133626 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 55586 132826 55642 133626 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 57150 132826 57206 133626 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 58714 132826 58770 133626 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 10414 132826 10470 133626 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 60278 132826 60334 133626 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 61750 132826 61806 133626 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 13542 132826 13598 133626 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 16670 132826 16726 133626 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 18970 132826 19026 133626 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 21362 132826 21418 133626 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 23662 132826 23718 133626 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 26054 132826 26110 133626 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 27526 132826 27582 133626 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 1858 132826 1914 133626 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 4986 132826 5042 133626 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 8114 132826 8170 133626 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 11242 132826 11298 133626 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 14370 132826 14426 133626 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 64878 132826 64934 133626 6 gpio_in[0]
port 81 nsew signal input
rlabel metal2 s 88246 132826 88302 133626 6 gpio_in[10]
port 82 nsew signal input
rlabel metal2 s 90546 132826 90602 133626 6 gpio_in[11]
port 83 nsew signal input
rlabel metal2 s 92938 132826 92994 133626 6 gpio_in[12]
port 84 nsew signal input
rlabel metal2 s 95238 132826 95294 133626 6 gpio_in[13]
port 85 nsew signal input
rlabel metal2 s 97538 132826 97594 133626 6 gpio_in[14]
port 86 nsew signal input
rlabel metal2 s 99930 132826 99986 133626 6 gpio_in[15]
port 87 nsew signal input
rlabel metal2 s 102230 132826 102286 133626 6 gpio_in[16]
port 88 nsew signal input
rlabel metal2 s 104622 132826 104678 133626 6 gpio_in[17]
port 89 nsew signal input
rlabel metal2 s 106922 132826 106978 133626 6 gpio_in[18]
port 90 nsew signal input
rlabel metal2 s 109222 132826 109278 133626 6 gpio_in[19]
port 91 nsew signal input
rlabel metal2 s 67270 132826 67326 133626 6 gpio_in[1]
port 92 nsew signal input
rlabel metal2 s 111614 132826 111670 133626 6 gpio_in[20]
port 93 nsew signal input
rlabel metal2 s 113914 132826 113970 133626 6 gpio_in[21]
port 94 nsew signal input
rlabel metal2 s 116214 132826 116270 133626 6 gpio_in[22]
port 95 nsew signal input
rlabel metal2 s 118606 132826 118662 133626 6 gpio_in[23]
port 96 nsew signal input
rlabel metal2 s 69570 132826 69626 133626 6 gpio_in[2]
port 97 nsew signal input
rlabel metal2 s 71870 132826 71926 133626 6 gpio_in[3]
port 98 nsew signal input
rlabel metal2 s 74262 132826 74318 133626 6 gpio_in[4]
port 99 nsew signal input
rlabel metal2 s 76562 132826 76618 133626 6 gpio_in[5]
port 100 nsew signal input
rlabel metal2 s 78954 132826 79010 133626 6 gpio_in[6]
port 101 nsew signal input
rlabel metal2 s 81254 132826 81310 133626 6 gpio_in[7]
port 102 nsew signal input
rlabel metal2 s 83554 132826 83610 133626 6 gpio_in[8]
port 103 nsew signal input
rlabel metal2 s 85946 132826 86002 133626 6 gpio_in[9]
port 104 nsew signal input
rlabel metal2 s 65706 132826 65762 133626 6 gpio_oeb[0]
port 105 nsew signal output
rlabel metal2 s 88982 132826 89038 133626 6 gpio_oeb[10]
port 106 nsew signal output
rlabel metal2 s 91374 132826 91430 133626 6 gpio_oeb[11]
port 107 nsew signal output
rlabel metal2 s 93674 132826 93730 133626 6 gpio_oeb[12]
port 108 nsew signal output
rlabel metal2 s 96066 132826 96122 133626 6 gpio_oeb[13]
port 109 nsew signal output
rlabel metal2 s 98366 132826 98422 133626 6 gpio_oeb[14]
port 110 nsew signal output
rlabel metal2 s 100666 132826 100722 133626 6 gpio_oeb[15]
port 111 nsew signal output
rlabel metal2 s 103058 132826 103114 133626 6 gpio_oeb[16]
port 112 nsew signal output
rlabel metal2 s 105358 132826 105414 133626 6 gpio_oeb[17]
port 113 nsew signal output
rlabel metal2 s 107658 132826 107714 133626 6 gpio_oeb[18]
port 114 nsew signal output
rlabel metal2 s 110050 132826 110106 133626 6 gpio_oeb[19]
port 115 nsew signal output
rlabel metal2 s 68006 132826 68062 133626 6 gpio_oeb[1]
port 116 nsew signal output
rlabel metal2 s 112350 132826 112406 133626 6 gpio_oeb[20]
port 117 nsew signal output
rlabel metal2 s 114650 132826 114706 133626 6 gpio_oeb[21]
port 118 nsew signal output
rlabel metal2 s 117042 132826 117098 133626 6 gpio_oeb[22]
port 119 nsew signal output
rlabel metal2 s 119342 132826 119398 133626 6 gpio_oeb[23]
port 120 nsew signal output
rlabel metal2 s 120906 132826 120962 133626 6 gpio_oeb[24]
port 121 nsew signal output
rlabel metal2 s 121734 132826 121790 133626 6 gpio_oeb[25]
port 122 nsew signal output
rlabel metal2 s 122470 132826 122526 133626 6 gpio_oeb[26]
port 123 nsew signal output
rlabel metal2 s 123206 132826 123262 133626 6 gpio_oeb[27]
port 124 nsew signal output
rlabel metal2 s 124034 132826 124090 133626 6 gpio_oeb[28]
port 125 nsew signal output
rlabel metal2 s 124770 132826 124826 133626 6 gpio_oeb[29]
port 126 nsew signal output
rlabel metal2 s 70398 132826 70454 133626 6 gpio_oeb[2]
port 127 nsew signal output
rlabel metal2 s 125598 132826 125654 133626 6 gpio_oeb[30]
port 128 nsew signal output
rlabel metal2 s 126334 132826 126390 133626 6 gpio_oeb[31]
port 129 nsew signal output
rlabel metal2 s 127162 132826 127218 133626 6 gpio_oeb[32]
port 130 nsew signal output
rlabel metal2 s 127898 132826 127954 133626 6 gpio_oeb[33]
port 131 nsew signal output
rlabel metal2 s 128726 132826 128782 133626 6 gpio_oeb[34]
port 132 nsew signal output
rlabel metal2 s 129462 132826 129518 133626 6 gpio_oeb[35]
port 133 nsew signal output
rlabel metal2 s 130290 132826 130346 133626 6 gpio_oeb[36]
port 134 nsew signal output
rlabel metal2 s 131026 132826 131082 133626 6 gpio_oeb[37]
port 135 nsew signal output
rlabel metal2 s 72698 132826 72754 133626 6 gpio_oeb[3]
port 136 nsew signal output
rlabel metal2 s 74998 132826 75054 133626 6 gpio_oeb[4]
port 137 nsew signal output
rlabel metal2 s 77390 132826 77446 133626 6 gpio_oeb[5]
port 138 nsew signal output
rlabel metal2 s 79690 132826 79746 133626 6 gpio_oeb[6]
port 139 nsew signal output
rlabel metal2 s 81990 132826 82046 133626 6 gpio_oeb[7]
port 140 nsew signal output
rlabel metal2 s 84382 132826 84438 133626 6 gpio_oeb[8]
port 141 nsew signal output
rlabel metal2 s 86682 132826 86738 133626 6 gpio_oeb[9]
port 142 nsew signal output
rlabel metal2 s 66442 132826 66498 133626 6 gpio_out[0]
port 143 nsew signal output
rlabel metal2 s 89810 132826 89866 133626 6 gpio_out[10]
port 144 nsew signal output
rlabel metal2 s 92110 132826 92166 133626 6 gpio_out[11]
port 145 nsew signal output
rlabel metal2 s 94502 132826 94558 133626 6 gpio_out[12]
port 146 nsew signal output
rlabel metal2 s 96802 132826 96858 133626 6 gpio_out[13]
port 147 nsew signal output
rlabel metal2 s 99102 132826 99158 133626 6 gpio_out[14]
port 148 nsew signal output
rlabel metal2 s 101494 132826 101550 133626 6 gpio_out[15]
port 149 nsew signal output
rlabel metal2 s 103794 132826 103850 133626 6 gpio_out[16]
port 150 nsew signal output
rlabel metal2 s 106094 132826 106150 133626 6 gpio_out[17]
port 151 nsew signal output
rlabel metal2 s 108486 132826 108542 133626 6 gpio_out[18]
port 152 nsew signal output
rlabel metal2 s 110786 132826 110842 133626 6 gpio_out[19]
port 153 nsew signal output
rlabel metal2 s 68834 132826 68890 133626 6 gpio_out[1]
port 154 nsew signal output
rlabel metal2 s 113178 132826 113234 133626 6 gpio_out[20]
port 155 nsew signal output
rlabel metal2 s 115478 132826 115534 133626 6 gpio_out[21]
port 156 nsew signal output
rlabel metal2 s 117778 132826 117834 133626 6 gpio_out[22]
port 157 nsew signal output
rlabel metal2 s 120170 132826 120226 133626 6 gpio_out[23]
port 158 nsew signal output
rlabel metal2 s 71134 132826 71190 133626 6 gpio_out[2]
port 159 nsew signal output
rlabel metal2 s 73434 132826 73490 133626 6 gpio_out[3]
port 160 nsew signal output
rlabel metal2 s 75826 132826 75882 133626 6 gpio_out[4]
port 161 nsew signal output
rlabel metal2 s 78126 132826 78182 133626 6 gpio_out[5]
port 162 nsew signal output
rlabel metal2 s 80426 132826 80482 133626 6 gpio_out[6]
port 163 nsew signal output
rlabel metal2 s 82818 132826 82874 133626 6 gpio_out[7]
port 164 nsew signal output
rlabel metal2 s 85118 132826 85174 133626 6 gpio_out[8]
port 165 nsew signal output
rlabel metal2 s 87510 132826 87566 133626 6 gpio_out[9]
port 166 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 iram_addr0[0]
port 167 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 iram_addr0[1]
port 168 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 iram_addr0[2]
port 169 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 iram_addr0[3]
port 170 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 iram_addr0[4]
port 171 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 iram_addr0[5]
port 172 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 iram_addr0[6]
port 173 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 iram_addr0[7]
port 174 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 iram_addr0[8]
port 175 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 iram_clk0
port 176 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 iram_csb0
port 177 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 iram_din0[0]
port 178 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 iram_din0[10]
port 179 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 iram_din0[11]
port 180 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 iram_din0[12]
port 181 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 iram_din0[13]
port 182 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 iram_din0[14]
port 183 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 iram_din0[15]
port 184 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 iram_din0[16]
port 185 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 iram_din0[17]
port 186 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 iram_din0[18]
port 187 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 iram_din0[19]
port 188 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 iram_din0[1]
port 189 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 iram_din0[20]
port 190 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 iram_din0[21]
port 191 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 iram_din0[22]
port 192 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 iram_din0[23]
port 193 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 iram_din0[24]
port 194 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 iram_din0[25]
port 195 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 iram_din0[26]
port 196 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 iram_din0[27]
port 197 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 iram_din0[28]
port 198 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 iram_din0[29]
port 199 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 iram_din0[2]
port 200 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 iram_din0[30]
port 201 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 iram_din0[31]
port 202 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 iram_din0[3]
port 203 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 iram_din0[4]
port 204 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 iram_din0[5]
port 205 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 iram_din0[6]
port 206 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 iram_din0[7]
port 207 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 iram_din0[8]
port 208 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 iram_din0[9]
port 209 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 iram_dout0[0]
port 210 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 iram_dout0[10]
port 211 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 iram_dout0[11]
port 212 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 iram_dout0[12]
port 213 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 iram_dout0[13]
port 214 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 iram_dout0[14]
port 215 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 iram_dout0[15]
port 216 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 iram_dout0[16]
port 217 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 iram_dout0[17]
port 218 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 iram_dout0[18]
port 219 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 iram_dout0[19]
port 220 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 iram_dout0[1]
port 221 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 iram_dout0[20]
port 222 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 iram_dout0[21]
port 223 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 iram_dout0[22]
port 224 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 iram_dout0[23]
port 225 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 iram_dout0[24]
port 226 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 iram_dout0[25]
port 227 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 iram_dout0[26]
port 228 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 iram_dout0[27]
port 229 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 iram_dout0[28]
port 230 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 iram_dout0[29]
port 231 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 iram_dout0[2]
port 232 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 iram_dout0[30]
port 233 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 iram_dout0[31]
port 234 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 iram_dout0[3]
port 235 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 iram_dout0[4]
port 236 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 iram_dout0[5]
port 237 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 iram_dout0[6]
port 238 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 iram_dout0[7]
port 239 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 iram_dout0[8]
port 240 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 iram_dout0[9]
port 241 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 iram_web0
port 242 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 iram_wmask0[0]
port 243 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 iram_wmask0[1]
port 244 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 iram_wmask0[2]
port 245 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 iram_wmask0[3]
port 246 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 la_data_in[0]
port 247 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[100]
port 248 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[101]
port 249 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[102]
port 250 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[103]
port 251 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[104]
port 252 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[105]
port 253 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[106]
port 254 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[107]
port 255 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[108]
port 256 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[109]
port 257 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[10]
port 258 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[110]
port 259 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[111]
port 260 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[112]
port 261 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[113]
port 262 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[114]
port 263 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[115]
port 264 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[116]
port 265 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[117]
port 266 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[118]
port 267 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[119]
port 268 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_in[11]
port 269 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[120]
port 270 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[121]
port 271 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[122]
port 272 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[123]
port 273 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[124]
port 274 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_data_in[125]
port 275 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[126]
port 276 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[127]
port 277 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_data_in[12]
port 278 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[13]
port 279 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[14]
port 280 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[15]
port 281 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[16]
port 282 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[17]
port 283 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[18]
port 284 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in[19]
port 285 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[1]
port 286 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[20]
port 287 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[21]
port 288 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[22]
port 289 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[23]
port 290 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[24]
port 291 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[25]
port 292 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[26]
port 293 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[27]
port 294 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[28]
port 295 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[29]
port 296 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[2]
port 297 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[30]
port 298 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[31]
port 299 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[32]
port 300 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[33]
port 301 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[34]
port 302 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[35]
port 303 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[36]
port 304 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[37]
port 305 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[38]
port 306 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[39]
port 307 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_data_in[3]
port 308 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[40]
port 309 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[41]
port 310 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[42]
port 311 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[43]
port 312 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[44]
port 313 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[45]
port 314 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[46]
port 315 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[47]
port 316 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[48]
port 317 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[49]
port 318 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_data_in[4]
port 319 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[50]
port 320 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[51]
port 321 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[52]
port 322 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[53]
port 323 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[54]
port 324 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[55]
port 325 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[56]
port 326 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[57]
port 327 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[58]
port 328 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[59]
port 329 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_data_in[5]
port 330 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[60]
port 331 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[61]
port 332 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[62]
port 333 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[63]
port 334 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[64]
port 335 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[65]
port 336 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[66]
port 337 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[67]
port 338 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[68]
port 339 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[69]
port 340 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_data_in[6]
port 341 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[70]
port 342 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[71]
port 343 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[72]
port 344 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[73]
port 345 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[74]
port 346 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[75]
port 347 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[76]
port 348 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[77]
port 349 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[78]
port 350 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[79]
port 351 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_data_in[7]
port 352 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[80]
port 353 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[81]
port 354 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[82]
port 355 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[83]
port 356 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[84]
port 357 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[85]
port 358 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[86]
port 359 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[87]
port 360 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[88]
port 361 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[89]
port 362 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[8]
port 363 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_data_in[90]
port 364 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[91]
port 365 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[92]
port 366 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[93]
port 367 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[94]
port 368 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[95]
port 369 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[96]
port 370 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[97]
port 371 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[98]
port 372 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[99]
port 373 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[9]
port 374 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_out[0]
port 375 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[100]
port 376 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[101]
port 377 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[102]
port 378 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[103]
port 379 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[104]
port 380 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[105]
port 381 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[106]
port 382 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[107]
port 383 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[108]
port 384 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[109]
port 385 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 la_data_out[10]
port 386 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[110]
port 387 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[111]
port 388 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[112]
port 389 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[113]
port 390 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[114]
port 391 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[115]
port 392 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[116]
port 393 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[117]
port 394 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[118]
port 395 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[119]
port 396 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 la_data_out[11]
port 397 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[120]
port 398 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[121]
port 399 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 la_data_out[122]
port 400 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[123]
port 401 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[124]
port 402 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[125]
port 403 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 la_data_out[126]
port 404 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[127]
port 405 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[12]
port 406 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[13]
port 407 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_out[14]
port 408 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[15]
port 409 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[16]
port 410 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[17]
port 411 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la_data_out[18]
port 412 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 la_data_out[19]
port 413 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 la_data_out[1]
port 414 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[20]
port 415 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[21]
port 416 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[22]
port 417 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[23]
port 418 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[24]
port 419 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[25]
port 420 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[26]
port 421 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_out[27]
port 422 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[28]
port 423 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[29]
port 424 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 la_data_out[2]
port 425 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[30]
port 426 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[31]
port 427 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[32]
port 428 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[33]
port 429 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[34]
port 430 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[35]
port 431 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 la_data_out[36]
port 432 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[37]
port 433 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[38]
port 434 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[39]
port 435 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[3]
port 436 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[40]
port 437 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[41]
port 438 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[42]
port 439 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[43]
port 440 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[44]
port 441 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[45]
port 442 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[46]
port 443 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[47]
port 444 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[48]
port 445 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[49]
port 446 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[4]
port 447 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[50]
port 448 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[51]
port 449 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[52]
port 450 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[53]
port 451 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[54]
port 452 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[55]
port 453 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[56]
port 454 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[57]
port 455 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[58]
port 456 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 la_data_out[59]
port 457 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 la_data_out[5]
port 458 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[60]
port 459 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[61]
port 460 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[62]
port 461 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[63]
port 462 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[64]
port 463 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[65]
port 464 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[66]
port 465 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[67]
port 466 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[68]
port 467 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[69]
port 468 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 la_data_out[6]
port 469 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[70]
port 470 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[71]
port 471 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[72]
port 472 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[73]
port 473 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[74]
port 474 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[75]
port 475 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[76]
port 476 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[77]
port 477 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[78]
port 478 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[79]
port 479 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[7]
port 480 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[80]
port 481 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[81]
port 482 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[82]
port 483 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[83]
port 484 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[84]
port 485 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[85]
port 486 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[86]
port 487 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[87]
port 488 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[88]
port 489 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[89]
port 490 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[8]
port 491 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[90]
port 492 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[91]
port 493 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[92]
port 494 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[93]
port 495 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[94]
port 496 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[95]
port 497 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[96]
port 498 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[97]
port 499 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[98]
port 500 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[99]
port 501 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[9]
port 502 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_oenb[0]
port 503 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[100]
port 504 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[101]
port 505 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[102]
port 506 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[103]
port 507 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[104]
port 508 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[105]
port 509 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[106]
port 510 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[107]
port 511 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[108]
port 512 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[109]
port 513 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_oenb[10]
port 514 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[110]
port 515 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[111]
port 516 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[112]
port 517 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[113]
port 518 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[114]
port 519 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_oenb[115]
port 520 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[116]
port 521 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[117]
port 522 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[118]
port 523 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[119]
port 524 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_oenb[11]
port 525 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_oenb[120]
port 526 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[121]
port 527 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[122]
port 528 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[123]
port 529 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_oenb[124]
port 530 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[125]
port 531 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[126]
port 532 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_oenb[127]
port 533 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[12]
port 534 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[13]
port 535 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[14]
port 536 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[15]
port 537 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[16]
port 538 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[17]
port 539 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[18]
port 540 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_oenb[19]
port 541 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[1]
port 542 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_oenb[20]
port 543 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[21]
port 544 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[22]
port 545 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[23]
port 546 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[24]
port 547 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[25]
port 548 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[26]
port 549 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_oenb[27]
port 550 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[28]
port 551 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[29]
port 552 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[2]
port 553 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[30]
port 554 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[31]
port 555 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[32]
port 556 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[33]
port 557 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[34]
port 558 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[35]
port 559 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_oenb[36]
port 560 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[37]
port 561 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[38]
port 562 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[39]
port 563 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_oenb[3]
port 564 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[40]
port 565 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_oenb[41]
port 566 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[42]
port 567 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[43]
port 568 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[44]
port 569 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[45]
port 570 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[46]
port 571 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[47]
port 572 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[48]
port 573 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[49]
port 574 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[4]
port 575 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[50]
port 576 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[51]
port 577 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[52]
port 578 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[53]
port 579 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[54]
port 580 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[55]
port 581 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_oenb[56]
port 582 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[57]
port 583 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[58]
port 584 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[59]
port 585 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[5]
port 586 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[60]
port 587 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[61]
port 588 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_oenb[62]
port 589 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[63]
port 590 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[64]
port 591 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[65]
port 592 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[66]
port 593 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[67]
port 594 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[68]
port 595 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[69]
port 596 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_oenb[6]
port 597 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[70]
port 598 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[71]
port 599 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[72]
port 600 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[73]
port 601 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[74]
port 602 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[75]
port 603 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[76]
port 604 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[77]
port 605 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[78]
port 606 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[79]
port 607 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_oenb[7]
port 608 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[80]
port 609 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[81]
port 610 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[82]
port 611 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[83]
port 612 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[84]
port 613 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[85]
port 614 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_oenb[86]
port 615 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[87]
port 616 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[88]
port 617 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[89]
port 618 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[8]
port 619 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[90]
port 620 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[91]
port 621 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[92]
port 622 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[93]
port 623 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[94]
port 624 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[95]
port 625 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[96]
port 626 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[97]
port 627 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[98]
port 628 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[99]
port 629 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[9]
port 630 nsew signal input
rlabel metal2 s 62578 132826 62634 133626 6 user_irq[0]
port 631 nsew signal output
rlabel metal2 s 63314 132826 63370 133626 6 user_irq[1]
port 632 nsew signal output
rlabel metal2 s 64142 132826 64198 133626 6 user_irq[2]
port 633 nsew signal output
rlabel metal4 s 4208 2128 4528 131152 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 131152 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 131152 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 131152 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 131152 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 131152 6 vssd1
port 635 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 131152 6 vssd1
port 635 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 131152 6 vssd1
port 635 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 131152 6 vssd1
port 635 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 636 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 637 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_ack_o
port 638 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 wbs_adr_i[0]
port 639 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[10]
port 640 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[11]
port 641 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[12]
port 642 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[13]
port 643 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[14]
port 644 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[15]
port 645 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[16]
port 646 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[17]
port 647 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[18]
port 648 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[19]
port 649 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_adr_i[1]
port 650 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[20]
port 651 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[21]
port 652 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[22]
port 653 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[23]
port 654 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[24]
port 655 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[25]
port 656 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[26]
port 657 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[27]
port 658 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[28]
port 659 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[29]
port 660 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[2]
port 661 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[30]
port 662 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[31]
port 663 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[3]
port 664 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[4]
port 665 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[5]
port 666 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[6]
port 667 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[7]
port 668 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[8]
port 669 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[9]
port 670 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 671 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_i[0]
port 672 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[10]
port 673 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[11]
port 674 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[12]
port 675 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[13]
port 676 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[14]
port 677 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[15]
port 678 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[16]
port 679 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[17]
port 680 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[18]
port 681 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[19]
port 682 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[1]
port 683 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[20]
port 684 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[21]
port 685 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[22]
port 686 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_i[23]
port 687 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[24]
port 688 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[25]
port 689 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[26]
port 690 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[27]
port 691 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[28]
port 692 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[29]
port 693 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_i[2]
port 694 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[30]
port 695 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[31]
port 696 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[3]
port 697 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[4]
port 698 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_i[5]
port 699 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[6]
port 700 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[7]
port 701 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[8]
port 702 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[9]
port 703 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[0]
port 704 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[10]
port 705 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[11]
port 706 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[12]
port 707 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[13]
port 708 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[14]
port 709 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[15]
port 710 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[16]
port 711 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[17]
port 712 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[18]
port 713 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[19]
port 714 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_o[1]
port 715 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[20]
port 716 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[21]
port 717 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[22]
port 718 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[23]
port 719 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[24]
port 720 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[25]
port 721 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[26]
port 722 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[27]
port 723 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[28]
port 724 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[29]
port 725 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_o[2]
port 726 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[30]
port 727 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[31]
port 728 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[3]
port 729 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_o[4]
port 730 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[5]
port 731 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_o[6]
port 732 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[7]
port 733 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[8]
port 734 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[9]
port 735 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wbs_sel_i[0]
port 736 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_sel_i[1]
port 737 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[2]
port 738 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[3]
port 739 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_stb_i
port 740 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_we_i
port 741 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 131482 133626
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44471376
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/rvj1_caravel_soc/runs/rvj1_caravel_soc/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1315206
<< end >>

