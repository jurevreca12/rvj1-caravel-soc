magic
tech sky130A
magscale 1 2
timestamp 1653944247
<< obsli1 >>
rect 1104 2159 127880 128945
<< obsm1 >>
rect 290 280 128970 129804
<< metal2 >>
rect 294 130344 350 131144
rect 938 130344 994 131144
rect 1582 130344 1638 131144
rect 2226 130344 2282 131144
rect 2870 130344 2926 131144
rect 3514 130344 3570 131144
rect 4158 130344 4214 131144
rect 4802 130344 4858 131144
rect 5446 130344 5502 131144
rect 6182 130344 6238 131144
rect 6826 130344 6882 131144
rect 7470 130344 7526 131144
rect 8114 130344 8170 131144
rect 8758 130344 8814 131144
rect 9402 130344 9458 131144
rect 10046 130344 10102 131144
rect 10690 130344 10746 131144
rect 11334 130344 11390 131144
rect 12070 130344 12126 131144
rect 12714 130344 12770 131144
rect 13358 130344 13414 131144
rect 14002 130344 14058 131144
rect 14646 130344 14702 131144
rect 15290 130344 15346 131144
rect 15934 130344 15990 131144
rect 16578 130344 16634 131144
rect 17314 130344 17370 131144
rect 17958 130344 18014 131144
rect 18602 130344 18658 131144
rect 19246 130344 19302 131144
rect 19890 130344 19946 131144
rect 20534 130344 20590 131144
rect 21178 130344 21234 131144
rect 21822 130344 21878 131144
rect 22466 130344 22522 131144
rect 23202 130344 23258 131144
rect 23846 130344 23902 131144
rect 24490 130344 24546 131144
rect 25134 130344 25190 131144
rect 25778 130344 25834 131144
rect 26422 130344 26478 131144
rect 27066 130344 27122 131144
rect 27710 130344 27766 131144
rect 28446 130344 28502 131144
rect 29090 130344 29146 131144
rect 29734 130344 29790 131144
rect 30378 130344 30434 131144
rect 31022 130344 31078 131144
rect 31666 130344 31722 131144
rect 32310 130344 32366 131144
rect 32954 130344 33010 131144
rect 33598 130344 33654 131144
rect 34334 130344 34390 131144
rect 34978 130344 35034 131144
rect 35622 130344 35678 131144
rect 36266 130344 36322 131144
rect 36910 130344 36966 131144
rect 37554 130344 37610 131144
rect 38198 130344 38254 131144
rect 38842 130344 38898 131144
rect 39578 130344 39634 131144
rect 40222 130344 40278 131144
rect 40866 130344 40922 131144
rect 41510 130344 41566 131144
rect 42154 130344 42210 131144
rect 42798 130344 42854 131144
rect 43442 130344 43498 131144
rect 44086 130344 44142 131144
rect 44730 130344 44786 131144
rect 45466 130344 45522 131144
rect 46110 130344 46166 131144
rect 46754 130344 46810 131144
rect 47398 130344 47454 131144
rect 48042 130344 48098 131144
rect 48686 130344 48742 131144
rect 49330 130344 49386 131144
rect 49974 130344 50030 131144
rect 50618 130344 50674 131144
rect 51354 130344 51410 131144
rect 51998 130344 52054 131144
rect 52642 130344 52698 131144
rect 53286 130344 53342 131144
rect 53930 130344 53986 131144
rect 54574 130344 54630 131144
rect 55218 130344 55274 131144
rect 55862 130344 55918 131144
rect 56598 130344 56654 131144
rect 57242 130344 57298 131144
rect 57886 130344 57942 131144
rect 58530 130344 58586 131144
rect 59174 130344 59230 131144
rect 59818 130344 59874 131144
rect 60462 130344 60518 131144
rect 61106 130344 61162 131144
rect 61750 130344 61806 131144
rect 62486 130344 62542 131144
rect 63130 130344 63186 131144
rect 63774 130344 63830 131144
rect 64418 130344 64474 131144
rect 65062 130344 65118 131144
rect 65706 130344 65762 131144
rect 66350 130344 66406 131144
rect 66994 130344 67050 131144
rect 67730 130344 67786 131144
rect 68374 130344 68430 131144
rect 69018 130344 69074 131144
rect 69662 130344 69718 131144
rect 70306 130344 70362 131144
rect 70950 130344 71006 131144
rect 71594 130344 71650 131144
rect 72238 130344 72294 131144
rect 72882 130344 72938 131144
rect 73618 130344 73674 131144
rect 74262 130344 74318 131144
rect 74906 130344 74962 131144
rect 75550 130344 75606 131144
rect 76194 130344 76250 131144
rect 76838 130344 76894 131144
rect 77482 130344 77538 131144
rect 78126 130344 78182 131144
rect 78862 130344 78918 131144
rect 79506 130344 79562 131144
rect 80150 130344 80206 131144
rect 80794 130344 80850 131144
rect 81438 130344 81494 131144
rect 82082 130344 82138 131144
rect 82726 130344 82782 131144
rect 83370 130344 83426 131144
rect 84014 130344 84070 131144
rect 84750 130344 84806 131144
rect 85394 130344 85450 131144
rect 86038 130344 86094 131144
rect 86682 130344 86738 131144
rect 87326 130344 87382 131144
rect 87970 130344 88026 131144
rect 88614 130344 88670 131144
rect 89258 130344 89314 131144
rect 89902 130344 89958 131144
rect 90638 130344 90694 131144
rect 91282 130344 91338 131144
rect 91926 130344 91982 131144
rect 92570 130344 92626 131144
rect 93214 130344 93270 131144
rect 93858 130344 93914 131144
rect 94502 130344 94558 131144
rect 95146 130344 95202 131144
rect 95882 130344 95938 131144
rect 96526 130344 96582 131144
rect 97170 130344 97226 131144
rect 97814 130344 97870 131144
rect 98458 130344 98514 131144
rect 99102 130344 99158 131144
rect 99746 130344 99802 131144
rect 100390 130344 100446 131144
rect 101034 130344 101090 131144
rect 101770 130344 101826 131144
rect 102414 130344 102470 131144
rect 103058 130344 103114 131144
rect 103702 130344 103758 131144
rect 104346 130344 104402 131144
rect 104990 130344 105046 131144
rect 105634 130344 105690 131144
rect 106278 130344 106334 131144
rect 107014 130344 107070 131144
rect 107658 130344 107714 131144
rect 108302 130344 108358 131144
rect 108946 130344 109002 131144
rect 109590 130344 109646 131144
rect 110234 130344 110290 131144
rect 110878 130344 110934 131144
rect 111522 130344 111578 131144
rect 112166 130344 112222 131144
rect 112902 130344 112958 131144
rect 113546 130344 113602 131144
rect 114190 130344 114246 131144
rect 114834 130344 114890 131144
rect 115478 130344 115534 131144
rect 116122 130344 116178 131144
rect 116766 130344 116822 131144
rect 117410 130344 117466 131144
rect 118146 130344 118202 131144
rect 118790 130344 118846 131144
rect 119434 130344 119490 131144
rect 120078 130344 120134 131144
rect 120722 130344 120778 131144
rect 121366 130344 121422 131144
rect 122010 130344 122066 131144
rect 122654 130344 122710 131144
rect 123298 130344 123354 131144
rect 124034 130344 124090 131144
rect 124678 130344 124734 131144
rect 125322 130344 125378 131144
rect 125966 130344 126022 131144
rect 126610 130344 126666 131144
rect 127254 130344 127310 131144
rect 127898 130344 127954 131144
rect 128542 130344 128598 131144
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7286 0 7342 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82082 0 82138 800
rect 82266 0 82322 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87418 0 87474 800
rect 87602 0 87658 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91466 0 91522 800
rect 91650 0 91706 800
rect 91834 0 91890 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 95882 0 95938 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97170 0 97226 800
rect 97354 0 97410 800
rect 97538 0 97594 800
rect 97722 0 97778 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98366 0 98422 800
rect 98550 0 98606 800
rect 98734 0 98790 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
rect 100022 0 100078 800
rect 100206 0 100262 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101034 0 101090 800
rect 101218 0 101274 800
rect 101402 0 101458 800
rect 101586 0 101642 800
rect 101770 0 101826 800
rect 101954 0 102010 800
rect 102138 0 102194 800
rect 102322 0 102378 800
rect 102506 0 102562 800
rect 102690 0 102746 800
rect 102874 0 102930 800
rect 103058 0 103114 800
rect 103334 0 103390 800
rect 103518 0 103574 800
rect 103702 0 103758 800
rect 103886 0 103942 800
rect 104070 0 104126 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104806 0 104862 800
rect 104990 0 105046 800
rect 105174 0 105230 800
rect 105358 0 105414 800
rect 105542 0 105598 800
rect 105726 0 105782 800
rect 106002 0 106058 800
rect 106186 0 106242 800
rect 106370 0 106426 800
rect 106554 0 106610 800
rect 106738 0 106794 800
rect 106922 0 106978 800
rect 107106 0 107162 800
rect 107290 0 107346 800
rect 107474 0 107530 800
rect 107658 0 107714 800
rect 107842 0 107898 800
rect 108026 0 108082 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108670 0 108726 800
rect 108854 0 108910 800
rect 109038 0 109094 800
rect 109222 0 109278 800
rect 109406 0 109462 800
rect 109590 0 109646 800
rect 109774 0 109830 800
rect 109958 0 110014 800
rect 110142 0 110198 800
rect 110326 0 110382 800
rect 110510 0 110566 800
rect 110694 0 110750 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111338 0 111394 800
rect 111522 0 111578 800
rect 111706 0 111762 800
rect 111890 0 111946 800
rect 112074 0 112130 800
rect 112258 0 112314 800
rect 112442 0 112498 800
rect 112626 0 112682 800
rect 112810 0 112866 800
rect 112994 0 113050 800
rect 113178 0 113234 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 113822 0 113878 800
rect 114006 0 114062 800
rect 114190 0 114246 800
rect 114374 0 114430 800
rect 114558 0 114614 800
rect 114742 0 114798 800
rect 114926 0 114982 800
rect 115110 0 115166 800
rect 115294 0 115350 800
rect 115478 0 115534 800
rect 115662 0 115718 800
rect 115846 0 115902 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116490 0 116546 800
rect 116674 0 116730 800
rect 116858 0 116914 800
rect 117042 0 117098 800
rect 117226 0 117282 800
rect 117410 0 117466 800
rect 117594 0 117650 800
rect 117778 0 117834 800
rect 117962 0 118018 800
rect 118146 0 118202 800
rect 118330 0 118386 800
rect 118514 0 118570 800
rect 118790 0 118846 800
rect 118974 0 119030 800
rect 119158 0 119214 800
rect 119342 0 119398 800
rect 119526 0 119582 800
rect 119710 0 119766 800
rect 119894 0 119950 800
rect 120078 0 120134 800
rect 120262 0 120318 800
rect 120446 0 120502 800
rect 120630 0 120686 800
rect 120814 0 120870 800
rect 120998 0 121054 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121642 0 121698 800
rect 121826 0 121882 800
rect 122010 0 122066 800
rect 122194 0 122250 800
rect 122378 0 122434 800
rect 122562 0 122618 800
rect 122746 0 122802 800
rect 122930 0 122986 800
rect 123114 0 123170 800
rect 123298 0 123354 800
rect 123482 0 123538 800
rect 123666 0 123722 800
rect 123942 0 123998 800
rect 124126 0 124182 800
rect 124310 0 124366 800
rect 124494 0 124550 800
rect 124678 0 124734 800
rect 124862 0 124918 800
rect 125046 0 125102 800
rect 125230 0 125286 800
rect 125414 0 125470 800
rect 125598 0 125654 800
rect 125782 0 125838 800
rect 125966 0 126022 800
rect 126150 0 126206 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126794 0 126850 800
rect 126978 0 127034 800
rect 127162 0 127218 800
rect 127346 0 127402 800
rect 127530 0 127586 800
rect 127714 0 127770 800
rect 127898 0 127954 800
rect 128082 0 128138 800
rect 128266 0 128322 800
rect 128450 0 128506 800
rect 128634 0 128690 800
rect 128818 0 128874 800
<< obsm2 >>
rect 18 130288 238 130506
rect 406 130288 882 130506
rect 1050 130288 1526 130506
rect 1694 130288 2170 130506
rect 2338 130288 2814 130506
rect 2982 130288 3458 130506
rect 3626 130288 4102 130506
rect 4270 130288 4746 130506
rect 4914 130288 5390 130506
rect 5558 130288 6126 130506
rect 6294 130288 6770 130506
rect 6938 130288 7414 130506
rect 7582 130288 8058 130506
rect 8226 130288 8702 130506
rect 8870 130288 9346 130506
rect 9514 130288 9990 130506
rect 10158 130288 10634 130506
rect 10802 130288 11278 130506
rect 11446 130288 12014 130506
rect 12182 130288 12658 130506
rect 12826 130288 13302 130506
rect 13470 130288 13946 130506
rect 14114 130288 14590 130506
rect 14758 130288 15234 130506
rect 15402 130288 15878 130506
rect 16046 130288 16522 130506
rect 16690 130288 17258 130506
rect 17426 130288 17902 130506
rect 18070 130288 18546 130506
rect 18714 130288 19190 130506
rect 19358 130288 19834 130506
rect 20002 130288 20478 130506
rect 20646 130288 21122 130506
rect 21290 130288 21766 130506
rect 21934 130288 22410 130506
rect 22578 130288 23146 130506
rect 23314 130288 23790 130506
rect 23958 130288 24434 130506
rect 24602 130288 25078 130506
rect 25246 130288 25722 130506
rect 25890 130288 26366 130506
rect 26534 130288 27010 130506
rect 27178 130288 27654 130506
rect 27822 130288 28390 130506
rect 28558 130288 29034 130506
rect 29202 130288 29678 130506
rect 29846 130288 30322 130506
rect 30490 130288 30966 130506
rect 31134 130288 31610 130506
rect 31778 130288 32254 130506
rect 32422 130288 32898 130506
rect 33066 130288 33542 130506
rect 33710 130288 34278 130506
rect 34446 130288 34922 130506
rect 35090 130288 35566 130506
rect 35734 130288 36210 130506
rect 36378 130288 36854 130506
rect 37022 130288 37498 130506
rect 37666 130288 38142 130506
rect 38310 130288 38786 130506
rect 38954 130288 39522 130506
rect 39690 130288 40166 130506
rect 40334 130288 40810 130506
rect 40978 130288 41454 130506
rect 41622 130288 42098 130506
rect 42266 130288 42742 130506
rect 42910 130288 43386 130506
rect 43554 130288 44030 130506
rect 44198 130288 44674 130506
rect 44842 130288 45410 130506
rect 45578 130288 46054 130506
rect 46222 130288 46698 130506
rect 46866 130288 47342 130506
rect 47510 130288 47986 130506
rect 48154 130288 48630 130506
rect 48798 130288 49274 130506
rect 49442 130288 49918 130506
rect 50086 130288 50562 130506
rect 50730 130288 51298 130506
rect 51466 130288 51942 130506
rect 52110 130288 52586 130506
rect 52754 130288 53230 130506
rect 53398 130288 53874 130506
rect 54042 130288 54518 130506
rect 54686 130288 55162 130506
rect 55330 130288 55806 130506
rect 55974 130288 56542 130506
rect 56710 130288 57186 130506
rect 57354 130288 57830 130506
rect 57998 130288 58474 130506
rect 58642 130288 59118 130506
rect 59286 130288 59762 130506
rect 59930 130288 60406 130506
rect 60574 130288 61050 130506
rect 61218 130288 61694 130506
rect 61862 130288 62430 130506
rect 62598 130288 63074 130506
rect 63242 130288 63718 130506
rect 63886 130288 64362 130506
rect 64530 130288 65006 130506
rect 65174 130288 65650 130506
rect 65818 130288 66294 130506
rect 66462 130288 66938 130506
rect 67106 130288 67674 130506
rect 67842 130288 68318 130506
rect 68486 130288 68962 130506
rect 69130 130288 69606 130506
rect 69774 130288 70250 130506
rect 70418 130288 70894 130506
rect 71062 130288 71538 130506
rect 71706 130288 72182 130506
rect 72350 130288 72826 130506
rect 72994 130288 73562 130506
rect 73730 130288 74206 130506
rect 74374 130288 74850 130506
rect 75018 130288 75494 130506
rect 75662 130288 76138 130506
rect 76306 130288 76782 130506
rect 76950 130288 77426 130506
rect 77594 130288 78070 130506
rect 78238 130288 78806 130506
rect 78974 130288 79450 130506
rect 79618 130288 80094 130506
rect 80262 130288 80738 130506
rect 80906 130288 81382 130506
rect 81550 130288 82026 130506
rect 82194 130288 82670 130506
rect 82838 130288 83314 130506
rect 83482 130288 83958 130506
rect 84126 130288 84694 130506
rect 84862 130288 85338 130506
rect 85506 130288 85982 130506
rect 86150 130288 86626 130506
rect 86794 130288 87270 130506
rect 87438 130288 87914 130506
rect 88082 130288 88558 130506
rect 88726 130288 89202 130506
rect 89370 130288 89846 130506
rect 90014 130288 90582 130506
rect 90750 130288 91226 130506
rect 91394 130288 91870 130506
rect 92038 130288 92514 130506
rect 92682 130288 93158 130506
rect 93326 130288 93802 130506
rect 93970 130288 94446 130506
rect 94614 130288 95090 130506
rect 95258 130288 95826 130506
rect 95994 130288 96470 130506
rect 96638 130288 97114 130506
rect 97282 130288 97758 130506
rect 97926 130288 98402 130506
rect 98570 130288 99046 130506
rect 99214 130288 99690 130506
rect 99858 130288 100334 130506
rect 100502 130288 100978 130506
rect 101146 130288 101714 130506
rect 101882 130288 102358 130506
rect 102526 130288 103002 130506
rect 103170 130288 103646 130506
rect 103814 130288 104290 130506
rect 104458 130288 104934 130506
rect 105102 130288 105578 130506
rect 105746 130288 106222 130506
rect 106390 130288 106958 130506
rect 107126 130288 107602 130506
rect 107770 130288 108246 130506
rect 108414 130288 108890 130506
rect 109058 130288 109534 130506
rect 109702 130288 110178 130506
rect 110346 130288 110822 130506
rect 110990 130288 111466 130506
rect 111634 130288 112110 130506
rect 112278 130288 112846 130506
rect 113014 130288 113490 130506
rect 113658 130288 114134 130506
rect 114302 130288 114778 130506
rect 114946 130288 115422 130506
rect 115590 130288 116066 130506
rect 116234 130288 116710 130506
rect 116878 130288 117354 130506
rect 117522 130288 118090 130506
rect 118258 130288 118734 130506
rect 118902 130288 119378 130506
rect 119546 130288 120022 130506
rect 120190 130288 120666 130506
rect 120834 130288 121310 130506
rect 121478 130288 121954 130506
rect 122122 130288 122598 130506
rect 122766 130288 123242 130506
rect 123410 130288 123978 130506
rect 124146 130288 124622 130506
rect 124790 130288 125266 130506
rect 125434 130288 125910 130506
rect 126078 130288 126554 130506
rect 126722 130288 127198 130506
rect 127366 130288 127842 130506
rect 128010 130288 128486 130506
rect 128654 130288 128964 130506
rect 18 856 128964 130288
rect 18 274 54 856
rect 222 274 238 856
rect 406 274 422 856
rect 590 274 606 856
rect 774 274 790 856
rect 958 274 974 856
rect 1142 274 1158 856
rect 1326 274 1342 856
rect 1510 274 1526 856
rect 1694 274 1710 856
rect 1878 274 1894 856
rect 2062 274 2078 856
rect 2246 274 2262 856
rect 2430 274 2446 856
rect 2614 274 2722 856
rect 2890 274 2906 856
rect 3074 274 3090 856
rect 3258 274 3274 856
rect 3442 274 3458 856
rect 3626 274 3642 856
rect 3810 274 3826 856
rect 3994 274 4010 856
rect 4178 274 4194 856
rect 4362 274 4378 856
rect 4546 274 4562 856
rect 4730 274 4746 856
rect 4914 274 4930 856
rect 5098 274 5114 856
rect 5282 274 5390 856
rect 5558 274 5574 856
rect 5742 274 5758 856
rect 5926 274 5942 856
rect 6110 274 6126 856
rect 6294 274 6310 856
rect 6478 274 6494 856
rect 6662 274 6678 856
rect 6846 274 6862 856
rect 7030 274 7046 856
rect 7214 274 7230 856
rect 7398 274 7414 856
rect 7582 274 7598 856
rect 7766 274 7874 856
rect 8042 274 8058 856
rect 8226 274 8242 856
rect 8410 274 8426 856
rect 8594 274 8610 856
rect 8778 274 8794 856
rect 8962 274 8978 856
rect 9146 274 9162 856
rect 9330 274 9346 856
rect 9514 274 9530 856
rect 9698 274 9714 856
rect 9882 274 9898 856
rect 10066 274 10082 856
rect 10250 274 10266 856
rect 10434 274 10542 856
rect 10710 274 10726 856
rect 10894 274 10910 856
rect 11078 274 11094 856
rect 11262 274 11278 856
rect 11446 274 11462 856
rect 11630 274 11646 856
rect 11814 274 11830 856
rect 11998 274 12014 856
rect 12182 274 12198 856
rect 12366 274 12382 856
rect 12550 274 12566 856
rect 12734 274 12750 856
rect 12918 274 13026 856
rect 13194 274 13210 856
rect 13378 274 13394 856
rect 13562 274 13578 856
rect 13746 274 13762 856
rect 13930 274 13946 856
rect 14114 274 14130 856
rect 14298 274 14314 856
rect 14482 274 14498 856
rect 14666 274 14682 856
rect 14850 274 14866 856
rect 15034 274 15050 856
rect 15218 274 15234 856
rect 15402 274 15418 856
rect 15586 274 15694 856
rect 15862 274 15878 856
rect 16046 274 16062 856
rect 16230 274 16246 856
rect 16414 274 16430 856
rect 16598 274 16614 856
rect 16782 274 16798 856
rect 16966 274 16982 856
rect 17150 274 17166 856
rect 17334 274 17350 856
rect 17518 274 17534 856
rect 17702 274 17718 856
rect 17886 274 17902 856
rect 18070 274 18178 856
rect 18346 274 18362 856
rect 18530 274 18546 856
rect 18714 274 18730 856
rect 18898 274 18914 856
rect 19082 274 19098 856
rect 19266 274 19282 856
rect 19450 274 19466 856
rect 19634 274 19650 856
rect 19818 274 19834 856
rect 20002 274 20018 856
rect 20186 274 20202 856
rect 20370 274 20386 856
rect 20554 274 20570 856
rect 20738 274 20846 856
rect 21014 274 21030 856
rect 21198 274 21214 856
rect 21382 274 21398 856
rect 21566 274 21582 856
rect 21750 274 21766 856
rect 21934 274 21950 856
rect 22118 274 22134 856
rect 22302 274 22318 856
rect 22486 274 22502 856
rect 22670 274 22686 856
rect 22854 274 22870 856
rect 23038 274 23054 856
rect 23222 274 23330 856
rect 23498 274 23514 856
rect 23682 274 23698 856
rect 23866 274 23882 856
rect 24050 274 24066 856
rect 24234 274 24250 856
rect 24418 274 24434 856
rect 24602 274 24618 856
rect 24786 274 24802 856
rect 24970 274 24986 856
rect 25154 274 25170 856
rect 25338 274 25354 856
rect 25522 274 25538 856
rect 25706 274 25722 856
rect 25890 274 25998 856
rect 26166 274 26182 856
rect 26350 274 26366 856
rect 26534 274 26550 856
rect 26718 274 26734 856
rect 26902 274 26918 856
rect 27086 274 27102 856
rect 27270 274 27286 856
rect 27454 274 27470 856
rect 27638 274 27654 856
rect 27822 274 27838 856
rect 28006 274 28022 856
rect 28190 274 28206 856
rect 28374 274 28482 856
rect 28650 274 28666 856
rect 28834 274 28850 856
rect 29018 274 29034 856
rect 29202 274 29218 856
rect 29386 274 29402 856
rect 29570 274 29586 856
rect 29754 274 29770 856
rect 29938 274 29954 856
rect 30122 274 30138 856
rect 30306 274 30322 856
rect 30490 274 30506 856
rect 30674 274 30690 856
rect 30858 274 30874 856
rect 31042 274 31150 856
rect 31318 274 31334 856
rect 31502 274 31518 856
rect 31686 274 31702 856
rect 31870 274 31886 856
rect 32054 274 32070 856
rect 32238 274 32254 856
rect 32422 274 32438 856
rect 32606 274 32622 856
rect 32790 274 32806 856
rect 32974 274 32990 856
rect 33158 274 33174 856
rect 33342 274 33358 856
rect 33526 274 33634 856
rect 33802 274 33818 856
rect 33986 274 34002 856
rect 34170 274 34186 856
rect 34354 274 34370 856
rect 34538 274 34554 856
rect 34722 274 34738 856
rect 34906 274 34922 856
rect 35090 274 35106 856
rect 35274 274 35290 856
rect 35458 274 35474 856
rect 35642 274 35658 856
rect 35826 274 35842 856
rect 36010 274 36026 856
rect 36194 274 36302 856
rect 36470 274 36486 856
rect 36654 274 36670 856
rect 36838 274 36854 856
rect 37022 274 37038 856
rect 37206 274 37222 856
rect 37390 274 37406 856
rect 37574 274 37590 856
rect 37758 274 37774 856
rect 37942 274 37958 856
rect 38126 274 38142 856
rect 38310 274 38326 856
rect 38494 274 38510 856
rect 38678 274 38786 856
rect 38954 274 38970 856
rect 39138 274 39154 856
rect 39322 274 39338 856
rect 39506 274 39522 856
rect 39690 274 39706 856
rect 39874 274 39890 856
rect 40058 274 40074 856
rect 40242 274 40258 856
rect 40426 274 40442 856
rect 40610 274 40626 856
rect 40794 274 40810 856
rect 40978 274 40994 856
rect 41162 274 41178 856
rect 41346 274 41454 856
rect 41622 274 41638 856
rect 41806 274 41822 856
rect 41990 274 42006 856
rect 42174 274 42190 856
rect 42358 274 42374 856
rect 42542 274 42558 856
rect 42726 274 42742 856
rect 42910 274 42926 856
rect 43094 274 43110 856
rect 43278 274 43294 856
rect 43462 274 43478 856
rect 43646 274 43662 856
rect 43830 274 43938 856
rect 44106 274 44122 856
rect 44290 274 44306 856
rect 44474 274 44490 856
rect 44658 274 44674 856
rect 44842 274 44858 856
rect 45026 274 45042 856
rect 45210 274 45226 856
rect 45394 274 45410 856
rect 45578 274 45594 856
rect 45762 274 45778 856
rect 45946 274 45962 856
rect 46130 274 46146 856
rect 46314 274 46330 856
rect 46498 274 46606 856
rect 46774 274 46790 856
rect 46958 274 46974 856
rect 47142 274 47158 856
rect 47326 274 47342 856
rect 47510 274 47526 856
rect 47694 274 47710 856
rect 47878 274 47894 856
rect 48062 274 48078 856
rect 48246 274 48262 856
rect 48430 274 48446 856
rect 48614 274 48630 856
rect 48798 274 48814 856
rect 48982 274 49090 856
rect 49258 274 49274 856
rect 49442 274 49458 856
rect 49626 274 49642 856
rect 49810 274 49826 856
rect 49994 274 50010 856
rect 50178 274 50194 856
rect 50362 274 50378 856
rect 50546 274 50562 856
rect 50730 274 50746 856
rect 50914 274 50930 856
rect 51098 274 51114 856
rect 51282 274 51298 856
rect 51466 274 51482 856
rect 51650 274 51758 856
rect 51926 274 51942 856
rect 52110 274 52126 856
rect 52294 274 52310 856
rect 52478 274 52494 856
rect 52662 274 52678 856
rect 52846 274 52862 856
rect 53030 274 53046 856
rect 53214 274 53230 856
rect 53398 274 53414 856
rect 53582 274 53598 856
rect 53766 274 53782 856
rect 53950 274 53966 856
rect 54134 274 54242 856
rect 54410 274 54426 856
rect 54594 274 54610 856
rect 54778 274 54794 856
rect 54962 274 54978 856
rect 55146 274 55162 856
rect 55330 274 55346 856
rect 55514 274 55530 856
rect 55698 274 55714 856
rect 55882 274 55898 856
rect 56066 274 56082 856
rect 56250 274 56266 856
rect 56434 274 56450 856
rect 56618 274 56634 856
rect 56802 274 56910 856
rect 57078 274 57094 856
rect 57262 274 57278 856
rect 57446 274 57462 856
rect 57630 274 57646 856
rect 57814 274 57830 856
rect 57998 274 58014 856
rect 58182 274 58198 856
rect 58366 274 58382 856
rect 58550 274 58566 856
rect 58734 274 58750 856
rect 58918 274 58934 856
rect 59102 274 59118 856
rect 59286 274 59394 856
rect 59562 274 59578 856
rect 59746 274 59762 856
rect 59930 274 59946 856
rect 60114 274 60130 856
rect 60298 274 60314 856
rect 60482 274 60498 856
rect 60666 274 60682 856
rect 60850 274 60866 856
rect 61034 274 61050 856
rect 61218 274 61234 856
rect 61402 274 61418 856
rect 61586 274 61602 856
rect 61770 274 61786 856
rect 61954 274 62062 856
rect 62230 274 62246 856
rect 62414 274 62430 856
rect 62598 274 62614 856
rect 62782 274 62798 856
rect 62966 274 62982 856
rect 63150 274 63166 856
rect 63334 274 63350 856
rect 63518 274 63534 856
rect 63702 274 63718 856
rect 63886 274 63902 856
rect 64070 274 64086 856
rect 64254 274 64270 856
rect 64438 274 64546 856
rect 64714 274 64730 856
rect 64898 274 64914 856
rect 65082 274 65098 856
rect 65266 274 65282 856
rect 65450 274 65466 856
rect 65634 274 65650 856
rect 65818 274 65834 856
rect 66002 274 66018 856
rect 66186 274 66202 856
rect 66370 274 66386 856
rect 66554 274 66570 856
rect 66738 274 66754 856
rect 66922 274 66938 856
rect 67106 274 67214 856
rect 67382 274 67398 856
rect 67566 274 67582 856
rect 67750 274 67766 856
rect 67934 274 67950 856
rect 68118 274 68134 856
rect 68302 274 68318 856
rect 68486 274 68502 856
rect 68670 274 68686 856
rect 68854 274 68870 856
rect 69038 274 69054 856
rect 69222 274 69238 856
rect 69406 274 69422 856
rect 69590 274 69606 856
rect 69774 274 69882 856
rect 70050 274 70066 856
rect 70234 274 70250 856
rect 70418 274 70434 856
rect 70602 274 70618 856
rect 70786 274 70802 856
rect 70970 274 70986 856
rect 71154 274 71170 856
rect 71338 274 71354 856
rect 71522 274 71538 856
rect 71706 274 71722 856
rect 71890 274 71906 856
rect 72074 274 72090 856
rect 72258 274 72366 856
rect 72534 274 72550 856
rect 72718 274 72734 856
rect 72902 274 72918 856
rect 73086 274 73102 856
rect 73270 274 73286 856
rect 73454 274 73470 856
rect 73638 274 73654 856
rect 73822 274 73838 856
rect 74006 274 74022 856
rect 74190 274 74206 856
rect 74374 274 74390 856
rect 74558 274 74574 856
rect 74742 274 74758 856
rect 74926 274 75034 856
rect 75202 274 75218 856
rect 75386 274 75402 856
rect 75570 274 75586 856
rect 75754 274 75770 856
rect 75938 274 75954 856
rect 76122 274 76138 856
rect 76306 274 76322 856
rect 76490 274 76506 856
rect 76674 274 76690 856
rect 76858 274 76874 856
rect 77042 274 77058 856
rect 77226 274 77242 856
rect 77410 274 77518 856
rect 77686 274 77702 856
rect 77870 274 77886 856
rect 78054 274 78070 856
rect 78238 274 78254 856
rect 78422 274 78438 856
rect 78606 274 78622 856
rect 78790 274 78806 856
rect 78974 274 78990 856
rect 79158 274 79174 856
rect 79342 274 79358 856
rect 79526 274 79542 856
rect 79710 274 79726 856
rect 79894 274 79910 856
rect 80078 274 80186 856
rect 80354 274 80370 856
rect 80538 274 80554 856
rect 80722 274 80738 856
rect 80906 274 80922 856
rect 81090 274 81106 856
rect 81274 274 81290 856
rect 81458 274 81474 856
rect 81642 274 81658 856
rect 81826 274 81842 856
rect 82010 274 82026 856
rect 82194 274 82210 856
rect 82378 274 82394 856
rect 82562 274 82670 856
rect 82838 274 82854 856
rect 83022 274 83038 856
rect 83206 274 83222 856
rect 83390 274 83406 856
rect 83574 274 83590 856
rect 83758 274 83774 856
rect 83942 274 83958 856
rect 84126 274 84142 856
rect 84310 274 84326 856
rect 84494 274 84510 856
rect 84678 274 84694 856
rect 84862 274 84878 856
rect 85046 274 85062 856
rect 85230 274 85338 856
rect 85506 274 85522 856
rect 85690 274 85706 856
rect 85874 274 85890 856
rect 86058 274 86074 856
rect 86242 274 86258 856
rect 86426 274 86442 856
rect 86610 274 86626 856
rect 86794 274 86810 856
rect 86978 274 86994 856
rect 87162 274 87178 856
rect 87346 274 87362 856
rect 87530 274 87546 856
rect 87714 274 87822 856
rect 87990 274 88006 856
rect 88174 274 88190 856
rect 88358 274 88374 856
rect 88542 274 88558 856
rect 88726 274 88742 856
rect 88910 274 88926 856
rect 89094 274 89110 856
rect 89278 274 89294 856
rect 89462 274 89478 856
rect 89646 274 89662 856
rect 89830 274 89846 856
rect 90014 274 90030 856
rect 90198 274 90214 856
rect 90382 274 90490 856
rect 90658 274 90674 856
rect 90842 274 90858 856
rect 91026 274 91042 856
rect 91210 274 91226 856
rect 91394 274 91410 856
rect 91578 274 91594 856
rect 91762 274 91778 856
rect 91946 274 91962 856
rect 92130 274 92146 856
rect 92314 274 92330 856
rect 92498 274 92514 856
rect 92682 274 92698 856
rect 92866 274 92974 856
rect 93142 274 93158 856
rect 93326 274 93342 856
rect 93510 274 93526 856
rect 93694 274 93710 856
rect 93878 274 93894 856
rect 94062 274 94078 856
rect 94246 274 94262 856
rect 94430 274 94446 856
rect 94614 274 94630 856
rect 94798 274 94814 856
rect 94982 274 94998 856
rect 95166 274 95182 856
rect 95350 274 95366 856
rect 95534 274 95642 856
rect 95810 274 95826 856
rect 95994 274 96010 856
rect 96178 274 96194 856
rect 96362 274 96378 856
rect 96546 274 96562 856
rect 96730 274 96746 856
rect 96914 274 96930 856
rect 97098 274 97114 856
rect 97282 274 97298 856
rect 97466 274 97482 856
rect 97650 274 97666 856
rect 97834 274 97850 856
rect 98018 274 98126 856
rect 98294 274 98310 856
rect 98478 274 98494 856
rect 98662 274 98678 856
rect 98846 274 98862 856
rect 99030 274 99046 856
rect 99214 274 99230 856
rect 99398 274 99414 856
rect 99582 274 99598 856
rect 99766 274 99782 856
rect 99950 274 99966 856
rect 100134 274 100150 856
rect 100318 274 100334 856
rect 100502 274 100518 856
rect 100686 274 100794 856
rect 100962 274 100978 856
rect 101146 274 101162 856
rect 101330 274 101346 856
rect 101514 274 101530 856
rect 101698 274 101714 856
rect 101882 274 101898 856
rect 102066 274 102082 856
rect 102250 274 102266 856
rect 102434 274 102450 856
rect 102618 274 102634 856
rect 102802 274 102818 856
rect 102986 274 103002 856
rect 103170 274 103278 856
rect 103446 274 103462 856
rect 103630 274 103646 856
rect 103814 274 103830 856
rect 103998 274 104014 856
rect 104182 274 104198 856
rect 104366 274 104382 856
rect 104550 274 104566 856
rect 104734 274 104750 856
rect 104918 274 104934 856
rect 105102 274 105118 856
rect 105286 274 105302 856
rect 105470 274 105486 856
rect 105654 274 105670 856
rect 105838 274 105946 856
rect 106114 274 106130 856
rect 106298 274 106314 856
rect 106482 274 106498 856
rect 106666 274 106682 856
rect 106850 274 106866 856
rect 107034 274 107050 856
rect 107218 274 107234 856
rect 107402 274 107418 856
rect 107586 274 107602 856
rect 107770 274 107786 856
rect 107954 274 107970 856
rect 108138 274 108154 856
rect 108322 274 108430 856
rect 108598 274 108614 856
rect 108782 274 108798 856
rect 108966 274 108982 856
rect 109150 274 109166 856
rect 109334 274 109350 856
rect 109518 274 109534 856
rect 109702 274 109718 856
rect 109886 274 109902 856
rect 110070 274 110086 856
rect 110254 274 110270 856
rect 110438 274 110454 856
rect 110622 274 110638 856
rect 110806 274 110822 856
rect 110990 274 111098 856
rect 111266 274 111282 856
rect 111450 274 111466 856
rect 111634 274 111650 856
rect 111818 274 111834 856
rect 112002 274 112018 856
rect 112186 274 112202 856
rect 112370 274 112386 856
rect 112554 274 112570 856
rect 112738 274 112754 856
rect 112922 274 112938 856
rect 113106 274 113122 856
rect 113290 274 113306 856
rect 113474 274 113582 856
rect 113750 274 113766 856
rect 113934 274 113950 856
rect 114118 274 114134 856
rect 114302 274 114318 856
rect 114486 274 114502 856
rect 114670 274 114686 856
rect 114854 274 114870 856
rect 115038 274 115054 856
rect 115222 274 115238 856
rect 115406 274 115422 856
rect 115590 274 115606 856
rect 115774 274 115790 856
rect 115958 274 115974 856
rect 116142 274 116250 856
rect 116418 274 116434 856
rect 116602 274 116618 856
rect 116786 274 116802 856
rect 116970 274 116986 856
rect 117154 274 117170 856
rect 117338 274 117354 856
rect 117522 274 117538 856
rect 117706 274 117722 856
rect 117890 274 117906 856
rect 118074 274 118090 856
rect 118258 274 118274 856
rect 118442 274 118458 856
rect 118626 274 118734 856
rect 118902 274 118918 856
rect 119086 274 119102 856
rect 119270 274 119286 856
rect 119454 274 119470 856
rect 119638 274 119654 856
rect 119822 274 119838 856
rect 120006 274 120022 856
rect 120190 274 120206 856
rect 120374 274 120390 856
rect 120558 274 120574 856
rect 120742 274 120758 856
rect 120926 274 120942 856
rect 121110 274 121126 856
rect 121294 274 121402 856
rect 121570 274 121586 856
rect 121754 274 121770 856
rect 121938 274 121954 856
rect 122122 274 122138 856
rect 122306 274 122322 856
rect 122490 274 122506 856
rect 122674 274 122690 856
rect 122858 274 122874 856
rect 123042 274 123058 856
rect 123226 274 123242 856
rect 123410 274 123426 856
rect 123594 274 123610 856
rect 123778 274 123886 856
rect 124054 274 124070 856
rect 124238 274 124254 856
rect 124422 274 124438 856
rect 124606 274 124622 856
rect 124790 274 124806 856
rect 124974 274 124990 856
rect 125158 274 125174 856
rect 125342 274 125358 856
rect 125526 274 125542 856
rect 125710 274 125726 856
rect 125894 274 125910 856
rect 126078 274 126094 856
rect 126262 274 126278 856
rect 126446 274 126554 856
rect 126722 274 126738 856
rect 126906 274 126922 856
rect 127090 274 127106 856
rect 127274 274 127290 856
rect 127458 274 127474 856
rect 127642 274 127658 856
rect 127826 274 127842 856
rect 128010 274 128026 856
rect 128194 274 128210 856
rect 128378 274 128394 856
rect 128562 274 128578 856
rect 128746 274 128762 856
rect 128930 274 128964 856
<< obsm3 >>
rect 13 579 128787 129709
<< metal4 >>
rect 4208 2128 4528 128976
rect 19568 2128 19888 128976
rect 34928 2128 35248 128976
rect 50288 2128 50608 128976
rect 65648 2128 65968 128976
rect 81008 2128 81328 128976
rect 96368 2128 96688 128976
rect 111728 2128 112048 128976
rect 127088 2128 127408 128976
<< obsm4 >>
rect 1899 129056 125981 129709
rect 1899 2048 4128 129056
rect 4608 2048 19488 129056
rect 19968 2048 34848 129056
rect 35328 2048 50208 129056
rect 50688 2048 65568 129056
rect 66048 2048 80928 129056
rect 81408 2048 96288 129056
rect 96768 2048 111648 129056
rect 112128 2048 125981 129056
rect 1899 851 125981 2048
<< labels >>
rlabel metal2 s 76838 130344 76894 131144 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 79506 130344 79562 131144 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 82082 130344 82138 131144 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 84750 130344 84806 131144 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 87326 130344 87382 131144 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 89258 130344 89314 131144 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 91282 130344 91338 131144 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 93214 130344 93270 131144 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 95146 130344 95202 131144 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 74906 130344 74962 131144 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 75550 130344 75606 131144 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 77482 130344 77538 131144 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 98458 130344 98514 131144 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 99746 130344 99802 131144 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 101034 130344 101090 131144 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 102414 130344 102470 131144 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 103702 130344 103758 131144 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 104990 130344 105046 131144 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 106278 130344 106334 131144 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 107658 130344 107714 131144 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 108946 130344 109002 131144 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 110234 130344 110290 131144 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 80150 130344 80206 131144 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 111522 130344 111578 131144 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 112902 130344 112958 131144 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 114190 130344 114246 131144 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 115478 130344 115534 131144 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 116766 130344 116822 131144 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 118146 130344 118202 131144 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 119434 130344 119490 131144 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 120722 130344 120778 131144 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 122010 130344 122066 131144 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 123298 130344 123354 131144 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 82726 130344 82782 131144 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 124678 130344 124734 131144 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 125966 130344 126022 131144 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 85394 130344 85450 131144 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 87970 130344 88026 131144 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 89902 130344 89958 131144 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 91926 130344 91982 131144 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 93858 130344 93914 131144 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 95882 130344 95938 131144 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 97170 130344 97226 131144 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 78126 130344 78182 131144 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 99102 130344 99158 131144 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 100390 130344 100446 131144 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 101770 130344 101826 131144 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 103058 130344 103114 131144 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 104346 130344 104402 131144 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 105634 130344 105690 131144 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 107014 130344 107070 131144 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 108302 130344 108358 131144 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 109590 130344 109646 131144 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 110878 130344 110934 131144 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 80794 130344 80850 131144 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 112166 130344 112222 131144 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 113546 130344 113602 131144 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 114834 130344 114890 131144 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 116122 130344 116178 131144 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 117410 130344 117466 131144 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 118790 130344 118846 131144 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 120078 130344 120134 131144 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 121366 130344 121422 131144 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 122654 130344 122710 131144 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 124034 130344 124090 131144 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 83370 130344 83426 131144 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 125322 130344 125378 131144 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 126610 130344 126666 131144 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 86038 130344 86094 131144 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 88614 130344 88670 131144 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 90638 130344 90694 131144 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 92570 130344 92626 131144 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 94502 130344 94558 131144 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 96526 130344 96582 131144 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 97814 130344 97870 131144 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 76194 130344 76250 131144 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 78862 130344 78918 131144 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 81438 130344 81494 131144 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 84014 130344 84070 131144 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 86682 130344 86738 131144 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 294 130344 350 131144 6 io_in[0]
port 81 nsew signal input
rlabel metal2 s 19890 130344 19946 131144 6 io_in[10]
port 82 nsew signal input
rlabel metal2 s 21822 130344 21878 131144 6 io_in[11]
port 83 nsew signal input
rlabel metal2 s 23846 130344 23902 131144 6 io_in[12]
port 84 nsew signal input
rlabel metal2 s 25778 130344 25834 131144 6 io_in[13]
port 85 nsew signal input
rlabel metal2 s 27710 130344 27766 131144 6 io_in[14]
port 86 nsew signal input
rlabel metal2 s 29734 130344 29790 131144 6 io_in[15]
port 87 nsew signal input
rlabel metal2 s 31666 130344 31722 131144 6 io_in[16]
port 88 nsew signal input
rlabel metal2 s 33598 130344 33654 131144 6 io_in[17]
port 89 nsew signal input
rlabel metal2 s 35622 130344 35678 131144 6 io_in[18]
port 90 nsew signal input
rlabel metal2 s 37554 130344 37610 131144 6 io_in[19]
port 91 nsew signal input
rlabel metal2 s 2226 130344 2282 131144 6 io_in[1]
port 92 nsew signal input
rlabel metal2 s 39578 130344 39634 131144 6 io_in[20]
port 93 nsew signal input
rlabel metal2 s 41510 130344 41566 131144 6 io_in[21]
port 94 nsew signal input
rlabel metal2 s 43442 130344 43498 131144 6 io_in[22]
port 95 nsew signal input
rlabel metal2 s 45466 130344 45522 131144 6 io_in[23]
port 96 nsew signal input
rlabel metal2 s 47398 130344 47454 131144 6 io_in[24]
port 97 nsew signal input
rlabel metal2 s 49330 130344 49386 131144 6 io_in[25]
port 98 nsew signal input
rlabel metal2 s 51354 130344 51410 131144 6 io_in[26]
port 99 nsew signal input
rlabel metal2 s 53286 130344 53342 131144 6 io_in[27]
port 100 nsew signal input
rlabel metal2 s 55218 130344 55274 131144 6 io_in[28]
port 101 nsew signal input
rlabel metal2 s 57242 130344 57298 131144 6 io_in[29]
port 102 nsew signal input
rlabel metal2 s 4158 130344 4214 131144 6 io_in[2]
port 103 nsew signal input
rlabel metal2 s 59174 130344 59230 131144 6 io_in[30]
port 104 nsew signal input
rlabel metal2 s 61106 130344 61162 131144 6 io_in[31]
port 105 nsew signal input
rlabel metal2 s 63130 130344 63186 131144 6 io_in[32]
port 106 nsew signal input
rlabel metal2 s 65062 130344 65118 131144 6 io_in[33]
port 107 nsew signal input
rlabel metal2 s 66994 130344 67050 131144 6 io_in[34]
port 108 nsew signal input
rlabel metal2 s 69018 130344 69074 131144 6 io_in[35]
port 109 nsew signal input
rlabel metal2 s 70950 130344 71006 131144 6 io_in[36]
port 110 nsew signal input
rlabel metal2 s 72882 130344 72938 131144 6 io_in[37]
port 111 nsew signal input
rlabel metal2 s 6182 130344 6238 131144 6 io_in[3]
port 112 nsew signal input
rlabel metal2 s 8114 130344 8170 131144 6 io_in[4]
port 113 nsew signal input
rlabel metal2 s 10046 130344 10102 131144 6 io_in[5]
port 114 nsew signal input
rlabel metal2 s 12070 130344 12126 131144 6 io_in[6]
port 115 nsew signal input
rlabel metal2 s 14002 130344 14058 131144 6 io_in[7]
port 116 nsew signal input
rlabel metal2 s 15934 130344 15990 131144 6 io_in[8]
port 117 nsew signal input
rlabel metal2 s 17958 130344 18014 131144 6 io_in[9]
port 118 nsew signal input
rlabel metal2 s 938 130344 994 131144 6 io_oeb[0]
port 119 nsew signal output
rlabel metal2 s 20534 130344 20590 131144 6 io_oeb[10]
port 120 nsew signal output
rlabel metal2 s 22466 130344 22522 131144 6 io_oeb[11]
port 121 nsew signal output
rlabel metal2 s 24490 130344 24546 131144 6 io_oeb[12]
port 122 nsew signal output
rlabel metal2 s 26422 130344 26478 131144 6 io_oeb[13]
port 123 nsew signal output
rlabel metal2 s 28446 130344 28502 131144 6 io_oeb[14]
port 124 nsew signal output
rlabel metal2 s 30378 130344 30434 131144 6 io_oeb[15]
port 125 nsew signal output
rlabel metal2 s 32310 130344 32366 131144 6 io_oeb[16]
port 126 nsew signal output
rlabel metal2 s 34334 130344 34390 131144 6 io_oeb[17]
port 127 nsew signal output
rlabel metal2 s 36266 130344 36322 131144 6 io_oeb[18]
port 128 nsew signal output
rlabel metal2 s 38198 130344 38254 131144 6 io_oeb[19]
port 129 nsew signal output
rlabel metal2 s 2870 130344 2926 131144 6 io_oeb[1]
port 130 nsew signal output
rlabel metal2 s 40222 130344 40278 131144 6 io_oeb[20]
port 131 nsew signal output
rlabel metal2 s 42154 130344 42210 131144 6 io_oeb[21]
port 132 nsew signal output
rlabel metal2 s 44086 130344 44142 131144 6 io_oeb[22]
port 133 nsew signal output
rlabel metal2 s 46110 130344 46166 131144 6 io_oeb[23]
port 134 nsew signal output
rlabel metal2 s 48042 130344 48098 131144 6 io_oeb[24]
port 135 nsew signal output
rlabel metal2 s 49974 130344 50030 131144 6 io_oeb[25]
port 136 nsew signal output
rlabel metal2 s 51998 130344 52054 131144 6 io_oeb[26]
port 137 nsew signal output
rlabel metal2 s 53930 130344 53986 131144 6 io_oeb[27]
port 138 nsew signal output
rlabel metal2 s 55862 130344 55918 131144 6 io_oeb[28]
port 139 nsew signal output
rlabel metal2 s 57886 130344 57942 131144 6 io_oeb[29]
port 140 nsew signal output
rlabel metal2 s 4802 130344 4858 131144 6 io_oeb[2]
port 141 nsew signal output
rlabel metal2 s 59818 130344 59874 131144 6 io_oeb[30]
port 142 nsew signal output
rlabel metal2 s 61750 130344 61806 131144 6 io_oeb[31]
port 143 nsew signal output
rlabel metal2 s 63774 130344 63830 131144 6 io_oeb[32]
port 144 nsew signal output
rlabel metal2 s 65706 130344 65762 131144 6 io_oeb[33]
port 145 nsew signal output
rlabel metal2 s 67730 130344 67786 131144 6 io_oeb[34]
port 146 nsew signal output
rlabel metal2 s 69662 130344 69718 131144 6 io_oeb[35]
port 147 nsew signal output
rlabel metal2 s 71594 130344 71650 131144 6 io_oeb[36]
port 148 nsew signal output
rlabel metal2 s 73618 130344 73674 131144 6 io_oeb[37]
port 149 nsew signal output
rlabel metal2 s 6826 130344 6882 131144 6 io_oeb[3]
port 150 nsew signal output
rlabel metal2 s 8758 130344 8814 131144 6 io_oeb[4]
port 151 nsew signal output
rlabel metal2 s 10690 130344 10746 131144 6 io_oeb[5]
port 152 nsew signal output
rlabel metal2 s 12714 130344 12770 131144 6 io_oeb[6]
port 153 nsew signal output
rlabel metal2 s 14646 130344 14702 131144 6 io_oeb[7]
port 154 nsew signal output
rlabel metal2 s 16578 130344 16634 131144 6 io_oeb[8]
port 155 nsew signal output
rlabel metal2 s 18602 130344 18658 131144 6 io_oeb[9]
port 156 nsew signal output
rlabel metal2 s 1582 130344 1638 131144 6 io_out[0]
port 157 nsew signal output
rlabel metal2 s 21178 130344 21234 131144 6 io_out[10]
port 158 nsew signal output
rlabel metal2 s 23202 130344 23258 131144 6 io_out[11]
port 159 nsew signal output
rlabel metal2 s 25134 130344 25190 131144 6 io_out[12]
port 160 nsew signal output
rlabel metal2 s 27066 130344 27122 131144 6 io_out[13]
port 161 nsew signal output
rlabel metal2 s 29090 130344 29146 131144 6 io_out[14]
port 162 nsew signal output
rlabel metal2 s 31022 130344 31078 131144 6 io_out[15]
port 163 nsew signal output
rlabel metal2 s 32954 130344 33010 131144 6 io_out[16]
port 164 nsew signal output
rlabel metal2 s 34978 130344 35034 131144 6 io_out[17]
port 165 nsew signal output
rlabel metal2 s 36910 130344 36966 131144 6 io_out[18]
port 166 nsew signal output
rlabel metal2 s 38842 130344 38898 131144 6 io_out[19]
port 167 nsew signal output
rlabel metal2 s 3514 130344 3570 131144 6 io_out[1]
port 168 nsew signal output
rlabel metal2 s 40866 130344 40922 131144 6 io_out[20]
port 169 nsew signal output
rlabel metal2 s 42798 130344 42854 131144 6 io_out[21]
port 170 nsew signal output
rlabel metal2 s 44730 130344 44786 131144 6 io_out[22]
port 171 nsew signal output
rlabel metal2 s 46754 130344 46810 131144 6 io_out[23]
port 172 nsew signal output
rlabel metal2 s 48686 130344 48742 131144 6 io_out[24]
port 173 nsew signal output
rlabel metal2 s 50618 130344 50674 131144 6 io_out[25]
port 174 nsew signal output
rlabel metal2 s 52642 130344 52698 131144 6 io_out[26]
port 175 nsew signal output
rlabel metal2 s 54574 130344 54630 131144 6 io_out[27]
port 176 nsew signal output
rlabel metal2 s 56598 130344 56654 131144 6 io_out[28]
port 177 nsew signal output
rlabel metal2 s 58530 130344 58586 131144 6 io_out[29]
port 178 nsew signal output
rlabel metal2 s 5446 130344 5502 131144 6 io_out[2]
port 179 nsew signal output
rlabel metal2 s 60462 130344 60518 131144 6 io_out[30]
port 180 nsew signal output
rlabel metal2 s 62486 130344 62542 131144 6 io_out[31]
port 181 nsew signal output
rlabel metal2 s 64418 130344 64474 131144 6 io_out[32]
port 182 nsew signal output
rlabel metal2 s 66350 130344 66406 131144 6 io_out[33]
port 183 nsew signal output
rlabel metal2 s 68374 130344 68430 131144 6 io_out[34]
port 184 nsew signal output
rlabel metal2 s 70306 130344 70362 131144 6 io_out[35]
port 185 nsew signal output
rlabel metal2 s 72238 130344 72294 131144 6 io_out[36]
port 186 nsew signal output
rlabel metal2 s 74262 130344 74318 131144 6 io_out[37]
port 187 nsew signal output
rlabel metal2 s 7470 130344 7526 131144 6 io_out[3]
port 188 nsew signal output
rlabel metal2 s 9402 130344 9458 131144 6 io_out[4]
port 189 nsew signal output
rlabel metal2 s 11334 130344 11390 131144 6 io_out[5]
port 190 nsew signal output
rlabel metal2 s 13358 130344 13414 131144 6 io_out[6]
port 191 nsew signal output
rlabel metal2 s 15290 130344 15346 131144 6 io_out[7]
port 192 nsew signal output
rlabel metal2 s 17314 130344 17370 131144 6 io_out[8]
port 193 nsew signal output
rlabel metal2 s 19246 130344 19302 131144 6 io_out[9]
port 194 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 iram_addr0[0]
port 195 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 iram_addr0[1]
port 196 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 iram_addr0[2]
port 197 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 iram_addr0[3]
port 198 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 iram_addr0[4]
port 199 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 iram_addr0[5]
port 200 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 iram_addr0[6]
port 201 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 iram_addr0[7]
port 202 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 iram_addr0[8]
port 203 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 iram_clk0
port 204 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 iram_csb0
port 205 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 iram_din0[0]
port 206 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 iram_din0[10]
port 207 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 iram_din0[11]
port 208 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 iram_din0[12]
port 209 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 iram_din0[13]
port 210 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 iram_din0[14]
port 211 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 iram_din0[15]
port 212 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 iram_din0[16]
port 213 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 iram_din0[17]
port 214 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 iram_din0[18]
port 215 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 iram_din0[19]
port 216 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 iram_din0[1]
port 217 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 iram_din0[20]
port 218 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 iram_din0[21]
port 219 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 iram_din0[22]
port 220 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 iram_din0[23]
port 221 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 iram_din0[24]
port 222 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 iram_din0[25]
port 223 nsew signal output
rlabel metal2 s 126794 0 126850 800 6 iram_din0[26]
port 224 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 iram_din0[27]
port 225 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 iram_din0[28]
port 226 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 iram_din0[29]
port 227 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 iram_din0[2]
port 228 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 iram_din0[30]
port 229 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 iram_din0[31]
port 230 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 iram_din0[3]
port 231 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 iram_din0[4]
port 232 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 iram_din0[5]
port 233 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 iram_din0[6]
port 234 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 iram_din0[7]
port 235 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 iram_din0[8]
port 236 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 iram_din0[9]
port 237 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 iram_dout0[0]
port 238 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 iram_dout0[10]
port 239 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 iram_dout0[11]
port 240 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 iram_dout0[12]
port 241 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 iram_dout0[13]
port 242 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 iram_dout0[14]
port 243 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 iram_dout0[15]
port 244 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 iram_dout0[16]
port 245 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 iram_dout0[17]
port 246 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 iram_dout0[18]
port 247 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 iram_dout0[19]
port 248 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 iram_dout0[1]
port 249 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 iram_dout0[20]
port 250 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 iram_dout0[21]
port 251 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 iram_dout0[22]
port 252 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 iram_dout0[23]
port 253 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 iram_dout0[24]
port 254 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 iram_dout0[25]
port 255 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 iram_dout0[26]
port 256 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 iram_dout0[27]
port 257 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 iram_dout0[28]
port 258 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 iram_dout0[29]
port 259 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 iram_dout0[2]
port 260 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 iram_dout0[30]
port 261 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 iram_dout0[31]
port 262 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 iram_dout0[3]
port 263 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 iram_dout0[4]
port 264 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 iram_dout0[5]
port 265 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 iram_dout0[6]
port 266 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 iram_dout0[7]
port 267 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 iram_dout0[8]
port 268 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 iram_dout0[9]
port 269 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 iram_web0
port 270 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 iram_wmask0[0]
port 271 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 iram_wmask0[1]
port 272 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 iram_wmask0[2]
port 273 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 iram_wmask0[3]
port 274 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_in[0]
port 275 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[100]
port 276 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[101]
port 277 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[102]
port 278 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[103]
port 279 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[104]
port 280 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[105]
port 281 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[106]
port 282 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[107]
port 283 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[108]
port 284 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_data_in[109]
port 285 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[10]
port 286 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[110]
port 287 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[111]
port 288 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[112]
port 289 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[113]
port 290 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[114]
port 291 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[115]
port 292 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[116]
port 293 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[117]
port 294 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[118]
port 295 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[119]
port 296 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[11]
port 297 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[120]
port 298 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[121]
port 299 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[122]
port 300 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[123]
port 301 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[124]
port 302 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[125]
port 303 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[126]
port 304 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[127]
port 305 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_data_in[12]
port 306 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[13]
port 307 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[14]
port 308 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[15]
port 309 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[16]
port 310 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[17]
port 311 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[18]
port 312 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[19]
port 313 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[1]
port 314 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[20]
port 315 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[21]
port 316 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[22]
port 317 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[23]
port 318 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[24]
port 319 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_data_in[25]
port 320 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[26]
port 321 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_data_in[27]
port 322 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[28]
port 323 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[29]
port 324 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[2]
port 325 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[30]
port 326 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[31]
port 327 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[32]
port 328 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[33]
port 329 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[34]
port 330 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[35]
port 331 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_data_in[36]
port 332 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[37]
port 333 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[38]
port 334 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[39]
port 335 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[3]
port 336 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[40]
port 337 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[41]
port 338 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[42]
port 339 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[43]
port 340 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[44]
port 341 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[45]
port 342 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[46]
port 343 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[47]
port 344 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[48]
port 345 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[49]
port 346 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[4]
port 347 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_data_in[50]
port 348 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[51]
port 349 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[52]
port 350 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[53]
port 351 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[54]
port 352 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[55]
port 353 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[56]
port 354 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[57]
port 355 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[58]
port 356 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[59]
port 357 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[5]
port 358 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[60]
port 359 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[61]
port 360 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[62]
port 361 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[63]
port 362 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[64]
port 363 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[65]
port 364 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[66]
port 365 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[67]
port 366 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[68]
port 367 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[69]
port 368 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_data_in[6]
port 369 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[70]
port 370 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[71]
port 371 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[72]
port 372 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[73]
port 373 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[74]
port 374 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[75]
port 375 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[76]
port 376 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[77]
port 377 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[78]
port 378 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[79]
port 379 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[7]
port 380 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[80]
port 381 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[81]
port 382 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[82]
port 383 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[83]
port 384 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[84]
port 385 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[85]
port 386 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[86]
port 387 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[87]
port 388 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[88]
port 389 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[89]
port 390 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[8]
port 391 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[90]
port 392 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[91]
port 393 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[92]
port 394 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[93]
port 395 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[94]
port 396 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[95]
port 397 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[96]
port 398 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[97]
port 399 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[98]
port 400 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[99]
port 401 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[9]
port 402 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_out[0]
port 403 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[100]
port 404 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[101]
port 405 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[102]
port 406 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 la_data_out[103]
port 407 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[104]
port 408 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[105]
port 409 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[106]
port 410 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[107]
port 411 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[108]
port 412 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[109]
port 413 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[10]
port 414 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[110]
port 415 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[111]
port 416 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 la_data_out[112]
port 417 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[113]
port 418 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[114]
port 419 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[115]
port 420 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[116]
port 421 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 la_data_out[117]
port 422 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[118]
port 423 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[119]
port 424 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[11]
port 425 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 la_data_out[120]
port 426 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[121]
port 427 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[122]
port 428 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[123]
port 429 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[124]
port 430 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[125]
port 431 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[126]
port 432 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[127]
port 433 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[12]
port 434 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[13]
port 435 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[14]
port 436 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[15]
port 437 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[16]
port 438 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[17]
port 439 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[18]
port 440 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[19]
port 441 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[1]
port 442 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[20]
port 443 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[21]
port 444 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[22]
port 445 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[23]
port 446 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[24]
port 447 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[25]
port 448 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 la_data_out[26]
port 449 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 la_data_out[27]
port 450 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[28]
port 451 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[29]
port 452 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[2]
port 453 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[30]
port 454 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[31]
port 455 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[32]
port 456 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[33]
port 457 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[34]
port 458 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[35]
port 459 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[36]
port 460 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[37]
port 461 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[38]
port 462 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[39]
port 463 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[3]
port 464 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[40]
port 465 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[41]
port 466 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[42]
port 467 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[43]
port 468 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[44]
port 469 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[45]
port 470 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[46]
port 471 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[47]
port 472 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[48]
port 473 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[49]
port 474 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[4]
port 475 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[50]
port 476 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[51]
port 477 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[52]
port 478 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[53]
port 479 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[54]
port 480 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[55]
port 481 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[56]
port 482 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[57]
port 483 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[58]
port 484 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[59]
port 485 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[5]
port 486 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[60]
port 487 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[61]
port 488 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[62]
port 489 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[63]
port 490 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[64]
port 491 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[65]
port 492 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[66]
port 493 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[67]
port 494 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[68]
port 495 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[69]
port 496 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[6]
port 497 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[70]
port 498 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[71]
port 499 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[72]
port 500 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[73]
port 501 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[74]
port 502 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[75]
port 503 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[76]
port 504 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[77]
port 505 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[78]
port 506 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[79]
port 507 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[7]
port 508 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[80]
port 509 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[81]
port 510 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[82]
port 511 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[83]
port 512 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[84]
port 513 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[85]
port 514 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[86]
port 515 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[87]
port 516 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[88]
port 517 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[89]
port 518 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[8]
port 519 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[90]
port 520 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[91]
port 521 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[92]
port 522 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[93]
port 523 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[94]
port 524 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[95]
port 525 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[96]
port 526 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[97]
port 527 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[98]
port 528 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[99]
port 529 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[9]
port 530 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_oenb[0]
port 531 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[100]
port 532 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_oenb[101]
port 533 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[102]
port 534 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[103]
port 535 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[104]
port 536 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_oenb[105]
port 537 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[106]
port 538 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_oenb[107]
port 539 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[108]
port 540 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[109]
port 541 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[10]
port 542 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[110]
port 543 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[111]
port 544 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[112]
port 545 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_oenb[113]
port 546 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[114]
port 547 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[115]
port 548 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[116]
port 549 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[117]
port 550 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[118]
port 551 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_oenb[119]
port 552 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[11]
port 553 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[120]
port 554 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[121]
port 555 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_oenb[122]
port 556 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[123]
port 557 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[124]
port 558 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[125]
port 559 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_oenb[126]
port 560 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[127]
port 561 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[12]
port 562 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[13]
port 563 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[14]
port 564 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_oenb[15]
port 565 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[16]
port 566 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[17]
port 567 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[18]
port 568 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[19]
port 569 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[1]
port 570 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[20]
port 571 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[21]
port 572 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[22]
port 573 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[23]
port 574 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_oenb[24]
port 575 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[25]
port 576 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[26]
port 577 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[27]
port 578 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[28]
port 579 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[29]
port 580 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[2]
port 581 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[30]
port 582 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[31]
port 583 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[32]
port 584 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[33]
port 585 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_oenb[34]
port 586 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[35]
port 587 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[36]
port 588 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[37]
port 589 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[38]
port 590 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[39]
port 591 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[3]
port 592 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[40]
port 593 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[41]
port 594 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[42]
port 595 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_oenb[43]
port 596 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[44]
port 597 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[45]
port 598 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[46]
port 599 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[47]
port 600 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[48]
port 601 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[49]
port 602 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[4]
port 603 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[50]
port 604 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[51]
port 605 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[52]
port 606 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[53]
port 607 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[54]
port 608 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[55]
port 609 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[56]
port 610 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[57]
port 611 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[58]
port 612 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[59]
port 613 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[5]
port 614 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_oenb[60]
port 615 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[61]
port 616 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[62]
port 617 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[63]
port 618 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[64]
port 619 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[65]
port 620 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[66]
port 621 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[67]
port 622 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[68]
port 623 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[69]
port 624 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[6]
port 625 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[70]
port 626 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[71]
port 627 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[72]
port 628 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[73]
port 629 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[74]
port 630 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[75]
port 631 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[76]
port 632 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[77]
port 633 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oenb[78]
port 634 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[79]
port 635 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[7]
port 636 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[80]
port 637 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[81]
port 638 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[82]
port 639 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[83]
port 640 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[84]
port 641 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[85]
port 642 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[86]
port 643 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[87]
port 644 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[88]
port 645 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_oenb[89]
port 646 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[8]
port 647 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[90]
port 648 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[91]
port 649 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[92]
port 650 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[93]
port 651 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[94]
port 652 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[95]
port 653 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[96]
port 654 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[97]
port 655 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[98]
port 656 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[99]
port 657 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[9]
port 658 nsew signal input
rlabel metal2 s 127254 130344 127310 131144 6 user_irq[0]
port 659 nsew signal output
rlabel metal2 s 127898 130344 127954 131144 6 user_irq[1]
port 660 nsew signal output
rlabel metal2 s 128542 130344 128598 131144 6 user_irq[2]
port 661 nsew signal output
rlabel metal4 s 4208 2128 4528 128976 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 128976 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 128976 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 128976 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 128976 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 128976 6 vssd1
port 663 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 128976 6 vssd1
port 663 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 128976 6 vssd1
port 663 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 128976 6 vssd1
port 663 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 664 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 665 nsew signal input
rlabel metal2 s 478 0 534 800 6 wb_uart_ack
port 666 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wb_uart_adr[0]
port 667 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wb_uart_adr[10]
port 668 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wb_uart_adr[11]
port 669 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wb_uart_adr[12]
port 670 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wb_uart_adr[13]
port 671 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wb_uart_adr[14]
port 672 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wb_uart_adr[15]
port 673 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wb_uart_adr[16]
port 674 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wb_uart_adr[17]
port 675 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wb_uart_adr[18]
port 676 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wb_uart_adr[19]
port 677 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 wb_uart_adr[1]
port 678 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wb_uart_adr[20]
port 679 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wb_uart_adr[21]
port 680 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 wb_uart_adr[22]
port 681 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wb_uart_adr[23]
port 682 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wb_uart_adr[24]
port 683 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wb_uart_adr[25]
port 684 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wb_uart_adr[26]
port 685 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wb_uart_adr[27]
port 686 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wb_uart_adr[28]
port 687 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wb_uart_adr[29]
port 688 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 wb_uart_adr[2]
port 689 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wb_uart_adr[30]
port 690 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wb_uart_adr[31]
port 691 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wb_uart_adr[3]
port 692 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wb_uart_adr[4]
port 693 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wb_uart_adr[5]
port 694 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wb_uart_adr[6]
port 695 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wb_uart_adr[7]
port 696 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wb_uart_adr[8]
port 697 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wb_uart_adr[9]
port 698 nsew signal output
rlabel metal2 s 662 0 718 800 6 wb_uart_clk
port 699 nsew signal output
rlabel metal2 s 846 0 902 800 6 wb_uart_cyc
port 700 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 wb_uart_dat_fromcpu[0]
port 701 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wb_uart_dat_fromcpu[10]
port 702 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wb_uart_dat_fromcpu[11]
port 703 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 wb_uart_dat_fromcpu[12]
port 704 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wb_uart_dat_fromcpu[13]
port 705 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wb_uart_dat_fromcpu[14]
port 706 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wb_uart_dat_fromcpu[15]
port 707 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wb_uart_dat_fromcpu[16]
port 708 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wb_uart_dat_fromcpu[17]
port 709 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wb_uart_dat_fromcpu[18]
port 710 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wb_uart_dat_fromcpu[19]
port 711 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wb_uart_dat_fromcpu[1]
port 712 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wb_uart_dat_fromcpu[20]
port 713 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wb_uart_dat_fromcpu[21]
port 714 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 wb_uart_dat_fromcpu[22]
port 715 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wb_uart_dat_fromcpu[23]
port 716 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wb_uart_dat_fromcpu[24]
port 717 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wb_uart_dat_fromcpu[25]
port 718 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wb_uart_dat_fromcpu[26]
port 719 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wb_uart_dat_fromcpu[27]
port 720 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wb_uart_dat_fromcpu[28]
port 721 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wb_uart_dat_fromcpu[29]
port 722 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wb_uart_dat_fromcpu[2]
port 723 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wb_uart_dat_fromcpu[30]
port 724 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wb_uart_dat_fromcpu[31]
port 725 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wb_uart_dat_fromcpu[3]
port 726 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wb_uart_dat_fromcpu[4]
port 727 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 wb_uart_dat_fromcpu[5]
port 728 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wb_uart_dat_fromcpu[6]
port 729 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wb_uart_dat_fromcpu[7]
port 730 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wb_uart_dat_fromcpu[8]
port 731 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wb_uart_dat_fromcpu[9]
port 732 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wb_uart_dat_tocpu[0]
port 733 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wb_uart_dat_tocpu[10]
port 734 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wb_uart_dat_tocpu[11]
port 735 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wb_uart_dat_tocpu[12]
port 736 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wb_uart_dat_tocpu[13]
port 737 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wb_uart_dat_tocpu[14]
port 738 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wb_uart_dat_tocpu[15]
port 739 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wb_uart_dat_tocpu[16]
port 740 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wb_uart_dat_tocpu[17]
port 741 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wb_uart_dat_tocpu[18]
port 742 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wb_uart_dat_tocpu[19]
port 743 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wb_uart_dat_tocpu[1]
port 744 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wb_uart_dat_tocpu[20]
port 745 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wb_uart_dat_tocpu[21]
port 746 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wb_uart_dat_tocpu[22]
port 747 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wb_uart_dat_tocpu[23]
port 748 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wb_uart_dat_tocpu[24]
port 749 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb_uart_dat_tocpu[25]
port 750 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wb_uart_dat_tocpu[26]
port 751 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wb_uart_dat_tocpu[27]
port 752 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wb_uart_dat_tocpu[28]
port 753 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wb_uart_dat_tocpu[29]
port 754 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wb_uart_dat_tocpu[2]
port 755 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wb_uart_dat_tocpu[30]
port 756 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wb_uart_dat_tocpu[31]
port 757 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wb_uart_dat_tocpu[3]
port 758 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wb_uart_dat_tocpu[4]
port 759 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wb_uart_dat_tocpu[5]
port 760 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wb_uart_dat_tocpu[6]
port 761 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wb_uart_dat_tocpu[7]
port 762 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_uart_dat_tocpu[8]
port 763 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wb_uart_dat_tocpu[9]
port 764 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wb_uart_rst
port 765 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wb_uart_sel[0]
port 766 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wb_uart_sel[1]
port 767 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wb_uart_sel[2]
port 768 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wb_uart_sel[3]
port 769 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wb_uart_stb
port 770 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wb_uart_we
port 771 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_ack_o
port 772 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[0]
port 773 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[10]
port 774 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[11]
port 775 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[12]
port 776 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[13]
port 777 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_adr_i[14]
port 778 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[15]
port 779 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[16]
port 780 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[17]
port 781 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[18]
port 782 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[19]
port 783 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[1]
port 784 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[20]
port 785 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[21]
port 786 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[22]
port 787 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[23]
port 788 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[24]
port 789 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[25]
port 790 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_adr_i[26]
port 791 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[27]
port 792 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[28]
port 793 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_adr_i[29]
port 794 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[2]
port 795 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[30]
port 796 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[31]
port 797 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[3]
port 798 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[4]
port 799 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[5]
port 800 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[6]
port 801 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[7]
port 802 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[8]
port 803 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[9]
port 804 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_cyc_i
port 805 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[0]
port 806 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[10]
port 807 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[11]
port 808 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[12]
port 809 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[13]
port 810 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[14]
port 811 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[15]
port 812 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[16]
port 813 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[17]
port 814 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[18]
port 815 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[19]
port 816 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[1]
port 817 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[20]
port 818 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_i[21]
port 819 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[22]
port 820 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[23]
port 821 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[24]
port 822 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_i[25]
port 823 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_i[26]
port 824 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[27]
port 825 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_i[28]
port 826 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_i[29]
port 827 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[2]
port 828 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_i[30]
port 829 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[31]
port 830 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[3]
port 831 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[4]
port 832 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[5]
port 833 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[6]
port 834 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[7]
port 835 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[8]
port 836 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[9]
port 837 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[0]
port 838 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[10]
port 839 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[11]
port 840 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[12]
port 841 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_o[13]
port 842 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[14]
port 843 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[15]
port 844 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[16]
port 845 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[17]
port 846 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[18]
port 847 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_o[19]
port 848 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[1]
port 849 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[20]
port 850 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[21]
port 851 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_o[22]
port 852 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[23]
port 853 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_o[24]
port 854 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[25]
port 855 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[26]
port 856 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[27]
port 857 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[28]
port 858 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[29]
port 859 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[2]
port 860 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_o[30]
port 861 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[31]
port 862 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[3]
port 863 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[4]
port 864 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[5]
port 865 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[6]
port 866 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_o[7]
port 867 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[8]
port 868 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[9]
port 869 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_sel_i[0]
port 870 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_sel_i[1]
port 871 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_sel_i[2]
port 872 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_sel_i[3]
port 873 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_stb_i
port 874 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_we_i
port 875 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 129000 131144
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 42944248
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/rvj1_caravel_soc/runs/rvj1_caravel_soc/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1315266
<< end >>

