magic
tech sky130A
magscale 1 2
timestamp 1654189623
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 348786 700476 348792 700528
rect 348844 700516 348850 700528
rect 357526 700516 357532 700528
rect 348844 700488 357532 700516
rect 348844 700476 348850 700488
rect 357526 700476 357532 700488
rect 357584 700476 357590 700528
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 358906 700448 358912 700460
rect 300176 700420 358912 700448
rect 300176 700408 300182 700420
rect 358906 700408 358912 700420
rect 358964 700408 358970 700460
rect 361022 700408 361028 700460
rect 361080 700448 361086 700460
rect 397454 700448 397460 700460
rect 361080 700420 397460 700448
rect 361080 700408 361086 700420
rect 397454 700408 397460 700420
rect 397512 700408 397518 700460
rect 283834 700340 283840 700392
rect 283892 700380 283898 700392
rect 357434 700380 357440 700392
rect 283892 700352 357440 700380
rect 283892 700340 283898 700352
rect 357434 700340 357440 700352
rect 357492 700340 357498 700392
rect 360930 700340 360936 700392
rect 360988 700380 360994 700392
rect 429838 700380 429844 700392
rect 360988 700352 429844 700380
rect 360988 700340 360994 700352
rect 429838 700340 429844 700352
rect 429896 700340 429902 700392
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 358814 700312 358820 700324
rect 267700 700284 358820 700312
rect 267700 700272 267706 700284
rect 358814 700272 358820 700284
rect 358872 700272 358878 700324
rect 360838 700272 360844 700324
rect 360896 700312 360902 700324
rect 559650 700312 559656 700324
rect 360896 700284 559656 700312
rect 360896 700272 360902 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 362218 696940 362224 696992
rect 362276 696980 362282 696992
rect 580166 696980 580172 696992
rect 362276 696952 580172 696980
rect 362276 696940 362282 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 359458 670692 359464 670744
rect 359516 670732 359522 670744
rect 580166 670732 580172 670744
rect 359516 670704 580172 670732
rect 359516 670692 359522 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 2774 656956 2780 657008
rect 2832 656996 2838 657008
rect 4890 656996 4896 657008
rect 2832 656968 4896 656996
rect 2832 656956 2838 656968
rect 4890 656956 4896 656968
rect 4948 656956 4954 657008
rect 361114 643084 361120 643136
rect 361172 643124 361178 643136
rect 580166 643124 580172 643136
rect 361172 643096 580172 643124
rect 361172 643084 361178 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4982 632108 4988 632120
rect 2832 632080 4988 632108
rect 2832 632068 2838 632080
rect 4982 632068 4988 632080
rect 5040 632068 5046 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 32398 618304 32404 618316
rect 3568 618276 32404 618304
rect 3568 618264 3574 618276
rect 32398 618264 32404 618276
rect 32456 618264 32462 618316
rect 358078 616836 358084 616888
rect 358136 616876 358142 616888
rect 580166 616876 580172 616888
rect 358136 616848 580172 616876
rect 358136 616836 358142 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 10318 605860 10324 605872
rect 3568 605832 10324 605860
rect 3568 605820 3574 605832
rect 10318 605820 10324 605832
rect 10376 605820 10382 605872
rect 3510 579776 3516 579828
rect 3568 579816 3574 579828
rect 8938 579816 8944 579828
rect 3568 579788 8944 579816
rect 3568 579776 3574 579788
rect 8938 579776 8944 579788
rect 8996 579776 9002 579828
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 84838 565876 84844 565888
rect 3292 565848 84844 565876
rect 3292 565836 3298 565848
rect 84838 565836 84844 565848
rect 84896 565836 84902 565888
rect 217962 565088 217968 565140
rect 218020 565128 218026 565140
rect 234614 565128 234620 565140
rect 218020 565100 234620 565128
rect 218020 565088 218026 565100
rect 234614 565088 234620 565100
rect 234672 565088 234678 565140
rect 331214 565088 331220 565140
rect 331272 565128 331278 565140
rect 358998 565128 359004 565140
rect 331272 565100 359004 565128
rect 331272 565088 331278 565100
rect 358998 565088 359004 565100
rect 359056 565088 359062 565140
rect 371878 563048 371884 563100
rect 371936 563088 371942 563100
rect 579798 563088 579804 563100
rect 371936 563060 579804 563088
rect 371936 563048 371942 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 2774 553664 2780 553716
rect 2832 553704 2838 553716
rect 5074 553704 5080 553716
rect 2832 553676 5080 553704
rect 2832 553664 2838 553676
rect 5074 553664 5080 553676
rect 5132 553664 5138 553716
rect 358170 536800 358176 536852
rect 358228 536840 358234 536852
rect 579614 536840 579620 536852
rect 358228 536812 579620 536840
rect 358228 536800 358234 536812
rect 579614 536800 579620 536812
rect 579672 536800 579678 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 10410 527184 10416 527196
rect 3016 527156 10416 527184
rect 3016 527144 3022 527156
rect 10410 527144 10416 527156
rect 10468 527144 10474 527196
rect 358262 484372 358268 484424
rect 358320 484412 358326 484424
rect 580166 484412 580172 484424
rect 358320 484384 580172 484412
rect 358320 484372 358326 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 219066 478184 219072 478236
rect 219124 478224 219130 478236
rect 248414 478224 248420 478236
rect 219124 478196 248420 478224
rect 219124 478184 219130 478196
rect 248414 478184 248420 478196
rect 248472 478184 248478 478236
rect 217686 478116 217692 478168
rect 217744 478156 217750 478168
rect 251174 478156 251180 478168
rect 217744 478128 251180 478156
rect 217744 478116 217750 478128
rect 251174 478116 251180 478128
rect 251232 478116 251238 478168
rect 311894 478116 311900 478168
rect 311952 478156 311958 478168
rect 357526 478156 357532 478168
rect 311952 478128 357532 478156
rect 311952 478116 311958 478128
rect 357526 478116 357532 478128
rect 357584 478116 357590 478168
rect 258350 476688 258356 476740
rect 258408 476728 258414 476740
rect 258408 476700 267734 476728
rect 258408 476688 258414 476700
rect 256602 476620 256608 476672
rect 256660 476660 256666 476672
rect 260098 476660 260104 476672
rect 256660 476632 260104 476660
rect 256660 476620 256666 476632
rect 260098 476620 260104 476632
rect 260156 476620 260162 476672
rect 241606 476552 241612 476604
rect 241664 476592 241670 476604
rect 252554 476592 252560 476604
rect 241664 476564 252560 476592
rect 241664 476552 241670 476564
rect 252554 476552 252560 476564
rect 252612 476552 252618 476604
rect 252646 476552 252652 476604
rect 252704 476592 252710 476604
rect 263594 476592 263600 476604
rect 252704 476564 263600 476592
rect 252704 476552 252710 476564
rect 263594 476552 263600 476564
rect 263652 476552 263658 476604
rect 247034 476524 247040 476536
rect 238726 476496 247040 476524
rect 236086 476416 236092 476468
rect 236144 476456 236150 476468
rect 238726 476456 238754 476496
rect 247034 476484 247040 476496
rect 247092 476484 247098 476536
rect 249794 476524 249800 476536
rect 248386 476496 249800 476524
rect 236144 476428 238754 476456
rect 236144 476416 236150 476428
rect 238846 476416 238852 476468
rect 238904 476456 238910 476468
rect 244274 476456 244280 476468
rect 238904 476428 244280 476456
rect 238904 476416 238910 476428
rect 244274 476416 244280 476428
rect 244332 476416 244338 476468
rect 248386 476456 248414 476496
rect 249794 476484 249800 476496
rect 249852 476484 249858 476536
rect 255314 476484 255320 476536
rect 255372 476524 255378 476536
rect 264974 476524 264980 476536
rect 255372 476496 264980 476524
rect 255372 476484 255378 476496
rect 264974 476484 264980 476496
rect 265032 476484 265038 476536
rect 244384 476428 248414 476456
rect 238754 476348 238760 476400
rect 238812 476388 238818 476400
rect 244384 476388 244412 476428
rect 253842 476416 253848 476468
rect 253900 476456 253906 476468
rect 258074 476456 258080 476468
rect 253900 476428 258080 476456
rect 253900 476416 253906 476428
rect 258074 476416 258080 476428
rect 258132 476416 258138 476468
rect 259546 476416 259552 476468
rect 259604 476456 259610 476468
rect 267706 476456 267734 476700
rect 278774 476688 278780 476740
rect 278832 476728 278838 476740
rect 302234 476728 302240 476740
rect 278832 476700 302240 476728
rect 278832 476688 278838 476700
rect 302234 476688 302240 476700
rect 302292 476688 302298 476740
rect 280338 476620 280344 476672
rect 280396 476660 280402 476672
rect 304994 476660 305000 476672
rect 280396 476632 305000 476660
rect 280396 476620 280402 476632
rect 304994 476620 305000 476632
rect 305052 476620 305058 476672
rect 284294 476552 284300 476604
rect 284352 476592 284358 476604
rect 310514 476592 310520 476604
rect 284352 476564 310520 476592
rect 284352 476552 284358 476564
rect 310514 476552 310520 476564
rect 310572 476552 310578 476604
rect 281534 476484 281540 476536
rect 281592 476524 281598 476536
rect 307754 476524 307760 476536
rect 281592 476496 307760 476524
rect 281592 476484 281598 476496
rect 307754 476484 307760 476496
rect 307812 476484 307818 476536
rect 267826 476456 267832 476468
rect 259604 476428 265848 476456
rect 267706 476428 267832 476456
rect 259604 476416 259610 476428
rect 238812 476360 244412 476388
rect 238812 476348 238818 476360
rect 245746 476348 245752 476400
rect 245804 476388 245810 476400
rect 255406 476388 255412 476400
rect 245804 476360 255412 476388
rect 245804 476348 245810 476360
rect 255406 476348 255412 476360
rect 255464 476348 255470 476400
rect 260926 476348 260932 476400
rect 260984 476388 260990 476400
rect 265820 476388 265848 476428
rect 267826 476416 267832 476428
rect 267884 476416 267890 476468
rect 285674 476416 285680 476468
rect 285732 476456 285738 476468
rect 313274 476456 313280 476468
rect 285732 476428 313280 476456
rect 285732 476416 285738 476428
rect 313274 476416 313280 476428
rect 313332 476416 313338 476468
rect 270494 476388 270500 476400
rect 260984 476360 265756 476388
rect 265820 476360 270500 476388
rect 260984 476348 260990 476360
rect 234614 476280 234620 476332
rect 234672 476320 234678 476332
rect 242894 476320 242900 476332
rect 234672 476292 242900 476320
rect 234672 476280 234678 476292
rect 242894 476280 242900 476292
rect 242952 476280 242958 476332
rect 248506 476280 248512 476332
rect 248564 476320 248570 476332
rect 258258 476320 258264 476332
rect 248564 476292 258264 476320
rect 248564 476280 248570 476292
rect 258258 476280 258264 476292
rect 258316 476280 258322 476332
rect 260742 476280 260748 476332
rect 260800 476320 260806 476332
rect 265618 476320 265624 476332
rect 260800 476292 265624 476320
rect 260800 476280 260806 476292
rect 265618 476280 265624 476292
rect 265676 476280 265682 476332
rect 265728 476320 265756 476360
rect 270494 476348 270500 476360
rect 270552 476348 270558 476400
rect 287054 476348 287060 476400
rect 287112 476388 287118 476400
rect 314654 476388 314660 476400
rect 287112 476360 314660 476388
rect 287112 476348 287118 476360
rect 314654 476348 314660 476360
rect 314712 476348 314718 476400
rect 273254 476320 273260 476332
rect 265728 476292 273260 476320
rect 273254 476280 273260 476292
rect 273312 476280 273318 476332
rect 288434 476280 288440 476332
rect 288492 476320 288498 476332
rect 317414 476320 317420 476332
rect 288492 476292 317420 476320
rect 288492 476280 288498 476292
rect 317414 476280 317420 476292
rect 317472 476280 317478 476332
rect 241514 476212 241520 476264
rect 241572 476252 241578 476264
rect 244274 476252 244280 476264
rect 241572 476224 244280 476252
rect 241572 476212 241578 476224
rect 244274 476212 244280 476224
rect 244332 476212 244338 476264
rect 251266 476212 251272 476264
rect 251324 476252 251330 476264
rect 260834 476252 260840 476264
rect 251324 476224 260840 476252
rect 251324 476212 251330 476224
rect 260834 476212 260840 476224
rect 260892 476212 260898 476264
rect 263686 476212 263692 476264
rect 263744 476252 263750 476264
rect 277762 476252 277768 476264
rect 263744 476224 277768 476252
rect 263744 476212 263750 476224
rect 277762 476212 277768 476224
rect 277820 476212 277826 476264
rect 289906 476212 289912 476264
rect 289964 476252 289970 476264
rect 320174 476252 320180 476264
rect 289964 476224 320180 476252
rect 289964 476212 289970 476224
rect 320174 476212 320180 476224
rect 320232 476212 320238 476264
rect 242802 476144 242808 476196
rect 242860 476184 242866 476196
rect 244918 476184 244924 476196
rect 242860 476156 244924 476184
rect 242860 476144 242866 476156
rect 244918 476144 244924 476156
rect 244976 476144 244982 476196
rect 251082 476144 251088 476196
rect 251140 476184 251146 476196
rect 252646 476184 252652 476196
rect 251140 476156 252652 476184
rect 251140 476144 251146 476156
rect 252646 476144 252652 476156
rect 252704 476144 252710 476196
rect 258166 476144 258172 476196
rect 258224 476184 258230 476196
rect 261478 476184 261484 476196
rect 258224 476156 261484 476184
rect 258224 476144 258230 476156
rect 261478 476144 261484 476156
rect 261536 476144 261542 476196
rect 262214 476144 262220 476196
rect 262272 476184 262278 476196
rect 262272 476156 262996 476184
rect 262272 476144 262278 476156
rect 234706 476076 234712 476128
rect 234764 476116 234770 476128
rect 235902 476116 235908 476128
rect 234764 476088 235908 476116
rect 234764 476076 234770 476088
rect 235902 476076 235908 476088
rect 235960 476076 235966 476128
rect 241422 476076 241428 476128
rect 241480 476116 241486 476128
rect 242894 476116 242900 476128
rect 241480 476088 242900 476116
rect 241480 476076 241486 476088
rect 242894 476076 242900 476088
rect 242952 476076 242958 476128
rect 244366 476076 244372 476128
rect 244424 476116 244430 476128
rect 245654 476116 245660 476128
rect 244424 476088 245660 476116
rect 244424 476076 244430 476088
rect 245654 476076 245660 476088
rect 245712 476076 245718 476128
rect 252370 476076 252376 476128
rect 252428 476116 252434 476128
rect 253934 476116 253940 476128
rect 252428 476088 253940 476116
rect 252428 476076 252434 476088
rect 253934 476076 253940 476088
rect 253992 476076 253998 476128
rect 260742 476076 260748 476128
rect 260800 476116 260806 476128
rect 262858 476116 262864 476128
rect 260800 476088 262864 476116
rect 260800 476076 260806 476088
rect 262858 476076 262864 476088
rect 262916 476076 262922 476128
rect 262968 476116 262996 476156
rect 265158 476144 265164 476196
rect 265216 476184 265222 476196
rect 280154 476184 280160 476196
rect 265216 476156 280160 476184
rect 265216 476144 265222 476156
rect 280154 476144 280160 476156
rect 280212 476144 280218 476196
rect 291194 476144 291200 476196
rect 291252 476184 291258 476196
rect 322934 476184 322940 476196
rect 291252 476156 322940 476184
rect 291252 476144 291258 476156
rect 322934 476144 322940 476156
rect 322992 476144 322998 476196
rect 276014 476116 276020 476128
rect 262968 476088 276020 476116
rect 276014 476076 276020 476088
rect 276072 476076 276078 476128
rect 292574 476076 292580 476128
rect 292632 476116 292638 476128
rect 325786 476116 325792 476128
rect 292632 476088 325792 476116
rect 292632 476076 292638 476088
rect 325786 476076 325792 476088
rect 325844 476076 325850 476128
rect 217318 475328 217324 475380
rect 217376 475368 217382 475380
rect 231854 475368 231860 475380
rect 217376 475340 231860 475368
rect 217376 475328 217382 475340
rect 231854 475328 231860 475340
rect 231912 475328 231918 475380
rect 273162 475328 273168 475380
rect 273220 475368 273226 475380
rect 282914 475368 282920 475380
rect 273220 475340 282920 475368
rect 273220 475328 273226 475340
rect 282914 475328 282920 475340
rect 282972 475328 282978 475380
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 332594 474756 332600 474768
rect 3108 474728 332600 474756
rect 3108 474716 3114 474728
rect 332594 474716 332600 474728
rect 332652 474716 332658 474768
rect 219158 474036 219164 474088
rect 219216 474076 219222 474088
rect 240226 474076 240232 474088
rect 219216 474048 240232 474076
rect 219216 474036 219222 474048
rect 240226 474036 240232 474048
rect 240284 474036 240290 474088
rect 3602 473968 3608 474020
rect 3660 474008 3666 474020
rect 353294 474008 353300 474020
rect 3660 473980 353300 474008
rect 3660 473968 3666 473980
rect 353294 473968 353300 473980
rect 353352 473968 353358 474020
rect 273254 471248 273260 471300
rect 273312 471288 273318 471300
rect 292666 471288 292672 471300
rect 273312 471260 292672 471288
rect 273312 471248 273318 471260
rect 292666 471248 292672 471260
rect 292724 471248 292730 471300
rect 277302 469956 277308 470008
rect 277360 469996 277366 470008
rect 289998 469996 290004 470008
rect 277360 469968 290004 469996
rect 277360 469956 277366 469968
rect 289998 469956 290004 469968
rect 290056 469956 290062 470008
rect 270402 469888 270408 469940
rect 270460 469928 270466 469940
rect 280246 469928 280252 469940
rect 270460 469900 280252 469928
rect 270460 469888 270466 469900
rect 280246 469888 280252 469900
rect 280304 469888 280310 469940
rect 271874 469820 271880 469872
rect 271932 469860 271938 469872
rect 289814 469860 289820 469872
rect 271932 469832 289820 469860
rect 271932 469820 271938 469832
rect 289814 469820 289820 469832
rect 289872 469820 289878 469872
rect 267642 468596 267648 468648
rect 267700 468636 267706 468648
rect 274634 468636 274640 468648
rect 267700 468608 274640 468636
rect 267700 468596 267706 468608
rect 274634 468596 274640 468608
rect 274692 468596 274698 468648
rect 275922 468596 275928 468648
rect 275980 468636 275986 468648
rect 287146 468636 287152 468648
rect 275980 468608 287152 468636
rect 275980 468596 275986 468608
rect 287146 468596 287152 468608
rect 287204 468596 287210 468648
rect 266262 468528 266268 468580
rect 266320 468568 266326 468580
rect 273346 468568 273352 468580
rect 266320 468540 273352 468568
rect 266320 468528 266326 468540
rect 273346 468528 273352 468540
rect 273404 468528 273410 468580
rect 274450 468528 274456 468580
rect 274508 468568 274514 468580
rect 285766 468568 285772 468580
rect 274508 468540 285772 468568
rect 274508 468528 274514 468540
rect 285766 468528 285772 468540
rect 285824 468528 285830 468580
rect 217778 468460 217784 468512
rect 217836 468500 217842 468512
rect 254026 468500 254032 468512
rect 217836 468472 254032 468500
rect 217836 468460 217842 468472
rect 254026 468460 254032 468472
rect 254084 468460 254090 468512
rect 267550 468460 267556 468512
rect 267608 468500 267614 468512
rect 277394 468500 277400 468512
rect 267608 468472 277400 468500
rect 267608 468460 267614 468472
rect 277394 468460 277400 468472
rect 277452 468460 277458 468512
rect 278682 468460 278688 468512
rect 278740 468500 278746 468512
rect 291286 468500 291292 468512
rect 278740 468472 291292 468500
rect 278740 468460 278746 468472
rect 291286 468460 291292 468472
rect 291344 468460 291350 468512
rect 262122 467780 262128 467832
rect 262180 467820 262186 467832
rect 269114 467820 269120 467832
rect 262180 467792 269120 467820
rect 262180 467780 262186 467792
rect 269114 467780 269120 467792
rect 269172 467780 269178 467832
rect 264882 467236 264888 467288
rect 264940 467276 264946 467288
rect 271966 467276 271972 467288
rect 264940 467248 271972 467276
rect 264940 467236 264946 467248
rect 271966 467236 271972 467248
rect 272024 467236 272030 467288
rect 274542 467236 274548 467288
rect 274600 467276 274606 467288
rect 284478 467276 284484 467288
rect 274600 467248 284484 467276
rect 274600 467236 274606 467248
rect 284478 467236 284484 467248
rect 284536 467236 284542 467288
rect 263502 467168 263508 467220
rect 263560 467208 263566 467220
rect 270678 467208 270684 467220
rect 263560 467180 270684 467208
rect 263560 467168 263566 467180
rect 270678 467168 270684 467180
rect 270736 467168 270742 467220
rect 271782 467168 271788 467220
rect 271840 467208 271846 467220
rect 281626 467208 281632 467220
rect 271840 467180 281632 467208
rect 271840 467168 271846 467180
rect 281626 467168 281632 467180
rect 281684 467168 281690 467220
rect 269022 467100 269028 467152
rect 269080 467140 269086 467152
rect 278866 467140 278872 467152
rect 269080 467112 278872 467140
rect 269080 467100 269086 467112
rect 278866 467100 278872 467112
rect 278924 467100 278930 467152
rect 280062 467100 280068 467152
rect 280120 467140 280126 467152
rect 292666 467140 292672 467152
rect 280120 467112 292672 467140
rect 280120 467100 280126 467112
rect 292666 467100 292672 467112
rect 292724 467100 292730 467152
rect 218054 465672 218060 465724
rect 218112 465712 218118 465724
rect 316034 465712 316040 465724
rect 218112 465684 316040 465712
rect 218112 465672 218118 465684
rect 316034 465672 316040 465684
rect 316092 465672 316098 465724
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 333974 462380 333980 462392
rect 3384 462352 333980 462380
rect 3384 462340 3390 462352
rect 333974 462340 333980 462352
rect 334032 462340 334038 462392
rect 274726 456152 274732 456204
rect 274784 456192 274790 456204
rect 295334 456192 295340 456204
rect 274784 456164 295340 456192
rect 274784 456152 274790 456164
rect 295334 456152 295340 456164
rect 295392 456152 295398 456204
rect 217594 456084 217600 456136
rect 217652 456124 217658 456136
rect 233234 456124 233240 456136
rect 217652 456096 233240 456124
rect 217652 456084 217658 456096
rect 233234 456084 233240 456096
rect 233292 456084 233298 456136
rect 276290 456084 276296 456136
rect 276348 456124 276354 456136
rect 298094 456124 298100 456136
rect 276348 456096 298100 456124
rect 276348 456084 276354 456096
rect 298094 456084 298100 456096
rect 298152 456084 298158 456136
rect 217502 456016 217508 456068
rect 217560 456056 217566 456068
rect 233326 456056 233332 456068
rect 217560 456028 233332 456056
rect 217560 456016 217566 456028
rect 233326 456016 233332 456028
rect 233384 456016 233390 456068
rect 277762 456016 277768 456068
rect 277820 456056 277826 456068
rect 300854 456056 300860 456068
rect 277820 456028 300860 456056
rect 277820 456016 277826 456028
rect 300854 456016 300860 456028
rect 300912 456016 300918 456068
rect 336826 454860 336832 454912
rect 336884 454900 336890 454912
rect 361022 454900 361028 454912
rect 336884 454872 361028 454900
rect 336884 454860 336890 454872
rect 361022 454860 361028 454872
rect 361080 454860 361086 454912
rect 219250 454792 219256 454844
rect 219308 454832 219314 454844
rect 244274 454832 244280 454844
rect 219308 454804 244280 454832
rect 219308 454792 219314 454804
rect 244274 454792 244280 454804
rect 244332 454792 244338 454844
rect 270586 454792 270592 454844
rect 270644 454832 270650 454844
rect 287238 454832 287244 454844
rect 270644 454804 287244 454832
rect 270644 454792 270650 454804
rect 287238 454792 287244 454804
rect 287296 454792 287302 454844
rect 302418 454792 302424 454844
rect 302476 454832 302482 454844
rect 580258 454832 580264 454844
rect 302476 454804 580264 454832
rect 302476 454792 302482 454804
rect 580258 454792 580264 454804
rect 580316 454792 580322 454844
rect 219342 454724 219348 454776
rect 219400 454764 219406 454776
rect 247126 454764 247132 454776
rect 219400 454736 247132 454764
rect 219400 454724 219406 454736
rect 247126 454724 247132 454736
rect 247184 454724 247190 454776
rect 267090 454724 267096 454776
rect 267148 454764 267154 454776
rect 283006 454764 283012 454776
rect 267148 454736 283012 454764
rect 267148 454724 267154 454736
rect 283006 454724 283012 454736
rect 283064 454724 283070 454776
rect 300210 454724 300216 454776
rect 300268 454764 300274 454776
rect 580350 454764 580356 454776
rect 300268 454736 580356 454764
rect 300268 454724 300274 454736
rect 580350 454724 580356 454736
rect 580408 454724 580414 454776
rect 217870 454656 217876 454708
rect 217928 454696 217934 454708
rect 255866 454696 255872 454708
rect 217928 454668 255872 454696
rect 217928 454656 217934 454668
rect 255866 454656 255872 454668
rect 255924 454656 255930 454708
rect 268562 454656 268568 454708
rect 268620 454696 268626 454708
rect 285858 454696 285864 454708
rect 268620 454668 285864 454696
rect 268620 454656 268626 454668
rect 285858 454656 285864 454668
rect 285916 454656 285922 454708
rect 298094 454656 298100 454708
rect 298152 454696 298158 454708
rect 580534 454696 580540 454708
rect 298152 454668 580540 454696
rect 298152 454656 298158 454668
rect 580534 454656 580540 454668
rect 580592 454656 580598 454708
rect 84838 453704 84844 453756
rect 84896 453744 84902 453756
rect 330202 453744 330208 453756
rect 84896 453716 330208 453744
rect 84896 453704 84902 453716
rect 330202 453704 330208 453716
rect 330260 453704 330266 453756
rect 320266 453636 320272 453688
rect 320324 453676 320330 453688
rect 358262 453676 358268 453688
rect 320324 453648 358268 453676
rect 320324 453636 320330 453648
rect 358262 453636 358268 453648
rect 358320 453636 358326 453688
rect 329926 453568 329932 453620
rect 329984 453608 329990 453620
rect 362218 453608 362224 453620
rect 329984 453580 362224 453608
rect 329984 453568 329990 453580
rect 362218 453568 362224 453580
rect 362276 453568 362282 453620
rect 32398 453500 32404 453552
rect 32456 453540 32462 453552
rect 327074 453540 327080 453552
rect 32456 453512 327080 453540
rect 32456 453500 32462 453512
rect 327074 453500 327080 453512
rect 327132 453500 327138 453552
rect 327166 453500 327172 453552
rect 327224 453540 327230 453552
rect 361114 453540 361120 453552
rect 327224 453512 361120 453540
rect 327224 453500 327230 453512
rect 361114 453500 361120 453512
rect 361172 453500 361178 453552
rect 10318 453432 10324 453484
rect 10376 453472 10382 453484
rect 351914 453472 351920 453484
rect 10376 453444 351920 453472
rect 10376 453432 10382 453444
rect 351914 453432 351920 453444
rect 351972 453432 351978 453484
rect 4890 453364 4896 453416
rect 4948 453404 4954 453416
rect 352006 453404 352012 453416
rect 4948 453376 352012 453404
rect 4948 453364 4954 453376
rect 352006 453364 352012 453376
rect 352064 453364 352070 453416
rect 5074 453296 5080 453348
rect 5132 453336 5138 453348
rect 353386 453336 353392 453348
rect 5132 453308 353392 453336
rect 5132 453296 5138 453308
rect 353386 453296 353392 453308
rect 353444 453296 353450 453348
rect 322934 452208 322940 452260
rect 322992 452248 322998 452260
rect 358170 452248 358176 452260
rect 322992 452220 358176 452248
rect 322992 452208 322998 452220
rect 358170 452208 358176 452220
rect 358228 452208 358234 452260
rect 307938 452140 307944 452192
rect 307996 452180 308002 452192
rect 360930 452180 360936 452192
rect 307996 452152 360936 452180
rect 307996 452140 308002 452152
rect 360930 452140 360936 452152
rect 360988 452140 360994 452192
rect 310514 452072 310520 452124
rect 310572 452112 310578 452124
rect 364334 452112 364340 452124
rect 310572 452084 364340 452112
rect 310572 452072 310578 452084
rect 364334 452072 364340 452084
rect 364392 452072 364398 452124
rect 71774 452004 71780 452056
rect 71832 452044 71838 452056
rect 347866 452044 347872 452056
rect 71832 452016 347872 452044
rect 71832 452004 71838 452016
rect 347866 452004 347872 452016
rect 347924 452004 347930 452056
rect 10410 451936 10416 451988
rect 10468 451976 10474 451988
rect 331214 451976 331220 451988
rect 10468 451948 331220 451976
rect 10468 451936 10474 451948
rect 331214 451936 331220 451948
rect 331272 451936 331278 451988
rect 6914 451868 6920 451920
rect 6972 451908 6978 451920
rect 350626 451908 350632 451920
rect 6972 451880 350632 451908
rect 6972 451868 6978 451880
rect 350626 451868 350632 451880
rect 350684 451868 350690 451920
rect 303614 450848 303620 450900
rect 303672 450888 303678 450900
rect 360838 450888 360844 450900
rect 303672 450860 360844 450888
rect 303672 450848 303678 450860
rect 360838 450848 360844 450860
rect 360896 450848 360902 450900
rect 301314 450780 301320 450832
rect 301372 450820 301378 450832
rect 359458 450820 359464 450832
rect 301372 450792 359464 450820
rect 301372 450780 301378 450792
rect 359458 450780 359464 450792
rect 359516 450780 359522 450832
rect 305914 450712 305920 450764
rect 305972 450752 305978 450764
rect 494054 450752 494060 450764
rect 305972 450724 494060 450752
rect 305972 450712 305978 450724
rect 494054 450712 494060 450724
rect 494112 450712 494118 450764
rect 8938 450644 8944 450696
rect 8996 450684 9002 450696
rect 329098 450684 329104 450696
rect 8996 450656 329104 450684
rect 8996 450644 9002 450656
rect 329098 450644 329104 450656
rect 329156 450644 329162 450696
rect 4798 450576 4804 450628
rect 4856 450616 4862 450628
rect 324498 450616 324504 450628
rect 4856 450588 324504 450616
rect 4856 450576 4862 450588
rect 324498 450576 324504 450588
rect 324556 450576 324562 450628
rect 4982 450508 4988 450560
rect 5040 450548 5046 450560
rect 326798 450548 326804 450560
rect 5040 450520 326804 450548
rect 5040 450508 5046 450520
rect 326798 450508 326804 450520
rect 326856 450508 326862 450560
rect 299014 449420 299020 449472
rect 299072 449460 299078 449472
rect 358078 449460 358084 449472
rect 299072 449432 358084 449460
rect 299072 449420 299078 449432
rect 358078 449420 358084 449432
rect 358136 449420 358142 449472
rect 296714 449352 296720 449404
rect 296772 449392 296778 449404
rect 371878 449392 371884 449404
rect 296772 449364 371884 449392
rect 296772 449352 296778 449364
rect 371878 449352 371884 449364
rect 371936 449352 371942 449404
rect 169754 449284 169760 449336
rect 169812 449324 169818 449336
rect 317506 449324 317512 449336
rect 169812 449296 317512 449324
rect 169812 449284 169818 449296
rect 317506 449284 317512 449296
rect 317564 449284 317570 449336
rect 106918 449216 106924 449268
rect 106976 449256 106982 449268
rect 319806 449256 319812 449268
rect 106976 449228 319812 449256
rect 106976 449216 106982 449228
rect 319806 449216 319812 449228
rect 319864 449216 319870 449268
rect 3418 449148 3424 449200
rect 3476 449188 3482 449200
rect 325786 449188 325792 449200
rect 3476 449160 325792 449188
rect 3476 449148 3482 449160
rect 325786 449148 325792 449160
rect 325844 449148 325850 449200
rect 332134 449148 332140 449200
rect 332192 449188 332198 449200
rect 527174 449188 527180 449200
rect 332192 449160 527180 449188
rect 332192 449148 332198 449160
rect 527174 449148 527180 449160
rect 527232 449148 527238 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 233142 448576 233148 448588
rect 3200 448548 233148 448576
rect 3200 448536 3206 448548
rect 233142 448536 233148 448548
rect 233200 448536 233206 448588
rect 309778 448196 309784 448248
rect 309836 448236 309842 448248
rect 412634 448236 412640 448248
rect 309836 448208 412640 448236
rect 309836 448196 309842 448208
rect 412634 448196 412640 448208
rect 412692 448196 412698 448248
rect 153194 448128 153200 448180
rect 153252 448168 153258 448180
rect 319070 448168 319076 448180
rect 153252 448140 319076 448168
rect 153252 448128 153258 448140
rect 319070 448128 319076 448140
rect 319128 448128 319134 448180
rect 307478 448060 307484 448112
rect 307536 448100 307542 448112
rect 477494 448100 477500 448112
rect 307536 448072 477500 448100
rect 307536 448060 307542 448072
rect 477494 448060 477500 448072
rect 477552 448060 477558 448112
rect 88334 447992 88340 448044
rect 88392 448032 88398 448044
rect 321370 448032 321376 448044
rect 88392 448004 321376 448032
rect 88392 447992 88398 448004
rect 321370 447992 321376 448004
rect 321428 447992 321434 448044
rect 305178 447924 305184 447976
rect 305236 447964 305242 447976
rect 542354 447964 542360 447976
rect 305236 447936 542360 447964
rect 305236 447924 305242 447936
rect 542354 447924 542360 447936
rect 542412 447924 542418 447976
rect 23474 447856 23480 447908
rect 23532 447896 23538 447908
rect 323670 447896 323676 447908
rect 23532 447868 323676 447896
rect 23532 447856 23538 447868
rect 323670 447856 323676 447868
rect 323728 447856 323734 447908
rect 3510 447788 3516 447840
rect 3568 447828 3574 447840
rect 332962 447828 332968 447840
rect 3568 447800 332968 447828
rect 3568 447788 3574 447800
rect 332962 447788 332968 447800
rect 333020 447788 333026 447840
rect 233142 446700 233148 446752
rect 233200 446740 233206 446752
rect 233200 446712 238754 446740
rect 233200 446700 233206 446712
rect 233234 446632 233240 446684
rect 233292 446672 233298 446684
rect 233878 446672 233884 446684
rect 233292 446644 233884 446672
rect 233292 446632 233298 446644
rect 233878 446632 233884 446644
rect 233936 446632 233942 446684
rect 234614 446632 234620 446684
rect 234672 446672 234678 446684
rect 235534 446672 235540 446684
rect 234672 446644 235540 446672
rect 234672 446632 234678 446644
rect 235534 446632 235540 446644
rect 235592 446632 235598 446684
rect 238726 446672 238754 446712
rect 248414 446700 248420 446752
rect 248472 446740 248478 446752
rect 249334 446740 249340 446752
rect 248472 446712 249340 446740
rect 248472 446700 248478 446712
rect 249334 446700 249340 446712
rect 249392 446700 249398 446752
rect 251174 446700 251180 446752
rect 251232 446740 251238 446752
rect 251726 446740 251732 446752
rect 251232 446712 251732 446740
rect 251232 446700 251238 446712
rect 251726 446700 251732 446712
rect 251784 446700 251790 446752
rect 252554 446700 252560 446752
rect 252612 446740 252618 446752
rect 253198 446740 253204 446752
rect 252612 446712 253204 446740
rect 252612 446700 252618 446712
rect 253198 446700 253204 446712
rect 253256 446700 253262 446752
rect 253934 446700 253940 446752
rect 253992 446740 253998 446752
rect 254670 446740 254676 446752
rect 253992 446712 254676 446740
rect 253992 446700 253998 446712
rect 254670 446700 254676 446712
rect 254728 446700 254734 446752
rect 258074 446700 258080 446752
rect 258132 446740 258138 446752
rect 258534 446740 258540 446752
rect 258132 446712 258540 446740
rect 258132 446700 258138 446712
rect 258534 446700 258540 446712
rect 258592 446700 258598 446752
rect 274634 446700 274640 446752
rect 274692 446740 274698 446752
rect 275646 446740 275652 446752
rect 274692 446712 275652 446740
rect 274692 446700 274698 446712
rect 275646 446700 275652 446712
rect 275704 446700 275710 446752
rect 278774 446700 278780 446752
rect 278832 446740 278838 446752
rect 279510 446740 279516 446752
rect 278832 446712 279516 446740
rect 278832 446700 278838 446712
rect 279510 446700 279516 446712
rect 279568 446700 279574 446752
rect 281534 446700 281540 446752
rect 281592 446740 281598 446752
rect 282454 446740 282460 446752
rect 281592 446712 282460 446740
rect 281592 446700 281598 446712
rect 282454 446700 282460 446712
rect 282512 446700 282518 446752
rect 289906 446700 289912 446752
rect 289964 446740 289970 446752
rect 290182 446740 290188 446752
rect 289964 446712 290188 446740
rect 289964 446700 289970 446712
rect 290182 446700 290188 446712
rect 290240 446700 290246 446752
rect 291194 446700 291200 446752
rect 291252 446740 291258 446752
rect 291838 446740 291844 446752
rect 291252 446712 291844 446740
rect 291252 446700 291258 446712
rect 291838 446700 291844 446712
rect 291896 446700 291902 446752
rect 292574 446700 292580 446752
rect 292632 446740 292638 446752
rect 293310 446740 293316 446752
rect 292632 446712 293316 446740
rect 292632 446700 292638 446712
rect 293310 446700 293316 446712
rect 293368 446700 293374 446752
rect 327074 446700 327080 446752
rect 327132 446740 327138 446752
rect 327902 446740 327908 446752
rect 327132 446712 327908 446740
rect 327132 446700 327138 446712
rect 327902 446700 327908 446712
rect 327960 446700 327966 446752
rect 351914 446700 351920 446752
rect 351972 446740 351978 446752
rect 352742 446740 352748 446752
rect 351972 446712 352748 446740
rect 351972 446700 351978 446712
rect 352742 446700 352748 446712
rect 352800 446700 352806 446752
rect 353294 446700 353300 446752
rect 353352 446740 353358 446752
rect 354214 446740 354220 446752
rect 353352 446712 354220 446740
rect 353352 446700 353358 446712
rect 354214 446700 354220 446712
rect 354272 446700 354278 446752
rect 355318 446672 355324 446684
rect 238726 446644 355324 446672
rect 355318 446632 355324 446644
rect 355376 446632 355382 446684
rect 238754 446564 238760 446616
rect 238812 446604 238818 446616
rect 239398 446604 239404 446616
rect 238812 446576 239404 446604
rect 238812 446564 238818 446576
rect 239398 446564 239404 446576
rect 239456 446564 239462 446616
rect 334434 446564 334440 446616
rect 334492 446604 334498 446616
rect 462314 446604 462320 446616
rect 334492 446576 462320 446604
rect 334492 446564 334498 446576
rect 462314 446564 462320 446576
rect 462372 446564 462378 446616
rect 201494 446496 201500 446548
rect 201552 446536 201558 446548
rect 343726 446536 343732 446548
rect 201552 446508 343732 446536
rect 201552 446496 201558 446508
rect 343726 446496 343732 446508
rect 343784 446496 343790 446548
rect 136634 446428 136640 446480
rect 136692 446468 136698 446480
rect 346026 446468 346032 446480
rect 136692 446440 346032 446468
rect 136692 446428 136698 446440
rect 346026 446428 346032 446440
rect 346084 446428 346090 446480
rect 40034 446360 40040 446412
rect 40092 446400 40098 446412
rect 322106 446400 322112 446412
rect 40092 446372 322112 446400
rect 40092 446360 40098 446372
rect 322106 446360 322112 446372
rect 322164 446360 322170 446412
rect 325234 446360 325240 446412
rect 325292 446400 325298 446412
rect 580442 446400 580448 446412
rect 325292 446372 580448 446400
rect 325292 446360 325298 446372
rect 580442 446360 580448 446372
rect 580500 446360 580506 446412
rect 255958 445680 255964 445732
rect 256016 445720 256022 445732
rect 256016 445692 258074 445720
rect 256016 445680 256022 445692
rect 258046 445652 258074 445692
rect 260098 445680 260104 445732
rect 260156 445720 260162 445732
rect 262030 445720 262036 445732
rect 260156 445692 262036 445720
rect 260156 445680 260162 445692
rect 262030 445680 262036 445692
rect 262088 445680 262094 445732
rect 262858 445680 262864 445732
rect 262916 445720 262922 445732
rect 266630 445720 266636 445732
rect 262916 445692 266636 445720
rect 262916 445680 262922 445692
rect 266630 445680 266636 445692
rect 266688 445680 266694 445732
rect 268194 445720 268200 445732
rect 267706 445692 268200 445720
rect 260466 445652 260472 445664
rect 258046 445624 260472 445652
rect 260466 445612 260472 445624
rect 260524 445612 260530 445664
rect 265618 445612 265624 445664
rect 265676 445652 265682 445664
rect 267706 445652 267734 445692
rect 268194 445680 268200 445692
rect 268252 445680 268258 445732
rect 265676 445624 267734 445652
rect 265676 445612 265682 445624
rect 313642 445476 313648 445528
rect 313700 445516 313706 445528
rect 340966 445516 340972 445528
rect 313700 445488 340972 445516
rect 313700 445476 313706 445488
rect 340966 445476 340972 445488
rect 341024 445476 341030 445528
rect 178770 445408 178776 445460
rect 178828 445448 178834 445460
rect 349154 445448 349160 445460
rect 178828 445420 349160 445448
rect 178828 445408 178834 445420
rect 349154 445408 349160 445420
rect 349212 445408 349218 445460
rect 7558 445340 7564 445392
rect 7616 445380 7622 445392
rect 351454 445380 351460 445392
rect 7616 445352 351460 445380
rect 7616 445340 7622 445352
rect 351454 445340 351460 445352
rect 351512 445340 351518 445392
rect 261478 445272 261484 445324
rect 261536 445312 261542 445324
rect 265066 445312 265072 445324
rect 261536 445284 265072 445312
rect 261536 445272 261542 445284
rect 265066 445272 265072 445284
rect 265124 445272 265130 445324
rect 341426 445272 341432 445324
rect 341484 445312 341490 445324
rect 358814 445312 358820 445324
rect 341484 445284 358820 445312
rect 341484 445272 341490 445284
rect 358814 445272 358820 445284
rect 358872 445272 358878 445324
rect 252462 445204 252468 445256
rect 252520 445244 252526 445256
rect 257430 445244 257436 445256
rect 252520 445216 257436 445244
rect 252520 445204 252526 445216
rect 257430 445204 257436 445216
rect 257488 445204 257494 445256
rect 339126 445204 339132 445256
rect 339184 445244 339190 445256
rect 358998 445244 359004 445256
rect 339184 445216 359004 445244
rect 339184 445204 339190 445216
rect 358998 445204 359004 445216
rect 359056 445204 359062 445256
rect 314470 445136 314476 445188
rect 314528 445176 314534 445188
rect 357434 445176 357440 445188
rect 314528 445148 357440 445176
rect 314528 445136 314534 445148
rect 357434 445136 357440 445148
rect 357492 445136 357498 445188
rect 257982 445068 257988 445120
rect 258040 445108 258046 445120
rect 263594 445108 263600 445120
rect 258040 445080 263600 445108
rect 258040 445068 258046 445080
rect 263594 445068 263600 445080
rect 263652 445068 263658 445120
rect 312906 445068 312912 445120
rect 312964 445108 312970 445120
rect 358906 445108 358912 445120
rect 312964 445080 358912 445108
rect 312964 445068 312970 445080
rect 358906 445068 358912 445080
rect 358964 445068 358970 445120
rect 217962 445000 217968 445052
rect 218020 445040 218026 445052
rect 315206 445040 315212 445052
rect 218020 445012 315212 445040
rect 218020 445000 218026 445012
rect 315206 445000 315212 445012
rect 315264 445000 315270 445052
rect 318794 445000 318800 445052
rect 318852 445040 318858 445052
rect 356790 445040 356796 445052
rect 318852 445012 356796 445040
rect 318852 445000 318858 445012
rect 356790 445000 356796 445012
rect 356848 445000 356854 445052
rect 244918 444932 244924 444984
rect 244976 444972 244982 444984
rect 246574 444972 246580 444984
rect 244976 444944 246580 444972
rect 244976 444932 244982 444944
rect 246574 444932 246580 444944
rect 246632 444932 246638 444984
rect 315850 444932 315856 444984
rect 315908 444972 315914 444984
rect 358354 444972 358360 444984
rect 315908 444944 358360 444972
rect 315908 444932 315914 444944
rect 358354 444932 358360 444944
rect 358412 444932 358418 444984
rect 304166 444864 304172 444916
rect 304224 444904 304230 444916
rect 359918 444904 359924 444916
rect 304224 444876 359924 444904
rect 304224 444864 304230 444876
rect 359918 444864 359924 444876
rect 359976 444864 359982 444916
rect 232406 444796 232412 444848
rect 232464 444836 232470 444848
rect 337562 444836 337568 444848
rect 232464 444808 337568 444836
rect 232464 444796 232470 444808
rect 337562 444796 337568 444808
rect 337620 444796 337626 444848
rect 231210 444728 231216 444780
rect 231268 444768 231274 444780
rect 339862 444768 339868 444780
rect 231268 444740 339868 444768
rect 231268 444728 231274 444740
rect 339862 444728 339868 444740
rect 339920 444728 339926 444780
rect 247034 444660 247040 444712
rect 247092 444700 247098 444712
rect 360654 444700 360660 444712
rect 247092 444672 360660 444700
rect 247092 444660 247098 444672
rect 360654 444660 360660 444672
rect 360712 444660 360718 444712
rect 232222 444592 232228 444644
rect 232280 444632 232286 444644
rect 346854 444632 346860 444644
rect 232280 444604 346860 444632
rect 232280 444592 232286 444604
rect 346854 444592 346860 444604
rect 346912 444592 346918 444644
rect 209038 444524 209044 444576
rect 209096 444564 209102 444576
rect 349890 444564 349896 444576
rect 209096 444536 349896 444564
rect 209096 444524 209102 444536
rect 349890 444524 349896 444536
rect 349948 444524 349954 444576
rect 309042 444456 309048 444508
rect 309100 444496 309106 444508
rect 321554 444496 321560 444508
rect 309100 444468 321560 444496
rect 309100 444456 309106 444468
rect 321554 444456 321560 444468
rect 321612 444456 321618 444508
rect 349798 444456 349804 444508
rect 349856 444496 349862 444508
rect 359182 444496 359188 444508
rect 349856 444468 359188 444496
rect 349856 444456 349862 444468
rect 359182 444456 359188 444468
rect 359240 444456 359246 444508
rect 340874 444388 340880 444440
rect 340932 444428 340938 444440
rect 357618 444428 357624 444440
rect 340932 444400 357624 444428
rect 340932 444388 340938 444400
rect 357618 444388 357624 444400
rect 357676 444388 357682 444440
rect 342254 443776 342260 443828
rect 342312 443816 342318 443828
rect 580994 443816 581000 443828
rect 342312 443788 581000 443816
rect 342312 443776 342318 443788
rect 580994 443776 581000 443788
rect 581052 443776 581058 443828
rect 340966 443708 340972 443760
rect 341024 443748 341030 443760
rect 580626 443748 580632 443760
rect 341024 443720 580632 443748
rect 341024 443708 341030 443720
rect 580626 443708 580632 443720
rect 580684 443708 580690 443760
rect 3418 443640 3424 443692
rect 3476 443680 3482 443692
rect 247034 443680 247040 443692
rect 3476 443652 247040 443680
rect 3476 443640 3482 443652
rect 247034 443640 247040 443652
rect 247092 443640 247098 443692
rect 321554 443640 321560 443692
rect 321612 443680 321618 443692
rect 580534 443680 580540 443692
rect 321612 443652 580540 443680
rect 321612 443640 321618 443652
rect 580534 443640 580540 443652
rect 580592 443640 580598 443692
rect 325970 443572 325976 443624
rect 326028 443612 326034 443624
rect 335998 443612 336004 443624
rect 326028 443584 336004 443612
rect 326028 443572 326034 443584
rect 335998 443572 336004 443584
rect 336056 443572 336062 443624
rect 231118 443504 231124 443556
rect 231176 443544 231182 443556
rect 342162 443544 342168 443556
rect 231176 443516 342168 443544
rect 231176 443504 231182 443516
rect 342162 443504 342168 443516
rect 342220 443504 342226 443556
rect 231302 443436 231308 443488
rect 231360 443476 231366 443488
rect 356054 443476 356060 443488
rect 231360 443448 356060 443476
rect 231360 443436 231366 443448
rect 356054 443436 356060 443448
rect 356112 443436 356118 443488
rect 174538 443368 174544 443420
rect 174596 443408 174602 443420
rect 342990 443408 342996 443420
rect 174596 443380 342996 443408
rect 174596 443368 174602 443380
rect 342990 443368 342996 443380
rect 343048 443368 343054 443420
rect 84838 443300 84844 443352
rect 84896 443340 84902 443352
rect 340690 443340 340696 443352
rect 84896 443312 340696 443340
rect 84896 443300 84902 443312
rect 340690 443300 340696 443312
rect 340748 443300 340754 443352
rect 302142 443232 302148 443284
rect 302200 443272 302206 443284
rect 580350 443272 580356 443284
rect 302200 443244 580356 443272
rect 302200 443232 302206 443244
rect 580350 443232 580356 443244
rect 580408 443232 580414 443284
rect 297450 443164 297456 443216
rect 297508 443204 297514 443216
rect 580258 443204 580264 443216
rect 297508 443176 580264 443204
rect 297508 443164 297514 443176
rect 580258 443164 580264 443176
rect 580316 443164 580322 443216
rect 32398 443096 32404 443148
rect 32456 443136 32462 443148
rect 338298 443136 338304 443148
rect 32456 443108 338304 443136
rect 32456 443096 32462 443108
rect 338298 443096 338304 443108
rect 338356 443096 338362 443148
rect 8938 443028 8944 443080
rect 8996 443068 9002 443080
rect 325970 443068 325976 443080
rect 8996 443040 325976 443068
rect 8996 443028 9002 443040
rect 325970 443028 325976 443040
rect 326028 443028 326034 443080
rect 4890 442960 4896 443012
rect 4948 443000 4954 443012
rect 344462 443000 344468 443012
rect 4948 442972 344468 443000
rect 4948 442960 4954 442972
rect 344462 442960 344468 442972
rect 344520 442960 344526 443012
rect 3510 442484 3516 442536
rect 3568 442524 3574 442536
rect 304166 442524 304172 442536
rect 3568 442496 304172 442524
rect 3568 442484 3574 442496
rect 304166 442484 304172 442496
rect 304224 442484 304230 442536
rect 315850 442524 315856 442536
rect 307036 442496 315856 442524
rect 3786 442416 3792 442468
rect 3844 442456 3850 442468
rect 307036 442456 307064 442496
rect 315850 442484 315856 442496
rect 315908 442484 315914 442536
rect 318794 442456 318800 442468
rect 3844 442428 307064 442456
rect 307128 442428 318800 442456
rect 3844 442416 3850 442428
rect 3970 442348 3976 442400
rect 4028 442388 4034 442400
rect 307128 442388 307156 442428
rect 318794 442416 318800 442428
rect 318852 442416 318858 442468
rect 4028 442360 307156 442388
rect 311866 442360 325694 442388
rect 4028 442348 4034 442360
rect 3878 442280 3884 442332
rect 3936 442320 3942 442332
rect 311526 442320 311532 442332
rect 3936 442292 311532 442320
rect 3936 442280 3942 442292
rect 311526 442280 311532 442292
rect 311584 442280 311590 442332
rect 311710 442280 311716 442332
rect 311768 442320 311774 442332
rect 311866 442320 311894 442360
rect 325666 442320 325694 442360
rect 340874 442320 340880 442332
rect 311768 442292 311894 442320
rect 312004 442292 321554 442320
rect 325666 442292 340880 442320
rect 311768 442280 311774 442292
rect 3602 442212 3608 442264
rect 3660 442252 3666 442264
rect 312004 442252 312032 442292
rect 3660 442224 302234 442252
rect 3660 442212 3666 442224
rect 302206 442184 302234 442224
rect 309106 442224 312032 442252
rect 309106 442184 309134 442224
rect 312078 442212 312084 442264
rect 312136 442212 312142 442264
rect 316034 442212 316040 442264
rect 316092 442252 316098 442264
rect 316092 442224 316724 442252
rect 316092 442212 316098 442224
rect 302206 442156 309134 442184
rect 304442 442076 304448 442128
rect 304500 442076 304506 442128
rect 304460 441640 304488 442076
rect 312096 441708 312124 442212
rect 316696 441776 316724 442224
rect 318518 442212 318524 442264
rect 318576 442212 318582 442264
rect 318536 441844 318564 442212
rect 321526 442184 321554 442292
rect 340874 442280 340880 442292
rect 340932 442280 340938 442332
rect 349798 442252 349804 442264
rect 325666 442224 349804 442252
rect 325666 442184 325694 442224
rect 349798 442212 349804 442224
rect 349856 442212 349862 442264
rect 321526 442156 325694 442184
rect 363690 441844 363696 441856
rect 318536 441816 363696 441844
rect 363690 441804 363696 441816
rect 363748 441804 363754 441856
rect 363598 441776 363604 441788
rect 316696 441748 363604 441776
rect 363598 441736 363604 441748
rect 363656 441736 363662 441788
rect 364978 441708 364984 441720
rect 312096 441680 364984 441708
rect 364978 441668 364984 441680
rect 365036 441668 365042 441720
rect 580442 441640 580448 441652
rect 304460 441612 580448 441640
rect 580442 441600 580448 441612
rect 580500 441600 580506 441652
rect 3694 439492 3700 439544
rect 3752 439532 3758 439544
rect 232222 439532 232228 439544
rect 3752 439504 232228 439532
rect 3752 439492 3758 439504
rect 232222 439492 232228 439504
rect 232280 439492 232286 439544
rect 363690 431876 363696 431928
rect 363748 431916 363754 431928
rect 580166 431916 580172 431928
rect 363748 431888 580172 431916
rect 363748 431876 363754 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 8938 423620 8944 423632
rect 3384 423592 8944 423620
rect 3384 423580 3390 423592
rect 8938 423580 8944 423592
rect 8996 423580 9002 423632
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 232222 411244 232228 411256
rect 3384 411216 232228 411244
rect 3384 411204 3390 411216
rect 232222 411204 232228 411216
rect 232280 411204 232286 411256
rect 2866 398760 2872 398812
rect 2924 398800 2930 398812
rect 231302 398800 231308 398812
rect 2924 398772 231308 398800
rect 2924 398760 2930 398772
rect 231302 398760 231308 398772
rect 231360 398760 231366 398812
rect 363598 379448 363604 379500
rect 363656 379488 363662 379500
rect 579614 379488 579620 379500
rect 363656 379460 579620 379488
rect 363656 379448 363662 379460
rect 579614 379448 579620 379460
rect 579672 379448 579678 379500
rect 2866 372512 2872 372564
rect 2924 372552 2930 372564
rect 32398 372552 32404 372564
rect 2924 372524 32404 372552
rect 2924 372512 2930 372524
rect 32398 372512 32404 372524
rect 32456 372512 32462 372564
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 231210 358748 231216 358760
rect 3384 358720 231216 358748
rect 3384 358708 3390 358720
rect 231210 358708 231216 358720
rect 231268 358708 231274 358760
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 84838 320124 84844 320136
rect 3384 320096 84844 320124
rect 3384 320084 3390 320096
rect 84838 320084 84844 320096
rect 84896 320084 84902 320136
rect 309410 310496 309416 310548
rect 309468 310536 309474 310548
rect 309778 310536 309784 310548
rect 309468 310508 309784 310536
rect 309468 310496 309474 310508
rect 309778 310496 309784 310508
rect 309836 310496 309842 310548
rect 310790 310496 310796 310548
rect 310848 310536 310854 310548
rect 311158 310536 311164 310548
rect 310848 310508 311164 310536
rect 310848 310496 310854 310508
rect 311158 310496 311164 310508
rect 311216 310496 311222 310548
rect 216122 309068 216128 309120
rect 216180 309108 216186 309120
rect 279970 309108 279976 309120
rect 216180 309080 279976 309108
rect 216180 309068 216186 309080
rect 279970 309068 279976 309080
rect 280028 309068 280034 309120
rect 354950 309068 354956 309120
rect 355008 309108 355014 309120
rect 369210 309108 369216 309120
rect 355008 309080 369216 309108
rect 355008 309068 355014 309080
rect 369210 309068 369216 309080
rect 369268 309068 369274 309120
rect 189718 309000 189724 309052
rect 189776 309040 189782 309052
rect 255774 309040 255780 309052
rect 189776 309012 255780 309040
rect 189776 309000 189782 309012
rect 255774 309000 255780 309012
rect 255832 309000 255838 309052
rect 353110 309000 353116 309052
rect 353168 309040 353174 309052
rect 366450 309040 366456 309052
rect 353168 309012 366456 309040
rect 353168 309000 353174 309012
rect 366450 309000 366456 309012
rect 366508 309000 366514 309052
rect 182818 308932 182824 308984
rect 182876 308972 182882 308984
rect 254394 308972 254400 308984
rect 182876 308944 254400 308972
rect 182876 308932 182882 308944
rect 254394 308932 254400 308944
rect 254452 308932 254458 308984
rect 318794 308932 318800 308984
rect 318852 308972 318858 308984
rect 319162 308972 319168 308984
rect 318852 308944 319168 308972
rect 318852 308932 318858 308944
rect 319162 308932 319168 308944
rect 319220 308932 319226 308984
rect 345382 308932 345388 308984
rect 345440 308972 345446 308984
rect 366542 308972 366548 308984
rect 345440 308944 366548 308972
rect 345440 308932 345446 308944
rect 366542 308932 366548 308944
rect 366600 308932 366606 308984
rect 213546 308864 213552 308916
rect 213604 308904 213610 308916
rect 286870 308904 286876 308916
rect 213604 308876 286876 308904
rect 213604 308864 213610 308876
rect 286870 308864 286876 308876
rect 286928 308864 286934 308916
rect 288894 308864 288900 308916
rect 288952 308904 288958 308916
rect 297266 308904 297272 308916
rect 288952 308876 297272 308904
rect 288952 308864 288958 308876
rect 297266 308864 297272 308876
rect 297324 308864 297330 308916
rect 311986 308864 311992 308916
rect 312044 308904 312050 308916
rect 312354 308904 312360 308916
rect 312044 308876 312360 308904
rect 312044 308864 312050 308876
rect 312354 308864 312360 308876
rect 312412 308864 312418 308916
rect 316126 308864 316132 308916
rect 316184 308904 316190 308916
rect 317046 308904 317052 308916
rect 316184 308876 317052 308904
rect 316184 308864 316190 308876
rect 317046 308864 317052 308876
rect 317104 308864 317110 308916
rect 317414 308864 317420 308916
rect 317472 308904 317478 308916
rect 317782 308904 317788 308916
rect 317472 308876 317788 308904
rect 317472 308864 317478 308876
rect 317782 308864 317788 308876
rect 317840 308864 317846 308916
rect 318978 308864 318984 308916
rect 319036 308904 319042 308916
rect 319530 308904 319536 308916
rect 319036 308876 319536 308904
rect 319036 308864 319042 308876
rect 319530 308864 319536 308876
rect 319588 308864 319594 308916
rect 320174 308864 320180 308916
rect 320232 308904 320238 308916
rect 320634 308904 320640 308916
rect 320232 308876 320640 308904
rect 320232 308864 320238 308876
rect 320634 308864 320640 308876
rect 320692 308864 320698 308916
rect 328454 308864 328460 308916
rect 328512 308904 328518 308916
rect 328822 308904 328828 308916
rect 328512 308876 328828 308904
rect 328512 308864 328518 308876
rect 328822 308864 328828 308876
rect 328880 308864 328886 308916
rect 346302 308864 346308 308916
rect 346360 308904 346366 308916
rect 368750 308904 368756 308916
rect 346360 308876 368756 308904
rect 346360 308864 346366 308876
rect 368750 308864 368756 308876
rect 368808 308864 368814 308916
rect 178678 308796 178684 308848
rect 178736 308836 178742 308848
rect 253014 308836 253020 308848
rect 178736 308808 253020 308836
rect 178736 308796 178742 308808
rect 253014 308796 253020 308808
rect 253072 308796 253078 308848
rect 293954 308796 293960 308848
rect 294012 308836 294018 308848
rect 354766 308836 354772 308848
rect 294012 308808 354772 308836
rect 294012 308796 294018 308808
rect 354766 308796 354772 308808
rect 354824 308796 354830 308848
rect 355410 308796 355416 308848
rect 355468 308836 355474 308848
rect 361298 308836 361304 308848
rect 355468 308808 361304 308836
rect 355468 308796 355474 308808
rect 361298 308796 361304 308808
rect 361356 308796 361362 308848
rect 68278 308728 68284 308780
rect 68336 308768 68342 308780
rect 240686 308768 240692 308780
rect 68336 308740 240692 308768
rect 68336 308728 68342 308740
rect 240686 308728 240692 308740
rect 240744 308728 240750 308780
rect 290734 308728 290740 308780
rect 290792 308768 290798 308780
rect 290792 308740 355456 308768
rect 290792 308728 290798 308740
rect 355428 308712 355456 308740
rect 43438 308660 43444 308712
rect 43496 308700 43502 308712
rect 236362 308700 236368 308712
rect 43496 308672 236368 308700
rect 43496 308660 43502 308672
rect 236362 308660 236368 308672
rect 236420 308660 236426 308712
rect 290918 308660 290924 308712
rect 290976 308700 290982 308712
rect 354674 308700 354680 308712
rect 290976 308672 354680 308700
rect 290976 308660 290982 308672
rect 354674 308660 354680 308672
rect 354732 308660 354738 308712
rect 355410 308660 355416 308712
rect 355468 308660 355474 308712
rect 357250 308660 357256 308712
rect 357308 308700 357314 308712
rect 357308 308672 364334 308700
rect 357308 308660 357314 308672
rect 46198 308592 46204 308644
rect 46256 308632 46262 308644
rect 239306 308632 239312 308644
rect 46256 308604 239312 308632
rect 46256 308592 46262 308604
rect 239306 308592 239312 308604
rect 239364 308592 239370 308644
rect 290274 308592 290280 308644
rect 290332 308632 290338 308644
rect 355686 308632 355692 308644
rect 290332 308604 355692 308632
rect 290332 308592 290338 308604
rect 355686 308592 355692 308604
rect 355744 308592 355750 308644
rect 364306 308632 364334 308672
rect 367462 308632 367468 308644
rect 364306 308604 367468 308632
rect 367462 308592 367468 308604
rect 367520 308592 367526 308644
rect 35158 308524 35164 308576
rect 35216 308564 35222 308576
rect 234522 308564 234528 308576
rect 35216 308536 234528 308564
rect 35216 308524 35222 308536
rect 234522 308524 234528 308536
rect 234580 308524 234586 308576
rect 263686 308524 263692 308576
rect 263744 308564 263750 308576
rect 264882 308564 264888 308576
rect 263744 308536 264888 308564
rect 263744 308524 263750 308536
rect 264882 308524 264888 308536
rect 264940 308524 264946 308576
rect 265066 308524 265072 308576
rect 265124 308564 265130 308576
rect 265526 308564 265532 308576
rect 265124 308536 265532 308564
rect 265124 308524 265130 308536
rect 265526 308524 265532 308536
rect 265584 308524 265590 308576
rect 267826 308524 267832 308576
rect 267884 308564 267890 308576
rect 268838 308564 268844 308576
rect 267884 308536 268844 308564
rect 267884 308524 267890 308536
rect 268838 308524 268844 308536
rect 268896 308524 268902 308576
rect 269114 308524 269120 308576
rect 269172 308564 269178 308576
rect 270218 308564 270224 308576
rect 269172 308536 270224 308564
rect 269172 308524 269178 308536
rect 270218 308524 270224 308536
rect 270276 308524 270282 308576
rect 270494 308524 270500 308576
rect 270552 308564 270558 308576
rect 271506 308564 271512 308576
rect 270552 308536 271512 308564
rect 270552 308524 270558 308536
rect 271506 308524 271512 308536
rect 271564 308524 271570 308576
rect 291378 308524 291384 308576
rect 291436 308564 291442 308576
rect 291436 308536 292574 308564
rect 291436 308524 291442 308536
rect 32398 308456 32404 308508
rect 32456 308496 32462 308508
rect 233142 308496 233148 308508
rect 32456 308468 233148 308496
rect 32456 308456 32462 308468
rect 233142 308456 233148 308468
rect 233200 308456 233206 308508
rect 233326 308456 233332 308508
rect 233384 308496 233390 308508
rect 234246 308496 234252 308508
rect 233384 308468 234252 308496
rect 233384 308456 233390 308468
rect 234246 308456 234252 308468
rect 234304 308456 234310 308508
rect 263594 308456 263600 308508
rect 263652 308496 263658 308508
rect 264054 308496 264060 308508
rect 263652 308468 264060 308496
rect 263652 308456 263658 308468
rect 264054 308456 264060 308468
rect 264112 308456 264118 308508
rect 265342 308456 265348 308508
rect 265400 308496 265406 308508
rect 265894 308496 265900 308508
rect 265400 308468 265900 308496
rect 265400 308456 265406 308468
rect 265894 308456 265900 308468
rect 265952 308456 265958 308508
rect 267734 308456 267740 308508
rect 267792 308496 267798 308508
rect 268194 308496 268200 308508
rect 267792 308468 268200 308496
rect 267792 308456 267798 308468
rect 268194 308456 268200 308468
rect 268252 308456 268258 308508
rect 269206 308456 269212 308508
rect 269264 308496 269270 308508
rect 269666 308496 269672 308508
rect 269264 308468 269672 308496
rect 269264 308456 269270 308468
rect 269666 308456 269672 308468
rect 269724 308456 269730 308508
rect 270678 308456 270684 308508
rect 270736 308496 270742 308508
rect 271598 308496 271604 308508
rect 270736 308468 271604 308496
rect 270736 308456 270742 308468
rect 271598 308456 271604 308468
rect 271656 308456 271662 308508
rect 271966 308456 271972 308508
rect 272024 308496 272030 308508
rect 272978 308496 272984 308508
rect 272024 308468 272984 308496
rect 272024 308456 272030 308468
rect 272978 308456 272984 308468
rect 273036 308456 273042 308508
rect 292546 308496 292574 308536
rect 297266 308524 297272 308576
rect 297324 308564 297330 308576
rect 355318 308564 355324 308576
rect 297324 308536 355324 308564
rect 297324 308524 297330 308536
rect 355318 308524 355324 308536
rect 355376 308524 355382 308576
rect 355778 308524 355784 308576
rect 355836 308564 355842 308576
rect 355962 308564 355968 308576
rect 355836 308536 355968 308564
rect 355836 308524 355842 308536
rect 355962 308524 355968 308536
rect 356020 308524 356026 308576
rect 356790 308524 356796 308576
rect 356848 308564 356854 308576
rect 367554 308564 367560 308576
rect 356848 308536 367560 308564
rect 356848 308524 356854 308536
rect 367554 308524 367560 308536
rect 367612 308524 367618 308576
rect 292546 308468 354536 308496
rect 25498 308388 25504 308440
rect 25556 308428 25562 308440
rect 231762 308428 231768 308440
rect 25556 308400 231768 308428
rect 25556 308388 25562 308400
rect 231762 308388 231768 308400
rect 231820 308388 231826 308440
rect 231946 308388 231952 308440
rect 232004 308428 232010 308440
rect 232866 308428 232872 308440
rect 232004 308400 232872 308428
rect 232004 308388 232010 308400
rect 232866 308388 232872 308400
rect 232924 308388 232930 308440
rect 233510 308388 233516 308440
rect 233568 308428 233574 308440
rect 233878 308428 233884 308440
rect 233568 308400 233884 308428
rect 233568 308388 233574 308400
rect 233878 308388 233884 308400
rect 233936 308388 233942 308440
rect 263870 308388 263876 308440
rect 263928 308428 263934 308440
rect 264422 308428 264428 308440
rect 263928 308400 264428 308428
rect 263928 308388 263934 308400
rect 264422 308388 264428 308400
rect 264480 308388 264486 308440
rect 265250 308388 265256 308440
rect 265308 308428 265314 308440
rect 265802 308428 265808 308440
rect 265308 308400 265808 308428
rect 265308 308388 265314 308400
rect 265802 308388 265808 308400
rect 265860 308388 265866 308440
rect 266538 308388 266544 308440
rect 266596 308428 266602 308440
rect 267182 308428 267188 308440
rect 266596 308400 267188 308428
rect 266596 308388 266602 308400
rect 267182 308388 267188 308400
rect 267240 308388 267246 308440
rect 268010 308388 268016 308440
rect 268068 308428 268074 308440
rect 268562 308428 268568 308440
rect 268068 308400 268568 308428
rect 268068 308388 268074 308400
rect 268562 308388 268568 308400
rect 268620 308388 268626 308440
rect 269298 308388 269304 308440
rect 269356 308428 269362 308440
rect 269758 308428 269764 308440
rect 269356 308400 269764 308428
rect 269356 308388 269362 308400
rect 269758 308388 269764 308400
rect 269816 308388 269822 308440
rect 270586 308388 270592 308440
rect 270644 308428 270650 308440
rect 271046 308428 271052 308440
rect 270644 308400 271052 308428
rect 270644 308388 270650 308400
rect 271046 308388 271052 308400
rect 271104 308388 271110 308440
rect 272150 308388 272156 308440
rect 272208 308428 272214 308440
rect 272518 308428 272524 308440
rect 272208 308400 272524 308428
rect 272208 308388 272214 308400
rect 272518 308388 272524 308400
rect 272576 308388 272582 308440
rect 354508 308428 354536 308468
rect 354674 308456 354680 308508
rect 354732 308496 354738 308508
rect 355594 308496 355600 308508
rect 354732 308468 355600 308496
rect 354732 308456 354738 308468
rect 355594 308456 355600 308468
rect 355652 308456 355658 308508
rect 355870 308456 355876 308508
rect 355928 308496 355934 308508
rect 358078 308496 358084 308508
rect 355928 308468 358084 308496
rect 355928 308456 355934 308468
rect 358078 308456 358084 308468
rect 358136 308456 358142 308508
rect 360304 308468 364334 308496
rect 358262 308428 358268 308440
rect 292546 308400 350534 308428
rect 354508 308400 358268 308428
rect 216214 308320 216220 308372
rect 216272 308360 216278 308372
rect 279326 308360 279332 308372
rect 216272 308332 279332 308360
rect 216272 308320 216278 308332
rect 279326 308320 279332 308332
rect 279384 308320 279390 308372
rect 289170 308320 289176 308372
rect 289228 308360 289234 308372
rect 292546 308360 292574 308400
rect 289228 308332 292574 308360
rect 289228 308320 289234 308332
rect 312078 308320 312084 308372
rect 312136 308360 312142 308372
rect 313090 308360 313096 308372
rect 312136 308332 313096 308360
rect 312136 308320 312142 308332
rect 313090 308320 313096 308332
rect 313148 308320 313154 308372
rect 314654 308320 314660 308372
rect 314712 308360 314718 308372
rect 315390 308360 315396 308372
rect 314712 308332 315396 308360
rect 314712 308320 314718 308332
rect 315390 308320 315396 308332
rect 315448 308320 315454 308372
rect 316126 308320 316132 308372
rect 316184 308360 316190 308372
rect 316770 308360 316776 308372
rect 316184 308332 316776 308360
rect 316184 308320 316190 308332
rect 316770 308320 316776 308332
rect 316828 308320 316834 308372
rect 321554 308320 321560 308372
rect 321612 308360 321618 308372
rect 322474 308360 322480 308372
rect 321612 308332 322480 308360
rect 321612 308320 321618 308332
rect 322474 308320 322480 308332
rect 322532 308320 322538 308372
rect 322934 308320 322940 308372
rect 322992 308360 322998 308372
rect 323854 308360 323860 308372
rect 322992 308332 323860 308360
rect 322992 308320 322998 308332
rect 323854 308320 323860 308332
rect 323912 308320 323918 308372
rect 324314 308320 324320 308372
rect 324372 308360 324378 308372
rect 324590 308360 324596 308372
rect 324372 308332 324596 308360
rect 324372 308320 324378 308332
rect 324590 308320 324596 308332
rect 324648 308320 324654 308372
rect 325786 308320 325792 308372
rect 325844 308360 325850 308372
rect 326798 308360 326804 308372
rect 325844 308332 326804 308360
rect 325844 308320 325850 308332
rect 326798 308320 326804 308332
rect 326856 308320 326862 308372
rect 327074 308320 327080 308372
rect 327132 308360 327138 308372
rect 327442 308360 327448 308372
rect 327132 308332 327448 308360
rect 327132 308320 327138 308332
rect 327442 308320 327448 308332
rect 327500 308320 327506 308372
rect 330110 308320 330116 308372
rect 330168 308360 330174 308372
rect 330478 308360 330484 308372
rect 330168 308332 330484 308360
rect 330168 308320 330174 308332
rect 330478 308320 330484 308332
rect 330536 308320 330542 308372
rect 216306 308252 216312 308304
rect 216364 308292 216370 308304
rect 278590 308292 278596 308304
rect 216364 308264 278596 308292
rect 216364 308252 216370 308264
rect 278590 308252 278596 308264
rect 278648 308252 278654 308304
rect 311986 308252 311992 308304
rect 312044 308292 312050 308304
rect 312722 308292 312728 308304
rect 312044 308264 312728 308292
rect 312044 308252 312050 308264
rect 312722 308252 312728 308264
rect 312780 308252 312786 308304
rect 316034 308252 316040 308304
rect 316092 308292 316098 308304
rect 316402 308292 316408 308304
rect 316092 308264 316408 308292
rect 316092 308252 316098 308264
rect 316402 308252 316408 308264
rect 316460 308252 316466 308304
rect 317506 308252 317512 308304
rect 317564 308292 317570 308304
rect 317874 308292 317880 308304
rect 317564 308264 317880 308292
rect 317564 308252 317570 308264
rect 317874 308252 317880 308264
rect 317932 308252 317938 308304
rect 318886 308252 318892 308304
rect 318944 308292 318950 308304
rect 319254 308292 319260 308304
rect 318944 308264 319260 308292
rect 318944 308252 318950 308264
rect 319254 308252 319260 308264
rect 319312 308252 319318 308304
rect 324406 308252 324412 308304
rect 324464 308292 324470 308304
rect 325326 308292 325332 308304
rect 324464 308264 325332 308292
rect 324464 308252 324470 308264
rect 325326 308252 325332 308264
rect 325384 308252 325390 308304
rect 325694 308252 325700 308304
rect 325752 308292 325758 308304
rect 326614 308292 326620 308304
rect 325752 308264 326620 308292
rect 325752 308252 325758 308264
rect 326614 308252 326620 308264
rect 326672 308252 326678 308304
rect 327258 308252 327264 308304
rect 327316 308292 327322 308304
rect 328178 308292 328184 308304
rect 327316 308264 328184 308292
rect 327316 308252 327322 308264
rect 328178 308252 328184 308264
rect 328236 308252 328242 308304
rect 328546 308252 328552 308304
rect 328604 308292 328610 308304
rect 329190 308292 329196 308304
rect 328604 308264 329196 308292
rect 328604 308252 328610 308264
rect 329190 308252 329196 308264
rect 329248 308252 329254 308304
rect 329834 308252 329840 308304
rect 329892 308292 329898 308304
rect 330294 308292 330300 308304
rect 329892 308264 330300 308292
rect 329892 308252 329898 308264
rect 330294 308252 330300 308264
rect 330352 308252 330358 308304
rect 264974 308184 264980 308236
rect 265032 308224 265038 308236
rect 266262 308224 266268 308236
rect 265032 308196 266268 308224
rect 265032 308184 265038 308196
rect 266262 308184 266268 308196
rect 266320 308184 266326 308236
rect 269482 308184 269488 308236
rect 269540 308224 269546 308236
rect 270126 308224 270132 308236
rect 269540 308196 270132 308224
rect 269540 308184 269546 308196
rect 270126 308184 270132 308196
rect 270184 308184 270190 308236
rect 270862 308184 270868 308236
rect 270920 308224 270926 308236
rect 271138 308224 271144 308236
rect 270920 308196 271144 308224
rect 270920 308184 270926 308196
rect 271138 308184 271144 308196
rect 271196 308184 271202 308236
rect 317690 308184 317696 308236
rect 317748 308224 317754 308236
rect 318242 308224 318248 308236
rect 317748 308196 318248 308224
rect 317748 308184 317754 308196
rect 318242 308184 318248 308196
rect 318300 308184 318306 308236
rect 324590 308184 324596 308236
rect 324648 308224 324654 308236
rect 325234 308224 325240 308236
rect 324648 308196 325240 308224
rect 324648 308184 324654 308196
rect 325234 308184 325240 308196
rect 325292 308184 325298 308236
rect 329926 308184 329932 308236
rect 329984 308224 329990 308236
rect 330938 308224 330944 308236
rect 329984 308196 330944 308224
rect 329984 308184 329990 308196
rect 330938 308184 330944 308196
rect 330996 308184 331002 308236
rect 350506 308224 350534 308400
rect 358262 308388 358268 308400
rect 358320 308388 358326 308440
rect 359642 308388 359648 308440
rect 359700 308428 359706 308440
rect 360194 308428 360200 308440
rect 359700 308400 360200 308428
rect 359700 308388 359706 308400
rect 360194 308388 360200 308400
rect 360252 308388 360258 308440
rect 356330 308320 356336 308372
rect 356388 308360 356394 308372
rect 360304 308360 360332 308468
rect 361022 308388 361028 308440
rect 361080 308428 361086 308440
rect 361574 308428 361580 308440
rect 361080 308400 361580 308428
rect 361080 308388 361086 308400
rect 361574 308388 361580 308400
rect 361632 308388 361638 308440
rect 364306 308428 364334 308468
rect 368842 308428 368848 308440
rect 364306 308400 368848 308428
rect 368842 308388 368848 308400
rect 368900 308388 368906 308440
rect 356388 308332 360332 308360
rect 356388 308320 356394 308332
rect 360378 308320 360384 308372
rect 360436 308360 360442 308372
rect 361114 308360 361120 308372
rect 360436 308332 361120 308360
rect 360436 308320 360442 308332
rect 361114 308320 361120 308332
rect 361172 308320 361178 308372
rect 361298 308320 361304 308372
rect 361356 308360 361362 308372
rect 368934 308360 368940 308372
rect 361356 308332 368940 308360
rect 361356 308320 361362 308332
rect 368934 308320 368940 308332
rect 368992 308320 368998 308372
rect 353570 308252 353576 308304
rect 353628 308292 353634 308304
rect 353628 308264 357296 308292
rect 353628 308252 353634 308264
rect 355778 308224 355784 308236
rect 350506 308196 355784 308224
rect 355778 308184 355784 308196
rect 355836 308184 355842 308236
rect 219066 308116 219072 308168
rect 219124 308156 219130 308168
rect 277946 308156 277952 308168
rect 219124 308128 277952 308156
rect 219124 308116 219130 308128
rect 277946 308116 277952 308128
rect 278004 308116 278010 308168
rect 313274 308116 313280 308168
rect 313332 308156 313338 308168
rect 313642 308156 313648 308168
rect 313332 308128 313648 308156
rect 313332 308116 313338 308128
rect 313642 308116 313648 308128
rect 313700 308116 313706 308168
rect 315022 308116 315028 308168
rect 315080 308156 315086 308168
rect 315850 308156 315856 308168
rect 315080 308128 315856 308156
rect 315080 308116 315086 308128
rect 315850 308116 315856 308128
rect 315908 308116 315914 308168
rect 317046 308116 317052 308168
rect 317104 308156 317110 308168
rect 318058 308156 318064 308168
rect 317104 308128 318064 308156
rect 317104 308116 317110 308128
rect 318058 308116 318064 308128
rect 318116 308116 318122 308168
rect 318886 308116 318892 308168
rect 318944 308156 318950 308168
rect 319806 308156 319812 308168
rect 318944 308128 319812 308156
rect 318944 308116 318950 308128
rect 319806 308116 319812 308128
rect 319864 308116 319870 308168
rect 320450 308116 320456 308168
rect 320508 308156 320514 308168
rect 321094 308156 321100 308168
rect 320508 308128 321100 308156
rect 320508 308116 320514 308128
rect 321094 308116 321100 308128
rect 321152 308116 321158 308168
rect 328730 308116 328736 308168
rect 328788 308156 328794 308168
rect 329558 308156 329564 308168
rect 328788 308128 329564 308156
rect 328788 308116 328794 308128
rect 329558 308116 329564 308128
rect 329616 308116 329622 308168
rect 354030 308116 354036 308168
rect 354088 308156 354094 308168
rect 357268 308156 357296 308264
rect 357526 308252 357532 308304
rect 357584 308292 357590 308304
rect 366266 308292 366272 308304
rect 357584 308264 366272 308292
rect 357584 308252 357590 308264
rect 366266 308252 366272 308264
rect 366324 308252 366330 308304
rect 358078 308184 358084 308236
rect 358136 308224 358142 308236
rect 367830 308224 367836 308236
rect 358136 308196 367836 308224
rect 358136 308184 358142 308196
rect 367830 308184 367836 308196
rect 367888 308184 367894 308236
rect 366174 308156 366180 308168
rect 354088 308128 357112 308156
rect 357268 308128 366180 308156
rect 354088 308116 354094 308128
rect 231762 308048 231768 308100
rect 231820 308088 231826 308100
rect 236086 308088 236092 308100
rect 231820 308060 236092 308088
rect 231820 308048 231826 308060
rect 236086 308048 236092 308060
rect 236144 308048 236150 308100
rect 313550 308048 313556 308100
rect 313608 308088 313614 308100
rect 314470 308088 314476 308100
rect 313608 308060 314476 308088
rect 313608 308048 313614 308060
rect 314470 308048 314476 308060
rect 314528 308048 314534 308100
rect 354766 308048 354772 308100
rect 354824 308088 354830 308100
rect 355502 308088 355508 308100
rect 354824 308060 355508 308088
rect 354824 308048 354830 308060
rect 355502 308048 355508 308060
rect 355560 308048 355566 308100
rect 357084 308088 357112 308128
rect 366174 308116 366180 308128
rect 366232 308116 366238 308168
rect 366358 308088 366364 308100
rect 357084 308060 366364 308088
rect 366358 308048 366364 308060
rect 366416 308048 366422 308100
rect 233142 307980 233148 308032
rect 233200 308020 233206 308032
rect 237926 308020 237932 308032
rect 233200 307992 237932 308020
rect 233200 307980 233206 307992
rect 237926 307980 237932 307992
rect 237984 307980 237990 308032
rect 314746 307980 314752 308032
rect 314804 308020 314810 308032
rect 315114 308020 315120 308032
rect 314804 307992 315120 308020
rect 314804 307980 314810 307992
rect 315114 307980 315120 307992
rect 315172 307980 315178 308032
rect 325878 307980 325884 308032
rect 325936 308020 325942 308032
rect 326246 308020 326252 308032
rect 325936 307992 326252 308020
rect 325936 307980 325942 307992
rect 326246 307980 326252 307992
rect 326304 307980 326310 308032
rect 354490 307980 354496 308032
rect 354548 308020 354554 308032
rect 365070 308020 365076 308032
rect 354548 307992 365076 308020
rect 354548 307980 354554 307992
rect 365070 307980 365076 307992
rect 365128 307980 365134 308032
rect 322290 307912 322296 307964
rect 322348 307952 322354 307964
rect 323578 307952 323584 307964
rect 322348 307924 323584 307952
rect 322348 307912 322354 307924
rect 323578 307912 323584 307924
rect 323636 307912 323642 307964
rect 327074 307912 327080 307964
rect 327132 307952 327138 307964
rect 327810 307952 327816 307964
rect 327132 307924 327816 307952
rect 327132 307912 327138 307924
rect 327810 307912 327816 307924
rect 327868 307912 327874 307964
rect 352650 307912 352656 307964
rect 352708 307952 352714 307964
rect 357526 307952 357532 307964
rect 352708 307924 357532 307952
rect 352708 307912 352714 307924
rect 357526 307912 357532 307924
rect 357584 307912 357590 307964
rect 360562 307912 360568 307964
rect 360620 307952 360626 307964
rect 361206 307952 361212 307964
rect 360620 307924 361212 307952
rect 360620 307912 360626 307924
rect 361206 307912 361212 307924
rect 361264 307912 361270 307964
rect 253198 307844 253204 307896
rect 253256 307884 253262 307896
rect 258074 307884 258080 307896
rect 253256 307856 258080 307884
rect 253256 307844 253262 307856
rect 258074 307844 258080 307856
rect 258132 307844 258138 307896
rect 360286 307844 360292 307896
rect 360344 307884 360350 307896
rect 360654 307884 360660 307896
rect 360344 307856 360660 307884
rect 360344 307844 360350 307856
rect 360654 307844 360660 307856
rect 360712 307844 360718 307896
rect 254762 307776 254768 307828
rect 254820 307816 254826 307828
rect 258718 307816 258724 307828
rect 254820 307788 258724 307816
rect 254820 307776 254826 307788
rect 258718 307776 258724 307788
rect 258776 307776 258782 307828
rect 260650 307776 260656 307828
rect 260708 307816 260714 307828
rect 263502 307816 263508 307828
rect 260708 307788 263508 307816
rect 260708 307776 260714 307788
rect 263502 307776 263508 307788
rect 263560 307776 263566 307828
rect 361666 307776 361672 307828
rect 361724 307816 361730 307828
rect 361942 307816 361948 307828
rect 361724 307788 361948 307816
rect 361724 307776 361730 307788
rect 361942 307776 361948 307788
rect 362000 307776 362006 307828
rect 314654 307708 314660 307760
rect 314712 307748 314718 307760
rect 315482 307748 315488 307760
rect 314712 307720 315488 307748
rect 314712 307708 314718 307720
rect 315482 307708 315488 307720
rect 315540 307708 315546 307760
rect 361850 307708 361856 307760
rect 361908 307748 361914 307760
rect 362494 307748 362500 307760
rect 361908 307720 362500 307748
rect 361908 307708 361914 307720
rect 362494 307708 362500 307720
rect 362552 307708 362558 307760
rect 317506 307504 317512 307556
rect 317564 307544 317570 307556
rect 318610 307544 318616 307556
rect 317564 307516 318616 307544
rect 317564 307504 317570 307516
rect 318610 307504 318616 307516
rect 318668 307504 318674 307556
rect 313274 307368 313280 307420
rect 313332 307408 313338 307420
rect 314102 307408 314108 307420
rect 313332 307380 314108 307408
rect 313332 307368 313338 307380
rect 314102 307368 314108 307380
rect 314160 307368 314166 307420
rect 312354 307232 312360 307284
rect 312412 307272 312418 307284
rect 377398 307272 377404 307284
rect 312412 307244 377404 307272
rect 312412 307232 312418 307244
rect 377398 307232 377404 307244
rect 377456 307232 377462 307284
rect 207014 307164 207020 307216
rect 207072 307204 207078 307216
rect 272426 307204 272432 307216
rect 207072 307176 272432 307204
rect 207072 307164 207078 307176
rect 272426 307164 272432 307176
rect 272484 307164 272490 307216
rect 314010 307164 314016 307216
rect 314068 307204 314074 307216
rect 422294 307204 422300 307216
rect 314068 307176 422300 307204
rect 314068 307164 314074 307176
rect 422294 307164 422300 307176
rect 422352 307164 422358 307216
rect 178034 307096 178040 307148
rect 178092 307136 178098 307148
rect 266998 307136 267004 307148
rect 178092 307108 267004 307136
rect 178092 307096 178098 307108
rect 266998 307096 267004 307108
rect 267056 307096 267062 307148
rect 326154 307096 326160 307148
rect 326212 307136 326218 307148
rect 484394 307136 484400 307148
rect 326212 307108 484400 307136
rect 326212 307096 326218 307108
rect 484394 307096 484400 307108
rect 484452 307096 484458 307148
rect 67634 307028 67640 307080
rect 67692 307068 67698 307080
rect 245470 307068 245476 307080
rect 67692 307040 245476 307068
rect 67692 307028 67698 307040
rect 245470 307028 245476 307040
rect 245528 307028 245534 307080
rect 330754 307028 330760 307080
rect 330812 307068 330818 307080
rect 507854 307068 507860 307080
rect 330812 307040 507860 307068
rect 330812 307028 330818 307040
rect 507854 307028 507860 307040
rect 507912 307028 507918 307080
rect 235166 306824 235172 306876
rect 235224 306824 235230 306876
rect 307754 306824 307760 306876
rect 307812 306864 307818 306876
rect 307938 306864 307944 306876
rect 307812 306836 307944 306864
rect 307812 306824 307818 306836
rect 307938 306824 307944 306836
rect 307996 306824 308002 306876
rect 235074 306620 235080 306672
rect 235132 306660 235138 306672
rect 235184 306660 235212 306824
rect 248598 306688 248604 306740
rect 248656 306688 248662 306740
rect 285950 306688 285956 306740
rect 286008 306688 286014 306740
rect 336918 306688 336924 306740
rect 336976 306688 336982 306740
rect 235132 306632 235212 306660
rect 235132 306620 235138 306632
rect 248616 306536 248644 306688
rect 249702 306620 249708 306672
rect 249760 306660 249766 306672
rect 250254 306660 250260 306672
rect 249760 306632 250260 306660
rect 249760 306620 249766 306632
rect 250254 306620 250260 306632
rect 250312 306620 250318 306672
rect 249886 306552 249892 306604
rect 249944 306592 249950 306604
rect 250346 306592 250352 306604
rect 249944 306564 250352 306592
rect 249944 306552 249950 306564
rect 250346 306552 250352 306564
rect 250404 306552 250410 306604
rect 285968 306536 285996 306688
rect 297174 306552 297180 306604
rect 297232 306552 297238 306604
rect 303798 306552 303804 306604
rect 303856 306592 303862 306604
rect 304166 306592 304172 306604
rect 303856 306564 304172 306592
rect 303856 306552 303862 306564
rect 304166 306552 304172 306564
rect 304224 306552 304230 306604
rect 306374 306552 306380 306604
rect 306432 306592 306438 306604
rect 306926 306592 306932 306604
rect 306432 306564 306932 306592
rect 306432 306552 306438 306564
rect 306926 306552 306932 306564
rect 306984 306552 306990 306604
rect 320358 306552 320364 306604
rect 320416 306592 320422 306604
rect 320726 306592 320732 306604
rect 320416 306564 320732 306592
rect 320416 306552 320422 306564
rect 320726 306552 320732 306564
rect 320784 306552 320790 306604
rect 248598 306484 248604 306536
rect 248656 306484 248662 306536
rect 285950 306484 285956 306536
rect 286008 306484 286014 306536
rect 287146 306484 287152 306536
rect 287204 306524 287210 306536
rect 287514 306524 287520 306536
rect 287204 306496 287520 306524
rect 287204 306484 287210 306496
rect 287514 306484 287520 306496
rect 287572 306484 287578 306536
rect 236086 306416 236092 306468
rect 236144 306456 236150 306468
rect 237098 306456 237104 306468
rect 236144 306428 237104 306456
rect 236144 306416 236150 306428
rect 237098 306416 237104 306428
rect 237156 306416 237162 306468
rect 243262 306416 243268 306468
rect 243320 306456 243326 306468
rect 243446 306456 243452 306468
rect 243320 306428 243452 306456
rect 243320 306416 243326 306428
rect 243446 306416 243452 306428
rect 243504 306416 243510 306468
rect 247218 306416 247224 306468
rect 247276 306456 247282 306468
rect 247954 306456 247960 306468
rect 247276 306428 247960 306456
rect 247276 306416 247282 306428
rect 247954 306416 247960 306428
rect 248012 306416 248018 306468
rect 259546 306416 259552 306468
rect 259604 306456 259610 306468
rect 260190 306456 260196 306468
rect 259604 306428 260196 306456
rect 259604 306416 259610 306428
rect 260190 306416 260196 306428
rect 260248 306416 260254 306468
rect 285674 306416 285680 306468
rect 285732 306456 285738 306468
rect 286226 306456 286232 306468
rect 285732 306428 286232 306456
rect 285732 306416 285738 306428
rect 286226 306416 286232 306428
rect 286284 306416 286290 306468
rect 236270 306348 236276 306400
rect 236328 306388 236334 306400
rect 237006 306388 237012 306400
rect 236328 306360 237012 306388
rect 236328 306348 236334 306360
rect 237006 306348 237012 306360
rect 237064 306348 237070 306400
rect 237742 306348 237748 306400
rect 237800 306388 237806 306400
rect 238478 306388 238484 306400
rect 237800 306360 238484 306388
rect 237800 306348 237806 306360
rect 238478 306348 238484 306360
rect 238536 306348 238542 306400
rect 239122 306348 239128 306400
rect 239180 306388 239186 306400
rect 239950 306388 239956 306400
rect 239180 306360 239956 306388
rect 239180 306348 239186 306360
rect 239950 306348 239956 306360
rect 240008 306348 240014 306400
rect 243078 306348 243084 306400
rect 243136 306388 243142 306400
rect 244090 306388 244096 306400
rect 243136 306360 244096 306388
rect 243136 306348 243142 306360
rect 244090 306348 244096 306360
rect 244148 306348 244154 306400
rect 247126 306348 247132 306400
rect 247184 306388 247190 306400
rect 247586 306388 247592 306400
rect 247184 306360 247592 306388
rect 247184 306348 247190 306360
rect 247586 306348 247592 306360
rect 247644 306348 247650 306400
rect 248506 306348 248512 306400
rect 248564 306388 248570 306400
rect 248690 306388 248696 306400
rect 248564 306360 248696 306388
rect 248564 306348 248570 306360
rect 248690 306348 248696 306360
rect 248748 306348 248754 306400
rect 251174 306348 251180 306400
rect 251232 306388 251238 306400
rect 252186 306388 252192 306400
rect 251232 306360 252192 306388
rect 251232 306348 251238 306360
rect 252186 306348 252192 306360
rect 252244 306348 252250 306400
rect 252738 306348 252744 306400
rect 252796 306388 252802 306400
rect 253474 306388 253480 306400
rect 252796 306360 253480 306388
rect 252796 306348 252802 306360
rect 253474 306348 253480 306360
rect 253532 306348 253538 306400
rect 254210 306348 254216 306400
rect 254268 306388 254274 306400
rect 254670 306388 254676 306400
rect 254268 306360 254676 306388
rect 254268 306348 254274 306360
rect 254670 306348 254676 306360
rect 254728 306348 254734 306400
rect 255682 306348 255688 306400
rect 255740 306388 255746 306400
rect 256418 306388 256424 306400
rect 255740 306360 256424 306388
rect 255740 306348 255746 306360
rect 256418 306348 256424 306360
rect 256476 306348 256482 306400
rect 262398 306348 262404 306400
rect 262456 306388 262462 306400
rect 263042 306388 263048 306400
rect 262456 306360 263048 306388
rect 262456 306348 262462 306360
rect 263042 306348 263048 306360
rect 263100 306348 263106 306400
rect 271690 306348 271696 306400
rect 271748 306388 271754 306400
rect 276750 306388 276756 306400
rect 271748 306360 276756 306388
rect 271748 306348 271754 306360
rect 276750 306348 276756 306360
rect 276808 306348 276814 306400
rect 284294 306348 284300 306400
rect 284352 306388 284358 306400
rect 285214 306388 285220 306400
rect 284352 306360 285220 306388
rect 284352 306348 284358 306360
rect 285214 306348 285220 306360
rect 285272 306348 285278 306400
rect 293954 306348 293960 306400
rect 294012 306388 294018 306400
rect 294690 306388 294696 306400
rect 294012 306360 294696 306388
rect 294012 306348 294018 306360
rect 294690 306348 294696 306360
rect 294748 306348 294754 306400
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 231118 306320 231124 306332
rect 3384 306292 231124 306320
rect 3384 306280 3390 306292
rect 231118 306280 231124 306292
rect 231176 306280 231182 306332
rect 234890 306280 234896 306332
rect 234948 306320 234954 306332
rect 235718 306320 235724 306332
rect 234948 306292 235724 306320
rect 234948 306280 234954 306292
rect 235718 306280 235724 306292
rect 235776 306280 235782 306332
rect 236178 306280 236184 306332
rect 236236 306320 236242 306332
rect 236638 306320 236644 306332
rect 236236 306292 236644 306320
rect 236236 306280 236242 306292
rect 236638 306280 236644 306292
rect 236696 306280 236702 306332
rect 237650 306280 237656 306332
rect 237708 306320 237714 306332
rect 238386 306320 238392 306332
rect 237708 306292 238392 306320
rect 237708 306280 237714 306292
rect 238386 306280 238392 306292
rect 238444 306280 238450 306332
rect 238938 306280 238944 306332
rect 238996 306320 239002 306332
rect 239398 306320 239404 306332
rect 238996 306292 239404 306320
rect 238996 306280 239002 306292
rect 239398 306280 239404 306292
rect 239456 306280 239462 306332
rect 240410 306280 240416 306332
rect 240468 306320 240474 306332
rect 240870 306320 240876 306332
rect 240468 306292 240876 306320
rect 240468 306280 240474 306292
rect 240870 306280 240876 306292
rect 240928 306280 240934 306332
rect 242986 306280 242992 306332
rect 243044 306320 243050 306332
rect 243630 306320 243636 306332
rect 243044 306292 243636 306320
rect 243044 306280 243050 306292
rect 243630 306280 243636 306292
rect 243688 306280 243694 306332
rect 244366 306280 244372 306332
rect 244424 306320 244430 306332
rect 244734 306320 244740 306332
rect 244424 306292 244740 306320
rect 244424 306280 244430 306292
rect 244734 306280 244740 306292
rect 244792 306280 244798 306332
rect 245654 306280 245660 306332
rect 245712 306320 245718 306332
rect 246390 306320 246396 306332
rect 245712 306292 246396 306320
rect 245712 306280 245718 306292
rect 246390 306280 246396 306292
rect 246448 306280 246454 306332
rect 247402 306280 247408 306332
rect 247460 306320 247466 306332
rect 248046 306320 248052 306332
rect 247460 306292 248052 306320
rect 247460 306280 247466 306292
rect 248046 306280 248052 306292
rect 248104 306280 248110 306332
rect 248414 306280 248420 306332
rect 248472 306320 248478 306332
rect 249426 306320 249432 306332
rect 248472 306292 249432 306320
rect 248472 306280 248478 306292
rect 249426 306280 249432 306292
rect 249484 306280 249490 306332
rect 251358 306280 251364 306332
rect 251416 306320 251422 306332
rect 251726 306320 251732 306332
rect 251416 306292 251732 306320
rect 251416 306280 251422 306292
rect 251726 306280 251732 306292
rect 251784 306280 251790 306332
rect 252922 306280 252928 306332
rect 252980 306320 252986 306332
rect 253566 306320 253572 306332
rect 252980 306292 253572 306320
rect 252980 306280 252986 306292
rect 253566 306280 253572 306292
rect 253624 306280 253630 306332
rect 254302 306280 254308 306332
rect 254360 306320 254366 306332
rect 255038 306320 255044 306332
rect 254360 306292 255044 306320
rect 254360 306280 254366 306292
rect 255038 306280 255044 306292
rect 255096 306280 255102 306332
rect 255590 306280 255596 306332
rect 255648 306320 255654 306332
rect 256050 306320 256056 306332
rect 255648 306292 256056 306320
rect 255648 306280 255654 306292
rect 256050 306280 256056 306292
rect 256108 306280 256114 306332
rect 258350 306280 258356 306332
rect 258408 306320 258414 306332
rect 259178 306320 259184 306332
rect 258408 306292 259184 306320
rect 258408 306280 258414 306292
rect 259178 306280 259184 306292
rect 259236 306280 259242 306332
rect 262490 306280 262496 306332
rect 262548 306320 262554 306332
rect 263134 306320 263140 306332
rect 262548 306292 263140 306320
rect 262548 306280 262554 306292
rect 263134 306280 263140 306292
rect 263192 306280 263198 306332
rect 281350 306320 281356 306332
rect 273226 306292 281356 306320
rect 218882 306212 218888 306264
rect 218940 306252 218946 306264
rect 273226 306252 273254 306292
rect 281350 306280 281356 306292
rect 281408 306280 281414 306332
rect 284386 306280 284392 306332
rect 284444 306320 284450 306332
rect 284754 306320 284760 306332
rect 284444 306292 284760 306320
rect 284444 306280 284450 306292
rect 284754 306280 284760 306292
rect 284812 306280 284818 306332
rect 287238 306280 287244 306332
rect 287296 306320 287302 306332
rect 287974 306320 287980 306332
rect 287296 306292 287980 306320
rect 287296 306280 287302 306292
rect 287974 306280 287980 306292
rect 288032 306280 288038 306332
rect 288434 306280 288440 306332
rect 288492 306320 288498 306332
rect 289354 306320 289360 306332
rect 288492 306292 289360 306320
rect 288492 306280 288498 306292
rect 289354 306280 289360 306292
rect 289412 306280 289418 306332
rect 289814 306280 289820 306332
rect 289872 306320 289878 306332
rect 290458 306320 290464 306332
rect 289872 306292 290464 306320
rect 289872 306280 289878 306292
rect 290458 306280 290464 306292
rect 290516 306280 290522 306332
rect 294138 306280 294144 306332
rect 294196 306320 294202 306332
rect 294598 306320 294604 306332
rect 294196 306292 294604 306320
rect 294196 306280 294202 306292
rect 294598 306280 294604 306292
rect 294656 306280 294662 306332
rect 218940 306224 273254 306252
rect 218940 306212 218946 306224
rect 285766 306212 285772 306264
rect 285824 306252 285830 306264
rect 286134 306252 286140 306264
rect 285824 306224 286140 306252
rect 285824 306212 285830 306224
rect 286134 306212 286140 306224
rect 286192 306212 286198 306264
rect 287330 306212 287336 306264
rect 287388 306252 287394 306264
rect 287606 306252 287612 306264
rect 287388 306224 287612 306252
rect 287388 306212 287394 306224
rect 287606 306212 287612 306224
rect 287664 306212 287670 306264
rect 291194 306212 291200 306264
rect 291252 306252 291258 306264
rect 292298 306252 292304 306264
rect 291252 306224 292304 306252
rect 291252 306212 291258 306224
rect 292298 306212 292304 306224
rect 292356 306212 292362 306264
rect 292758 306212 292764 306264
rect 292816 306252 292822 306264
rect 293218 306252 293224 306264
rect 292816 306224 293224 306252
rect 292816 306212 292822 306224
rect 293218 306212 293224 306224
rect 293276 306212 293282 306264
rect 295334 306212 295340 306264
rect 295392 306252 295398 306264
rect 295794 306252 295800 306264
rect 295392 306224 295800 306252
rect 295392 306212 295398 306224
rect 295794 306212 295800 306224
rect 295852 306212 295858 306264
rect 296714 306212 296720 306264
rect 296772 306252 296778 306264
rect 297192 306252 297220 306552
rect 336936 306468 336964 306688
rect 357710 306552 357716 306604
rect 357768 306592 357774 306604
rect 358078 306592 358084 306604
rect 357768 306564 358084 306592
rect 357768 306552 357774 306564
rect 358078 306552 358084 306564
rect 358136 306552 358142 306604
rect 358906 306484 358912 306536
rect 358964 306524 358970 306536
rect 359274 306524 359280 306536
rect 358964 306496 359280 306524
rect 358964 306484 358970 306496
rect 359274 306484 359280 306496
rect 359332 306484 359338 306536
rect 299474 306416 299480 306468
rect 299532 306456 299538 306468
rect 299842 306456 299848 306468
rect 299532 306428 299848 306456
rect 299532 306416 299538 306428
rect 299842 306416 299848 306428
rect 299900 306416 299906 306468
rect 336918 306416 336924 306468
rect 336976 306416 336982 306468
rect 359090 306416 359096 306468
rect 359148 306456 359154 306468
rect 359458 306456 359464 306468
rect 359148 306428 359464 306456
rect 359148 306416 359154 306428
rect 359458 306416 359464 306428
rect 359516 306416 359522 306468
rect 298186 306348 298192 306400
rect 298244 306388 298250 306400
rect 299382 306388 299388 306400
rect 298244 306360 299388 306388
rect 298244 306348 298250 306360
rect 299382 306348 299388 306360
rect 299440 306348 299446 306400
rect 306650 306348 306656 306400
rect 306708 306388 306714 306400
rect 307478 306388 307484 306400
rect 306708 306360 307484 306388
rect 306708 306348 306714 306360
rect 307478 306348 307484 306360
rect 307536 306348 307542 306400
rect 334158 306348 334164 306400
rect 334216 306388 334222 306400
rect 334894 306388 334900 306400
rect 334216 306360 334900 306388
rect 334216 306348 334222 306360
rect 334894 306348 334900 306360
rect 334952 306348 334958 306400
rect 335446 306348 335452 306400
rect 335504 306388 335510 306400
rect 335722 306388 335728 306400
rect 335504 306360 335728 306388
rect 335504 306348 335510 306360
rect 335722 306348 335728 306360
rect 335780 306348 335786 306400
rect 336826 306348 336832 306400
rect 336884 306388 336890 306400
rect 338022 306388 338028 306400
rect 336884 306360 338028 306388
rect 336884 306348 336890 306360
rect 338022 306348 338028 306360
rect 338080 306348 338086 306400
rect 342254 306348 342260 306400
rect 342312 306388 342318 306400
rect 342806 306388 342812 306400
rect 342312 306360 342812 306388
rect 342312 306348 342318 306360
rect 342806 306348 342812 306360
rect 342864 306348 342870 306400
rect 358722 306348 358728 306400
rect 358780 306388 358786 306400
rect 358780 306360 367094 306388
rect 358780 306348 358786 306360
rect 298094 306280 298100 306332
rect 298152 306320 298158 306332
rect 299014 306320 299020 306332
rect 298152 306292 299020 306320
rect 298152 306280 298158 306292
rect 299014 306280 299020 306292
rect 299072 306280 299078 306332
rect 299566 306280 299572 306332
rect 299624 306320 299630 306332
rect 300762 306320 300768 306332
rect 299624 306292 300768 306320
rect 299624 306280 299630 306292
rect 300762 306280 300768 306292
rect 300820 306280 300826 306332
rect 300946 306280 300952 306332
rect 301004 306320 301010 306332
rect 301314 306320 301320 306332
rect 301004 306292 301320 306320
rect 301004 306280 301010 306292
rect 301314 306280 301320 306292
rect 301372 306280 301378 306332
rect 303614 306280 303620 306332
rect 303672 306320 303678 306332
rect 304534 306320 304540 306332
rect 303672 306292 304540 306320
rect 303672 306280 303678 306292
rect 304534 306280 304540 306292
rect 304592 306280 304598 306332
rect 306466 306280 306472 306332
rect 306524 306320 306530 306332
rect 306742 306320 306748 306332
rect 306524 306292 306748 306320
rect 306524 306280 306530 306292
rect 306742 306280 306748 306292
rect 306800 306280 306806 306332
rect 309226 306280 309232 306332
rect 309284 306320 309290 306332
rect 310146 306320 310152 306332
rect 309284 306292 310152 306320
rect 309284 306280 309290 306292
rect 310146 306280 310152 306292
rect 310204 306280 310210 306332
rect 310606 306280 310612 306332
rect 310664 306320 310670 306332
rect 311526 306320 311532 306332
rect 310664 306292 311532 306320
rect 310664 306280 310670 306292
rect 311526 306280 311532 306292
rect 311584 306280 311590 306332
rect 331582 306280 331588 306332
rect 331640 306320 331646 306332
rect 332318 306320 332324 306332
rect 331640 306292 332324 306320
rect 331640 306280 331646 306292
rect 332318 306280 332324 306292
rect 332376 306280 332382 306332
rect 332778 306280 332784 306332
rect 332836 306320 332842 306332
rect 333238 306320 333244 306332
rect 332836 306292 333244 306320
rect 332836 306280 332842 306292
rect 333238 306280 333244 306292
rect 333296 306280 333302 306332
rect 334066 306280 334072 306332
rect 334124 306320 334130 306332
rect 334802 306320 334808 306332
rect 334124 306292 334808 306320
rect 334124 306280 334130 306292
rect 334802 306280 334808 306292
rect 334860 306280 334866 306332
rect 335354 306280 335360 306332
rect 335412 306320 335418 306332
rect 336274 306320 336280 306332
rect 335412 306292 336280 306320
rect 335412 306280 335418 306292
rect 336274 306280 336280 306292
rect 336332 306280 336338 306332
rect 337010 306280 337016 306332
rect 337068 306320 337074 306332
rect 337562 306320 337568 306332
rect 337068 306292 337568 306320
rect 337068 306280 337074 306292
rect 337562 306280 337568 306292
rect 337620 306280 337626 306332
rect 338206 306280 338212 306332
rect 338264 306320 338270 306332
rect 338942 306320 338948 306332
rect 338264 306292 338948 306320
rect 338264 306280 338270 306292
rect 338942 306280 338948 306292
rect 339000 306280 339006 306332
rect 339494 306280 339500 306332
rect 339552 306320 339558 306332
rect 340322 306320 340328 306332
rect 339552 306292 340328 306320
rect 339552 306280 339558 306292
rect 340322 306280 340328 306292
rect 340380 306280 340386 306332
rect 340966 306280 340972 306332
rect 341024 306320 341030 306332
rect 341518 306320 341524 306332
rect 341024 306292 341524 306320
rect 341024 306280 341030 306292
rect 341518 306280 341524 306292
rect 341576 306280 341582 306332
rect 342438 306280 342444 306332
rect 342496 306320 342502 306332
rect 342898 306320 342904 306332
rect 342496 306292 342904 306320
rect 342496 306280 342502 306292
rect 342898 306280 342904 306292
rect 342956 306280 342962 306332
rect 347774 306280 347780 306332
rect 347832 306320 347838 306332
rect 348602 306320 348608 306332
rect 347832 306292 348608 306320
rect 347832 306280 347838 306292
rect 348602 306280 348608 306292
rect 348660 306280 348666 306332
rect 354858 306280 354864 306332
rect 354916 306320 354922 306332
rect 367066 306320 367094 306360
rect 370130 306320 370136 306332
rect 354916 306292 358860 306320
rect 367066 306292 370136 306320
rect 354916 306280 354922 306292
rect 296772 306224 297220 306252
rect 296772 306212 296778 306224
rect 298278 306212 298284 306264
rect 298336 306252 298342 306264
rect 298554 306252 298560 306264
rect 298336 306224 298560 306252
rect 298336 306212 298342 306224
rect 298554 306212 298560 306224
rect 298612 306212 298618 306264
rect 301038 306212 301044 306264
rect 301096 306252 301102 306264
rect 301222 306252 301228 306264
rect 301096 306224 301228 306252
rect 301096 306212 301102 306224
rect 301222 306212 301228 306224
rect 301280 306212 301286 306264
rect 302510 306212 302516 306264
rect 302568 306252 302574 306264
rect 303154 306252 303160 306264
rect 302568 306224 303160 306252
rect 302568 306212 302574 306224
rect 303154 306212 303160 306224
rect 303212 306212 303218 306264
rect 304994 306212 305000 306264
rect 305052 306252 305058 306264
rect 305362 306252 305368 306264
rect 305052 306224 305368 306252
rect 305052 306212 305058 306224
rect 305362 306212 305368 306224
rect 305420 306212 305426 306264
rect 341150 306212 341156 306264
rect 341208 306252 341214 306264
rect 341886 306252 341892 306264
rect 341208 306224 341892 306252
rect 341208 306212 341214 306224
rect 341886 306212 341892 306224
rect 341944 306212 341950 306264
rect 353386 306212 353392 306264
rect 353444 306252 353450 306264
rect 358722 306252 358728 306264
rect 353444 306224 358728 306252
rect 353444 306212 353450 306224
rect 358722 306212 358728 306224
rect 358780 306212 358786 306264
rect 358832 306252 358860 306292
rect 370130 306280 370136 306292
rect 370188 306280 370194 306332
rect 371694 306252 371700 306264
rect 358832 306224 371700 306252
rect 371694 306212 371700 306224
rect 371752 306212 371758 306264
rect 214558 306144 214564 306196
rect 214616 306184 214622 306196
rect 271690 306184 271696 306196
rect 214616 306156 271696 306184
rect 214616 306144 214622 306156
rect 271690 306144 271696 306156
rect 271748 306144 271754 306196
rect 287422 306144 287428 306196
rect 287480 306184 287486 306196
rect 288066 306184 288072 306196
rect 287480 306156 288072 306184
rect 287480 306144 287486 306156
rect 288066 306144 288072 306156
rect 288124 306144 288130 306196
rect 292574 306144 292580 306196
rect 292632 306184 292638 306196
rect 293034 306184 293040 306196
rect 292632 306156 293040 306184
rect 292632 306144 292638 306156
rect 293034 306144 293040 306156
rect 293092 306144 293098 306196
rect 296898 306144 296904 306196
rect 296956 306184 296962 306196
rect 297818 306184 297824 306196
rect 296956 306156 297824 306184
rect 296956 306144 296962 306156
rect 297818 306144 297824 306156
rect 297876 306144 297882 306196
rect 302418 306144 302424 306196
rect 302476 306184 302482 306196
rect 303062 306184 303068 306196
rect 302476 306156 303068 306184
rect 302476 306144 302482 306156
rect 303062 306144 303068 306156
rect 303120 306144 303126 306196
rect 306466 306144 306472 306196
rect 306524 306184 306530 306196
rect 307386 306184 307392 306196
rect 306524 306156 307392 306184
rect 306524 306144 306530 306156
rect 307386 306144 307392 306156
rect 307444 306144 307450 306196
rect 331398 306144 331404 306196
rect 331456 306184 331462 306196
rect 331950 306184 331956 306196
rect 331456 306156 331956 306184
rect 331456 306144 331462 306156
rect 331950 306144 331956 306156
rect 332008 306144 332014 306196
rect 332594 306144 332600 306196
rect 332652 306184 332658 306196
rect 333698 306184 333704 306196
rect 332652 306156 333704 306184
rect 332652 306144 332658 306156
rect 333698 306144 333704 306156
rect 333756 306144 333762 306196
rect 338390 306144 338396 306196
rect 338448 306184 338454 306196
rect 339034 306184 339040 306196
rect 338448 306156 339040 306184
rect 338448 306144 338454 306156
rect 339034 306144 339040 306156
rect 339092 306144 339098 306196
rect 339770 306144 339776 306196
rect 339828 306184 339834 306196
rect 340414 306184 340420 306196
rect 339828 306156 340420 306184
rect 339828 306144 339834 306156
rect 340414 306144 340420 306156
rect 340472 306144 340478 306196
rect 341242 306144 341248 306196
rect 341300 306184 341306 306196
rect 341978 306184 341984 306196
rect 341300 306156 341984 306184
rect 341300 306144 341306 306156
rect 341978 306144 341984 306156
rect 342036 306144 342042 306196
rect 353846 306144 353852 306196
rect 353904 306184 353910 306196
rect 371510 306184 371516 306196
rect 353904 306156 358952 306184
rect 353904 306144 353910 306156
rect 216582 306076 216588 306128
rect 216640 306116 216646 306128
rect 278866 306116 278872 306128
rect 216640 306088 278872 306116
rect 216640 306076 216646 306088
rect 278866 306076 278872 306088
rect 278924 306076 278930 306128
rect 284478 306076 284484 306128
rect 284536 306116 284542 306128
rect 284846 306116 284852 306128
rect 284536 306088 284852 306116
rect 284536 306076 284542 306088
rect 284846 306076 284852 306088
rect 284904 306076 284910 306128
rect 292666 306076 292672 306128
rect 292724 306116 292730 306128
rect 293678 306116 293684 306128
rect 292724 306088 293684 306116
rect 292724 306076 292730 306088
rect 293678 306076 293684 306088
rect 293736 306076 293742 306128
rect 296806 306076 296812 306128
rect 296864 306116 296870 306128
rect 298002 306116 298008 306128
rect 296864 306088 298008 306116
rect 296864 306076 296870 306088
rect 298002 306076 298008 306088
rect 298060 306076 298066 306128
rect 299658 306076 299664 306128
rect 299716 306116 299722 306128
rect 299934 306116 299940 306128
rect 299716 306088 299940 306116
rect 299716 306076 299722 306088
rect 299934 306076 299940 306088
rect 299992 306076 299998 306128
rect 301038 306076 301044 306128
rect 301096 306116 301102 306128
rect 302142 306116 302148 306128
rect 301096 306088 302148 306116
rect 301096 306076 301102 306088
rect 302142 306076 302148 306088
rect 302200 306076 302206 306128
rect 303890 306076 303896 306128
rect 303948 306116 303954 306128
rect 304902 306116 304908 306128
rect 303948 306088 304908 306116
rect 303948 306076 303954 306088
rect 304902 306076 304908 306088
rect 304960 306076 304966 306128
rect 304994 306076 305000 306128
rect 305052 306116 305058 306128
rect 306098 306116 306104 306128
rect 305052 306088 306104 306116
rect 305052 306076 305058 306088
rect 306098 306076 306104 306088
rect 306156 306076 306162 306128
rect 331214 306076 331220 306128
rect 331272 306116 331278 306128
rect 331674 306116 331680 306128
rect 331272 306088 331680 306116
rect 331272 306076 331278 306088
rect 331674 306076 331680 306088
rect 331732 306076 331738 306128
rect 350350 306076 350356 306128
rect 350408 306116 350414 306128
rect 358630 306116 358636 306128
rect 350408 306088 358636 306116
rect 350408 306076 350414 306088
rect 358630 306076 358636 306088
rect 358688 306076 358694 306128
rect 358924 306116 358952 306156
rect 359752 306156 371516 306184
rect 359752 306116 359780 306156
rect 371510 306144 371516 306156
rect 371568 306144 371574 306196
rect 358924 306088 359780 306116
rect 360102 306076 360108 306128
rect 360160 306116 360166 306128
rect 367738 306116 367744 306128
rect 360160 306088 367744 306116
rect 360160 306076 360166 306088
rect 367738 306076 367744 306088
rect 367796 306076 367802 306128
rect 214834 306008 214840 306060
rect 214892 306048 214898 306060
rect 278130 306048 278136 306060
rect 214892 306020 278136 306048
rect 214892 306008 214898 306020
rect 278130 306008 278136 306020
rect 278188 306008 278194 306060
rect 352190 306008 352196 306060
rect 352248 306048 352254 306060
rect 352248 306020 357848 306048
rect 352248 306008 352254 306020
rect 215202 305940 215208 305992
rect 215260 305980 215266 305992
rect 279510 305980 279516 305992
rect 215260 305952 279516 305980
rect 215260 305940 215266 305952
rect 279510 305940 279516 305952
rect 279568 305940 279574 305992
rect 299658 305940 299664 305992
rect 299716 305980 299722 305992
rect 300394 305980 300400 305992
rect 299716 305952 300400 305980
rect 299716 305940 299722 305952
rect 300394 305940 300400 305952
rect 300452 305940 300458 305992
rect 331214 305940 331220 305992
rect 331272 305980 331278 305992
rect 331858 305980 331864 305992
rect 331272 305952 331864 305980
rect 331272 305940 331278 305952
rect 331858 305940 331864 305952
rect 331916 305940 331922 305992
rect 335722 305940 335728 305992
rect 335780 305980 335786 305992
rect 336642 305980 336648 305992
rect 335780 305952 336648 305980
rect 335780 305940 335786 305952
rect 336642 305940 336648 305952
rect 336700 305940 336706 305992
rect 357820 305980 357848 306020
rect 359918 306008 359924 306060
rect 359976 306048 359982 306060
rect 371326 306048 371332 306060
rect 359976 306020 371332 306048
rect 359976 306008 359982 306020
rect 371326 306008 371332 306020
rect 371384 306008 371390 306060
rect 371418 305980 371424 305992
rect 357820 305952 371424 305980
rect 371418 305940 371424 305952
rect 371476 305940 371482 305992
rect 215938 305872 215944 305924
rect 215996 305912 216002 305924
rect 280246 305912 280252 305924
rect 215996 305884 280252 305912
rect 215996 305872 216002 305884
rect 280246 305872 280252 305884
rect 280304 305872 280310 305924
rect 348970 305872 348976 305924
rect 349028 305912 349034 305924
rect 367646 305912 367652 305924
rect 349028 305884 367652 305912
rect 349028 305872 349034 305884
rect 367646 305872 367652 305884
rect 367704 305872 367710 305924
rect 212442 305804 212448 305856
rect 212500 305844 212506 305856
rect 282270 305844 282276 305856
rect 212500 305816 282276 305844
rect 212500 305804 212506 305816
rect 282270 305804 282276 305816
rect 282328 305804 282334 305856
rect 335538 305804 335544 305856
rect 335596 305844 335602 305856
rect 336182 305844 336188 305856
rect 335596 305816 336188 305844
rect 335596 305804 335602 305816
rect 336182 305804 336188 305816
rect 336240 305804 336246 305856
rect 349706 305804 349712 305856
rect 349764 305844 349770 305856
rect 369118 305844 369124 305856
rect 349764 305816 369124 305844
rect 349764 305804 349770 305816
rect 369118 305804 369124 305816
rect 369176 305804 369182 305856
rect 217870 305736 217876 305788
rect 217928 305776 217934 305788
rect 287146 305776 287152 305788
rect 217928 305748 287152 305776
rect 217928 305736 217934 305748
rect 287146 305736 287152 305748
rect 287204 305736 287210 305788
rect 294046 305736 294052 305788
rect 294104 305776 294110 305788
rect 295058 305776 295064 305788
rect 294104 305748 295064 305776
rect 294104 305736 294110 305748
rect 295058 305736 295064 305748
rect 295116 305736 295122 305788
rect 357710 305736 357716 305788
rect 357768 305776 357774 305788
rect 358354 305776 358360 305788
rect 357768 305748 358360 305776
rect 357768 305736 357774 305748
rect 358354 305736 358360 305748
rect 358412 305736 358418 305788
rect 358446 305736 358452 305788
rect 358504 305776 358510 305788
rect 370406 305776 370412 305788
rect 358504 305748 370412 305776
rect 358504 305736 358510 305748
rect 370406 305736 370412 305748
rect 370464 305736 370470 305788
rect 212350 305668 212356 305720
rect 212408 305708 212414 305720
rect 281626 305708 281632 305720
rect 212408 305680 281632 305708
rect 212408 305668 212414 305680
rect 281626 305668 281632 305680
rect 281684 305668 281690 305720
rect 352926 305668 352932 305720
rect 352984 305708 352990 305720
rect 359918 305708 359924 305720
rect 352984 305680 359924 305708
rect 352984 305668 352990 305680
rect 359918 305668 359924 305680
rect 359976 305668 359982 305720
rect 360010 305668 360016 305720
rect 360068 305708 360074 305720
rect 371602 305708 371608 305720
rect 360068 305680 371608 305708
rect 360068 305668 360074 305680
rect 371602 305668 371608 305680
rect 371660 305668 371666 305720
rect 217686 305600 217692 305652
rect 217744 305640 217750 305652
rect 344462 305640 344468 305652
rect 217744 305612 344468 305640
rect 217744 305600 217750 305612
rect 344462 305600 344468 305612
rect 344520 305600 344526 305652
rect 345566 305600 345572 305652
rect 345624 305640 345630 305652
rect 370222 305640 370228 305652
rect 345624 305612 370228 305640
rect 345624 305600 345630 305612
rect 370222 305600 370228 305612
rect 370280 305600 370286 305652
rect 214926 305532 214932 305584
rect 214984 305572 214990 305584
rect 276106 305572 276112 305584
rect 214984 305544 276112 305572
rect 214984 305532 214990 305544
rect 276106 305532 276112 305544
rect 276164 305532 276170 305584
rect 354306 305532 354312 305584
rect 354364 305572 354370 305584
rect 370038 305572 370044 305584
rect 354364 305544 370044 305572
rect 354364 305532 354370 305544
rect 370038 305532 370044 305544
rect 370096 305532 370102 305584
rect 215110 305464 215116 305516
rect 215168 305504 215174 305516
rect 276290 305504 276296 305516
rect 215168 305476 276296 305504
rect 215168 305464 215174 305476
rect 276290 305464 276296 305476
rect 276348 305464 276354 305516
rect 347222 305464 347228 305516
rect 347280 305504 347286 305516
rect 362402 305504 362408 305516
rect 347280 305476 362408 305504
rect 347280 305464 347286 305476
rect 362402 305464 362408 305476
rect 362460 305464 362466 305516
rect 215018 305396 215024 305448
rect 215076 305436 215082 305448
rect 275462 305436 275468 305448
rect 215076 305408 275468 305436
rect 215076 305396 215082 305408
rect 275462 305396 275468 305408
rect 275520 305396 275526 305448
rect 355226 305396 355232 305448
rect 355284 305436 355290 305448
rect 365162 305436 365168 305448
rect 355284 305408 365168 305436
rect 355284 305396 355290 305408
rect 365162 305396 365168 305408
rect 365220 305396 365226 305448
rect 234706 305328 234712 305380
rect 234764 305368 234770 305380
rect 235626 305368 235632 305380
rect 234764 305340 235632 305368
rect 234764 305328 234770 305340
rect 235626 305328 235632 305340
rect 235684 305328 235690 305380
rect 240226 305328 240232 305380
rect 240284 305368 240290 305380
rect 241330 305368 241336 305380
rect 240284 305340 241336 305368
rect 240284 305328 240290 305340
rect 241330 305328 241336 305340
rect 241388 305328 241394 305380
rect 241790 305328 241796 305380
rect 241848 305368 241854 305380
rect 242342 305368 242348 305380
rect 241848 305340 242348 305368
rect 241848 305328 241854 305340
rect 242342 305328 242348 305340
rect 242400 305328 242406 305380
rect 244550 305328 244556 305380
rect 244608 305368 244614 305380
rect 245102 305368 245108 305380
rect 244608 305340 245108 305368
rect 244608 305328 244614 305340
rect 245102 305328 245108 305340
rect 245160 305328 245166 305380
rect 245930 305328 245936 305380
rect 245988 305368 245994 305380
rect 246482 305368 246488 305380
rect 245988 305340 246488 305368
rect 245988 305328 245994 305340
rect 246482 305328 246488 305340
rect 246540 305328 246546 305380
rect 248690 305328 248696 305380
rect 248748 305368 248754 305380
rect 248966 305368 248972 305380
rect 248748 305340 248972 305368
rect 248748 305328 248754 305340
rect 248966 305328 248972 305340
rect 249024 305328 249030 305380
rect 249794 305328 249800 305380
rect 249852 305368 249858 305380
rect 250254 305368 250260 305380
rect 249852 305340 250260 305368
rect 249852 305328 249858 305340
rect 250254 305328 250260 305340
rect 250312 305328 250318 305380
rect 251450 305328 251456 305380
rect 251508 305368 251514 305380
rect 252094 305368 252100 305380
rect 251508 305340 252100 305368
rect 251508 305328 251514 305340
rect 252094 305328 252100 305340
rect 252152 305328 252158 305380
rect 256694 305328 256700 305380
rect 256752 305368 256758 305380
rect 257430 305368 257436 305380
rect 256752 305340 257436 305368
rect 256752 305328 256758 305340
rect 257430 305328 257436 305340
rect 257488 305328 257494 305380
rect 258258 305328 258264 305380
rect 258316 305368 258322 305380
rect 258810 305368 258816 305380
rect 258316 305340 258816 305368
rect 258316 305328 258322 305340
rect 258810 305328 258816 305340
rect 258868 305328 258874 305380
rect 259454 305328 259460 305380
rect 259512 305368 259518 305380
rect 260098 305368 260104 305380
rect 259512 305340 260104 305368
rect 259512 305328 259518 305340
rect 260098 305328 260104 305340
rect 260156 305328 260162 305380
rect 260834 305328 260840 305380
rect 260892 305368 260898 305380
rect 261018 305368 261024 305380
rect 260892 305340 261024 305368
rect 260892 305328 260898 305340
rect 261018 305328 261024 305340
rect 261076 305328 261082 305380
rect 261202 305328 261208 305380
rect 261260 305368 261266 305380
rect 262122 305368 262128 305380
rect 261260 305340 262128 305368
rect 261260 305328 261266 305340
rect 262122 305328 262128 305340
rect 262180 305328 262186 305380
rect 307938 305328 307944 305380
rect 307996 305368 308002 305380
rect 308858 305368 308864 305380
rect 307996 305340 308864 305368
rect 307996 305328 308002 305340
rect 308858 305328 308864 305340
rect 308916 305328 308922 305380
rect 342346 305328 342352 305380
rect 342404 305368 342410 305380
rect 343358 305368 343364 305380
rect 342404 305340 343364 305368
rect 342404 305328 342410 305340
rect 343358 305328 343364 305340
rect 343416 305328 343422 305380
rect 351730 305328 351736 305380
rect 351788 305368 351794 305380
rect 358446 305368 358452 305380
rect 351788 305340 358452 305368
rect 351788 305328 351794 305340
rect 358446 305328 358452 305340
rect 358504 305328 358510 305380
rect 359274 305328 359280 305380
rect 359332 305368 359338 305380
rect 359826 305368 359832 305380
rect 359332 305340 359832 305368
rect 359332 305328 359338 305340
rect 359826 305328 359832 305340
rect 359884 305328 359890 305380
rect 244366 305260 244372 305312
rect 244424 305300 244430 305312
rect 245010 305300 245016 305312
rect 244424 305272 245016 305300
rect 244424 305260 244430 305272
rect 245010 305260 245016 305272
rect 245068 305260 245074 305312
rect 351086 305260 351092 305312
rect 351144 305300 351150 305312
rect 360010 305300 360016 305312
rect 351144 305272 360016 305300
rect 351144 305260 351150 305272
rect 360010 305260 360016 305272
rect 360068 305260 360074 305312
rect 260834 305192 260840 305244
rect 260892 305232 260898 305244
rect 261662 305232 261668 305244
rect 260892 305204 261668 305232
rect 260892 305192 260898 305204
rect 261662 305192 261668 305204
rect 261720 305192 261726 305244
rect 357802 305192 357808 305244
rect 357860 305232 357866 305244
rect 358538 305232 358544 305244
rect 357860 305204 358544 305232
rect 357860 305192 357866 305204
rect 358538 305192 358544 305204
rect 358596 305192 358602 305244
rect 357434 305124 357440 305176
rect 357492 305164 357498 305176
rect 357986 305164 357992 305176
rect 357492 305136 357992 305164
rect 357492 305124 357498 305136
rect 357986 305124 357992 305136
rect 358044 305124 358050 305176
rect 241514 305056 241520 305108
rect 241572 305096 241578 305108
rect 242250 305096 242256 305108
rect 241572 305068 242256 305096
rect 241572 305056 241578 305068
rect 242250 305056 242256 305068
rect 242308 305056 242314 305108
rect 295518 304920 295524 304972
rect 295576 304960 295582 304972
rect 296438 304960 296444 304972
rect 295576 304932 296444 304960
rect 295576 304920 295582 304932
rect 296438 304920 296444 304932
rect 296496 304920 296502 304972
rect 300854 304920 300860 304972
rect 300912 304960 300918 304972
rect 301682 304960 301688 304972
rect 300912 304932 301688 304960
rect 300912 304920 300918 304932
rect 301682 304920 301688 304932
rect 301740 304920 301746 304972
rect 309962 304444 309968 304496
rect 310020 304484 310026 304496
rect 400214 304484 400220 304496
rect 310020 304456 400220 304484
rect 310020 304444 310026 304456
rect 400214 304444 400220 304456
rect 400272 304444 400278 304496
rect 311158 304376 311164 304428
rect 311216 304416 311222 304428
rect 404354 304416 404360 304428
rect 311216 304388 404360 304416
rect 311216 304376 311222 304388
rect 404354 304376 404360 304388
rect 404412 304376 404418 304428
rect 297082 304308 297088 304360
rect 297140 304348 297146 304360
rect 297358 304348 297364 304360
rect 297140 304320 297364 304348
rect 297140 304308 297146 304320
rect 297358 304308 297364 304320
rect 297416 304308 297422 304360
rect 315114 304308 315120 304360
rect 315172 304348 315178 304360
rect 425054 304348 425060 304360
rect 315172 304320 425060 304348
rect 315172 304308 315178 304320
rect 425054 304308 425060 304320
rect 425112 304308 425118 304360
rect 217502 304240 217508 304292
rect 217560 304280 217566 304292
rect 351546 304280 351552 304292
rect 217560 304252 351552 304280
rect 217560 304240 217566 304252
rect 351546 304240 351552 304252
rect 351604 304240 351610 304292
rect 332962 304172 332968 304224
rect 333020 304212 333026 304224
rect 333330 304212 333336 304224
rect 333020 304184 333336 304212
rect 333020 304172 333026 304184
rect 333330 304172 333336 304184
rect 333388 304172 333394 304224
rect 261110 303968 261116 304020
rect 261168 304008 261174 304020
rect 261478 304008 261484 304020
rect 261168 303980 261484 304008
rect 261168 303968 261174 303980
rect 261478 303968 261484 303980
rect 261536 303968 261542 304020
rect 256786 303696 256792 303748
rect 256844 303736 256850 303748
rect 257154 303736 257160 303748
rect 256844 303708 257160 303736
rect 256844 303696 256850 303708
rect 257154 303696 257160 303708
rect 257212 303696 257218 303748
rect 273438 303696 273444 303748
rect 273496 303736 273502 303748
rect 274358 303736 274364 303748
rect 273496 303708 274364 303736
rect 273496 303696 273502 303708
rect 274358 303696 274364 303708
rect 274416 303696 274422 303748
rect 343634 303696 343640 303748
rect 343692 303736 343698 303748
rect 344646 303736 344652 303748
rect 343692 303708 344652 303736
rect 343692 303696 343698 303708
rect 344646 303696 344652 303708
rect 344704 303696 344710 303748
rect 213822 303560 213828 303612
rect 213880 303600 213886 303612
rect 279786 303600 279792 303612
rect 213880 303572 279792 303600
rect 213880 303560 213886 303572
rect 279786 303560 279792 303572
rect 279844 303560 279850 303612
rect 291286 303560 291292 303612
rect 291344 303600 291350 303612
rect 291470 303600 291476 303612
rect 291344 303572 291476 303600
rect 291344 303560 291350 303572
rect 291470 303560 291476 303572
rect 291528 303560 291534 303612
rect 352466 303560 352472 303612
rect 352524 303600 352530 303612
rect 371786 303600 371792 303612
rect 352524 303572 371792 303600
rect 352524 303560 352530 303572
rect 371786 303560 371792 303572
rect 371844 303560 371850 303612
rect 214466 303492 214472 303544
rect 214524 303532 214530 303544
rect 282086 303532 282092 303544
rect 214524 303504 282092 303532
rect 214524 303492 214530 303504
rect 282086 303492 282092 303504
rect 282144 303492 282150 303544
rect 348510 303492 348516 303544
rect 348568 303532 348574 303544
rect 367922 303532 367928 303544
rect 348568 303504 367928 303532
rect 348568 303492 348574 303504
rect 367922 303492 367928 303504
rect 367980 303492 367986 303544
rect 216030 303424 216036 303476
rect 216088 303464 216094 303476
rect 283374 303464 283380 303476
rect 216088 303436 283380 303464
rect 216088 303424 216094 303436
rect 283374 303424 283380 303436
rect 283432 303424 283438 303476
rect 291470 303424 291476 303476
rect 291528 303464 291534 303476
rect 291930 303464 291936 303476
rect 291528 303436 291936 303464
rect 291528 303424 291534 303436
rect 291930 303424 291936 303436
rect 291988 303424 291994 303476
rect 352006 303424 352012 303476
rect 352064 303464 352070 303476
rect 373074 303464 373080 303476
rect 352064 303436 373080 303464
rect 352064 303424 352070 303436
rect 373074 303424 373080 303436
rect 373132 303424 373138 303476
rect 213730 303356 213736 303408
rect 213788 303396 213794 303408
rect 282730 303396 282736 303408
rect 213788 303368 282736 303396
rect 213788 303356 213794 303368
rect 282730 303356 282736 303368
rect 282788 303356 282794 303408
rect 351270 303356 351276 303408
rect 351328 303396 351334 303408
rect 372706 303396 372712 303408
rect 351328 303368 372712 303396
rect 351328 303356 351334 303368
rect 372706 303356 372712 303368
rect 372764 303356 372770 303408
rect 213178 303288 213184 303340
rect 213236 303328 213242 303340
rect 282546 303328 282552 303340
rect 213236 303300 282552 303328
rect 213236 303288 213242 303300
rect 282546 303288 282552 303300
rect 282604 303288 282610 303340
rect 337102 303288 337108 303340
rect 337160 303328 337166 303340
rect 337654 303328 337660 303340
rect 337160 303300 337660 303328
rect 337160 303288 337166 303300
rect 337654 303288 337660 303300
rect 337712 303288 337718 303340
rect 347682 303288 347688 303340
rect 347740 303328 347746 303340
rect 369302 303328 369308 303340
rect 347740 303300 369308 303328
rect 347740 303288 347746 303300
rect 369302 303288 369308 303300
rect 369360 303288 369366 303340
rect 213362 303220 213368 303272
rect 213420 303260 213426 303272
rect 283006 303260 283012 303272
rect 213420 303232 283012 303260
rect 213420 303220 213426 303232
rect 283006 303220 283012 303232
rect 283064 303220 283070 303272
rect 349890 303220 349896 303272
rect 349948 303260 349954 303272
rect 372798 303260 372804 303272
rect 349948 303232 372804 303260
rect 349948 303220 349954 303232
rect 372798 303220 372804 303232
rect 372856 303220 372862 303272
rect 211706 303152 211712 303204
rect 211764 303192 211770 303204
rect 281810 303192 281816 303204
rect 211764 303164 281816 303192
rect 211764 303152 211770 303164
rect 281810 303152 281816 303164
rect 281868 303152 281874 303204
rect 295610 303152 295616 303204
rect 295668 303192 295674 303204
rect 295978 303192 295984 303204
rect 295668 303164 295984 303192
rect 295668 303152 295674 303164
rect 295978 303152 295984 303164
rect 296036 303152 296042 303204
rect 305178 303152 305184 303204
rect 305236 303192 305242 303204
rect 306006 303192 306012 303204
rect 305236 303164 306012 303192
rect 305236 303152 305242 303164
rect 306006 303152 306012 303164
rect 306064 303152 306070 303204
rect 349246 303152 349252 303204
rect 349304 303192 349310 303204
rect 373166 303192 373172 303204
rect 349304 303164 373172 303192
rect 349304 303152 349310 303164
rect 373166 303152 373172 303164
rect 373224 303152 373230 303204
rect 214650 303084 214656 303136
rect 214708 303124 214714 303136
rect 287054 303124 287060 303136
rect 214708 303096 287060 303124
rect 214708 303084 214714 303096
rect 287054 303084 287060 303096
rect 287112 303084 287118 303136
rect 346486 303084 346492 303136
rect 346544 303124 346550 303136
rect 370498 303124 370504 303136
rect 346544 303096 370504 303124
rect 346544 303084 346550 303096
rect 370498 303084 370504 303096
rect 370556 303084 370562 303136
rect 211982 303016 211988 303068
rect 212040 303056 212046 303068
rect 345842 303056 345848 303068
rect 212040 303028 345848 303056
rect 212040 303016 212046 303028
rect 345842 303016 345848 303028
rect 345900 303016 345906 303068
rect 347406 303016 347412 303068
rect 347464 303056 347470 303068
rect 370682 303056 370688 303068
rect 347464 303028 370688 303056
rect 347464 303016 347470 303028
rect 370682 303016 370688 303028
rect 370740 303016 370746 303068
rect 256970 302948 256976 303000
rect 257028 302988 257034 303000
rect 257338 302988 257344 303000
rect 257028 302960 257344 302988
rect 257028 302948 257034 302960
rect 257338 302948 257344 302960
rect 257396 302948 257402 303000
rect 350626 302948 350632 303000
rect 350684 302988 350690 303000
rect 372890 302988 372896 303000
rect 350684 302960 372896 302988
rect 350684 302948 350690 302960
rect 372890 302948 372896 302960
rect 372948 302948 372954 303000
rect 213086 302880 213092 302932
rect 213144 302920 213150 302932
rect 346762 302920 346768 302932
rect 213144 302892 346768 302920
rect 213144 302880 213150 302892
rect 346762 302880 346768 302892
rect 346820 302880 346826 302932
rect 348326 302880 348332 302932
rect 348384 302920 348390 302932
rect 372982 302920 372988 302932
rect 348384 302892 372988 302920
rect 348384 302880 348390 302892
rect 372982 302880 372988 302892
rect 373040 302880 373046 302932
rect 217962 302812 217968 302864
rect 218020 302852 218026 302864
rect 283650 302852 283656 302864
rect 218020 302824 283656 302852
rect 218020 302812 218026 302824
rect 283650 302812 283656 302824
rect 283708 302812 283714 302864
rect 356054 302812 356060 302864
rect 356112 302852 356118 302864
rect 371878 302852 371884 302864
rect 356112 302824 371884 302852
rect 356112 302812 356118 302824
rect 371878 302812 371884 302824
rect 371936 302812 371942 302864
rect 215846 302744 215852 302796
rect 215904 302784 215910 302796
rect 280430 302784 280436 302796
rect 215904 302756 280436 302784
rect 215904 302744 215910 302756
rect 280430 302744 280436 302756
rect 280488 302744 280494 302796
rect 307846 302744 307852 302796
rect 307904 302784 307910 302796
rect 308766 302784 308772 302796
rect 307904 302756 308772 302784
rect 307904 302744 307910 302756
rect 308766 302744 308772 302756
rect 308824 302744 308830 302796
rect 355962 302744 355968 302796
rect 356020 302784 356026 302796
rect 370314 302784 370320 302796
rect 356020 302756 370320 302784
rect 356020 302744 356026 302756
rect 370314 302744 370320 302756
rect 370372 302744 370378 302796
rect 218974 302676 218980 302728
rect 219032 302716 219038 302728
rect 281166 302716 281172 302728
rect 219032 302688 281172 302716
rect 219032 302676 219038 302688
rect 281166 302676 281172 302688
rect 281224 302676 281230 302728
rect 356974 302676 356980 302728
rect 357032 302716 357038 302728
rect 370590 302716 370596 302728
rect 357032 302688 370596 302716
rect 357032 302676 357038 302688
rect 370590 302676 370596 302688
rect 370648 302676 370654 302728
rect 217410 302608 217416 302660
rect 217468 302648 217474 302660
rect 350810 302648 350816 302660
rect 217468 302620 350816 302648
rect 217468 302608 217474 302620
rect 350810 302608 350816 302620
rect 350868 302608 350874 302660
rect 358998 302608 359004 302660
rect 359056 302648 359062 302660
rect 359734 302648 359740 302660
rect 359056 302620 359740 302648
rect 359056 302608 359062 302620
rect 359734 302608 359740 302620
rect 359792 302608 359798 302660
rect 234982 302200 234988 302252
rect 235040 302240 235046 302252
rect 235258 302240 235264 302252
rect 235040 302212 235264 302240
rect 235040 302200 235046 302212
rect 235258 302200 235264 302212
rect 235316 302200 235322 302252
rect 306742 301656 306748 301708
rect 306800 301696 306806 301708
rect 382274 301696 382280 301708
rect 306800 301668 382280 301696
rect 306800 301656 306806 301668
rect 382274 301656 382280 301668
rect 382332 301656 382338 301708
rect 317874 301588 317880 301640
rect 317932 301628 317938 301640
rect 440234 301628 440240 301640
rect 317932 301600 440240 301628
rect 317932 301588 317938 301600
rect 440234 301588 440240 301600
rect 440292 301588 440298 301640
rect 340782 301520 340788 301572
rect 340840 301560 340846 301572
rect 560294 301560 560300 301572
rect 340840 301532 560300 301560
rect 340840 301520 340846 301532
rect 560294 301520 560300 301532
rect 560352 301520 560358 301572
rect 341426 301452 341432 301504
rect 341484 301492 341490 301504
rect 564434 301492 564440 301504
rect 341484 301464 564440 301492
rect 341484 301452 341490 301464
rect 564434 301452 564440 301464
rect 564492 301452 564498 301504
rect 213270 300772 213276 300824
rect 213328 300812 213334 300824
rect 283926 300812 283932 300824
rect 213328 300784 283932 300812
rect 213328 300772 213334 300784
rect 283926 300772 283932 300784
rect 283984 300772 283990 300824
rect 215754 300704 215760 300756
rect 215812 300744 215818 300756
rect 285858 300744 285864 300756
rect 215812 300716 285864 300744
rect 215812 300704 215818 300716
rect 285858 300704 285864 300716
rect 285916 300704 285922 300756
rect 216398 300636 216404 300688
rect 216456 300676 216462 300688
rect 287514 300676 287520 300688
rect 216456 300648 287520 300676
rect 216456 300636 216462 300648
rect 287514 300636 287520 300648
rect 287572 300636 287578 300688
rect 213454 300568 213460 300620
rect 213512 300608 213518 300620
rect 284294 300608 284300 300620
rect 213512 300580 284300 300608
rect 213512 300568 213518 300580
rect 284294 300568 284300 300580
rect 284352 300568 284358 300620
rect 214374 300500 214380 300552
rect 214432 300540 214438 300552
rect 286134 300540 286140 300552
rect 214432 300512 286140 300540
rect 214432 300500 214438 300512
rect 286134 300500 286140 300512
rect 286192 300500 286198 300552
rect 305362 300500 305368 300552
rect 305420 300540 305426 300552
rect 375374 300540 375380 300552
rect 305420 300512 375380 300540
rect 305420 300500 305426 300512
rect 375374 300500 375380 300512
rect 375432 300500 375438 300552
rect 217042 300432 217048 300484
rect 217100 300472 217106 300484
rect 349246 300472 349252 300484
rect 217100 300444 349252 300472
rect 217100 300432 217106 300444
rect 349246 300432 349252 300444
rect 349304 300432 349310 300484
rect 210786 300364 210792 300416
rect 210844 300404 210850 300416
rect 346946 300404 346952 300416
rect 210844 300376 346952 300404
rect 210844 300364 210850 300376
rect 346946 300364 346952 300376
rect 347004 300364 347010 300416
rect 210694 300296 210700 300348
rect 210752 300336 210758 300348
rect 349154 300336 349160 300348
rect 210752 300308 349160 300336
rect 210752 300296 210758 300308
rect 349154 300296 349160 300308
rect 349212 300296 349218 300348
rect 212166 300228 212172 300280
rect 212224 300268 212230 300280
rect 284386 300268 284392 300280
rect 212224 300240 284392 300268
rect 212224 300228 212230 300240
rect 284386 300228 284392 300240
rect 284444 300228 284450 300280
rect 337194 300228 337200 300280
rect 337252 300268 337258 300280
rect 542354 300268 542360 300280
rect 337252 300240 542360 300268
rect 337252 300228 337258 300240
rect 542354 300228 542360 300240
rect 542412 300228 542418 300280
rect 211062 300160 211068 300212
rect 211120 300200 211126 300212
rect 284478 300200 284484 300212
rect 211120 300172 284484 300200
rect 211120 300160 211126 300172
rect 284478 300160 284484 300172
rect 284536 300160 284542 300212
rect 339402 300160 339408 300212
rect 339460 300200 339466 300212
rect 553394 300200 553400 300212
rect 339460 300172 553400 300200
rect 339460 300160 339466 300172
rect 553394 300160 553400 300172
rect 553452 300160 553458 300212
rect 209682 300092 209688 300144
rect 209740 300132 209746 300144
rect 284662 300132 284668 300144
rect 209740 300104 284668 300132
rect 209740 300092 209746 300104
rect 284662 300092 284668 300104
rect 284720 300092 284726 300144
rect 339862 300092 339868 300144
rect 339920 300132 339926 300144
rect 556154 300132 556160 300144
rect 339920 300104 556160 300132
rect 339920 300092 339926 300104
rect 556154 300092 556160 300104
rect 556212 300092 556218 300144
rect 216490 300024 216496 300076
rect 216548 300064 216554 300076
rect 285950 300064 285956 300076
rect 216548 300036 285956 300064
rect 216548 300024 216554 300036
rect 285950 300024 285956 300036
rect 286008 300024 286014 300076
rect 219342 299956 219348 300008
rect 219400 299996 219406 300008
rect 287238 299996 287244 300008
rect 219400 299968 287244 299996
rect 219400 299956 219406 299968
rect 287238 299956 287244 299968
rect 287296 299956 287302 300008
rect 217778 299888 217784 299940
rect 217836 299928 217842 299940
rect 285306 299928 285312 299940
rect 217836 299900 285312 299928
rect 217836 299888 217842 299900
rect 285306 299888 285312 299900
rect 285364 299888 285370 299940
rect 304442 298936 304448 298988
rect 304500 298976 304506 298988
rect 372614 298976 372620 298988
rect 304500 298948 372620 298976
rect 304500 298936 304506 298948
rect 372614 298936 372620 298948
rect 372672 298936 372678 298988
rect 335262 298868 335268 298920
rect 335320 298908 335326 298920
rect 531314 298908 531320 298920
rect 335320 298880 531320 298908
rect 335320 298868 335326 298880
rect 531314 298868 531320 298880
rect 531372 298868 531378 298920
rect 335814 298800 335820 298852
rect 335872 298840 335878 298852
rect 535454 298840 535460 298852
rect 335872 298812 535460 298840
rect 335872 298800 335878 298812
rect 535454 298800 535460 298812
rect 535512 298800 535518 298852
rect 335722 298732 335728 298784
rect 335780 298772 335786 298784
rect 539594 298772 539600 298784
rect 335780 298744 539600 298772
rect 335780 298732 335786 298744
rect 539594 298732 539600 298744
rect 539652 298732 539658 298784
rect 323578 297576 323584 297628
rect 323636 297616 323642 297628
rect 465074 297616 465080 297628
rect 323636 297588 465080 297616
rect 323636 297576 323642 297588
rect 465074 297576 465080 297588
rect 465132 297576 465138 297628
rect 330110 297508 330116 297560
rect 330168 297548 330174 297560
rect 506474 297548 506480 297560
rect 330168 297520 506480 297548
rect 330168 297508 330174 297520
rect 506474 297508 506480 297520
rect 506532 297508 506538 297560
rect 331674 297440 331680 297492
rect 331732 297480 331738 297492
rect 510614 297480 510620 297492
rect 331732 297452 510620 297480
rect 331732 297440 331738 297452
rect 510614 297440 510620 297452
rect 510672 297440 510678 297492
rect 333882 297372 333888 297424
rect 333940 297412 333946 297424
rect 524414 297412 524420 297424
rect 333940 297384 524420 297412
rect 333940 297372 333946 297384
rect 524414 297372 524420 297384
rect 524472 297372 524478 297424
rect 217594 296284 217600 296336
rect 217652 296324 217658 296336
rect 343634 296324 343640 296336
rect 217652 296296 343640 296324
rect 217652 296284 217658 296296
rect 343634 296284 343640 296296
rect 343692 296284 343698 296336
rect 218698 296216 218704 296268
rect 218756 296256 218762 296268
rect 347866 296256 347872 296268
rect 218756 296228 347872 296256
rect 218756 296216 218762 296228
rect 347866 296216 347872 296228
rect 347924 296216 347930 296268
rect 327534 296148 327540 296200
rect 327592 296188 327598 296200
rect 492674 296188 492680 296200
rect 327592 296160 492680 296188
rect 327592 296148 327598 296160
rect 492674 296148 492680 296160
rect 492732 296148 492738 296200
rect 328914 296080 328920 296132
rect 328972 296120 328978 296132
rect 499574 296120 499580 296132
rect 328972 296092 499580 296120
rect 328972 296080 328978 296092
rect 499574 296080 499580 296092
rect 499632 296080 499638 296132
rect 330018 296012 330024 296064
rect 330076 296052 330082 296064
rect 503714 296052 503720 296064
rect 330076 296024 503720 296052
rect 330076 296012 330082 296024
rect 503714 296012 503720 296024
rect 503772 296012 503778 296064
rect 341242 295944 341248 295996
rect 341300 295984 341306 295996
rect 567194 295984 567200 295996
rect 341300 295956 567200 295984
rect 341300 295944 341306 295956
rect 567194 295944 567200 295956
rect 567252 295944 567258 295996
rect 325970 294788 325976 294840
rect 326028 294828 326034 294840
rect 481634 294828 481640 294840
rect 326028 294800 481640 294828
rect 326028 294788 326034 294800
rect 481634 294788 481640 294800
rect 481692 294788 481698 294840
rect 325878 294720 325884 294772
rect 325936 294760 325942 294772
rect 485774 294760 485780 294772
rect 325936 294732 485780 294760
rect 325936 294720 325942 294732
rect 485774 294720 485780 294732
rect 485832 294720 485838 294772
rect 327442 294652 327448 294704
rect 327500 294692 327506 294704
rect 489914 294692 489920 294704
rect 327500 294664 489920 294692
rect 327500 294652 327506 294664
rect 489914 294652 489920 294664
rect 489972 294652 489978 294704
rect 124214 294584 124220 294636
rect 124272 294624 124278 294636
rect 255682 294624 255688 294636
rect 124272 294596 255688 294624
rect 124272 294584 124278 294596
rect 255682 294584 255688 294596
rect 255740 294584 255746 294636
rect 338482 294584 338488 294636
rect 338540 294624 338546 294636
rect 549254 294624 549260 294636
rect 338540 294596 549260 294624
rect 338540 294584 338546 294596
rect 549254 294584 549260 294596
rect 549312 294584 549318 294636
rect 321922 293428 321928 293480
rect 321980 293468 321986 293480
rect 466454 293468 466460 293480
rect 321980 293440 466460 293468
rect 321980 293428 321986 293440
rect 466454 293428 466460 293440
rect 466512 293428 466518 293480
rect 117314 293360 117320 293412
rect 117372 293400 117378 293412
rect 254302 293400 254308 293412
rect 117372 293372 254308 293400
rect 117372 293360 117378 293372
rect 254302 293360 254308 293372
rect 254360 293360 254366 293412
rect 323302 293360 323308 293412
rect 323360 293400 323366 293412
rect 473354 293400 473360 293412
rect 323360 293372 473360 293400
rect 323360 293360 323366 293372
rect 473354 293360 473360 293372
rect 473412 293360 473418 293412
rect 110414 293292 110420 293344
rect 110472 293332 110478 293344
rect 252922 293332 252928 293344
rect 110472 293304 252928 293332
rect 110472 293292 110478 293304
rect 252922 293292 252928 293304
rect 252980 293292 252986 293344
rect 324682 293292 324688 293344
rect 324740 293332 324746 293344
rect 477494 293332 477500 293344
rect 324740 293304 477500 293332
rect 324740 293292 324746 293304
rect 477494 293292 477500 293304
rect 477552 293292 477558 293344
rect 102134 293224 102140 293276
rect 102192 293264 102198 293276
rect 251174 293264 251180 293276
rect 102192 293236 251180 293264
rect 102192 293224 102198 293236
rect 251174 293224 251180 293236
rect 251232 293224 251238 293276
rect 328822 293224 328828 293276
rect 328880 293264 328886 293276
rect 496814 293264 496820 293276
rect 328880 293236 496820 293264
rect 328880 293224 328886 293236
rect 496814 293224 496820 293236
rect 496872 293224 496878 293276
rect 315022 292000 315028 292052
rect 315080 292040 315086 292052
rect 431954 292040 431960 292052
rect 315080 292012 431960 292040
rect 315080 292000 315086 292012
rect 431954 292000 431960 292012
rect 432012 292000 432018 292052
rect 95234 291932 95240 291984
rect 95292 291972 95298 291984
rect 250162 291972 250168 291984
rect 95292 291944 250168 291972
rect 95292 291932 95298 291944
rect 250162 291932 250168 291944
rect 250220 291932 250226 291984
rect 320634 291932 320640 291984
rect 320692 291972 320698 291984
rect 459554 291972 459560 291984
rect 320692 291944 459560 291972
rect 320692 291932 320698 291944
rect 459554 291932 459560 291944
rect 459612 291932 459618 291984
rect 92474 291864 92480 291916
rect 92532 291904 92538 291916
rect 249794 291904 249800 291916
rect 92532 291876 249800 291904
rect 92532 291864 92538 291876
rect 249794 291864 249800 291876
rect 249852 291864 249858 291916
rect 321830 291864 321836 291916
rect 321888 291904 321894 291916
rect 463694 291904 463700 291916
rect 321888 291876 463700 291904
rect 321888 291864 321894 291876
rect 463694 291864 463700 291876
rect 463752 291864 463758 291916
rect 88334 291796 88340 291848
rect 88392 291836 88398 291848
rect 248414 291836 248420 291848
rect 88392 291808 248420 291836
rect 88392 291796 88398 291808
rect 248414 291796 248420 291808
rect 248472 291796 248478 291848
rect 323210 291796 323216 291848
rect 323268 291836 323274 291848
rect 470594 291836 470600 291848
rect 323268 291808 470600 291836
rect 323268 291796 323274 291808
rect 470594 291796 470600 291808
rect 470652 291796 470658 291848
rect 106918 290640 106924 290692
rect 106976 290680 106982 290692
rect 248782 290680 248788 290692
rect 106976 290652 248788 290680
rect 106976 290640 106982 290652
rect 248782 290640 248788 290652
rect 248840 290640 248846 290692
rect 312170 290640 312176 290692
rect 312228 290680 312234 290692
rect 414014 290680 414020 290692
rect 312228 290652 414020 290680
rect 312228 290640 312234 290652
rect 414014 290640 414020 290652
rect 414072 290640 414078 290692
rect 81434 290572 81440 290624
rect 81492 290612 81498 290624
rect 247402 290612 247408 290624
rect 81492 290584 247408 290612
rect 81492 290572 81498 290584
rect 247402 290572 247408 290584
rect 247460 290572 247466 290624
rect 313550 290572 313556 290624
rect 313608 290612 313614 290624
rect 423674 290612 423680 290624
rect 313608 290584 423680 290612
rect 313608 290572 313614 290584
rect 423674 290572 423680 290584
rect 423732 290572 423738 290624
rect 77294 290504 77300 290556
rect 77352 290544 77358 290556
rect 247494 290544 247500 290556
rect 77352 290516 247500 290544
rect 77352 290504 77358 290516
rect 247494 290504 247500 290516
rect 247552 290504 247558 290556
rect 314930 290504 314936 290556
rect 314988 290544 314994 290556
rect 427814 290544 427820 290556
rect 314988 290516 427820 290544
rect 314988 290504 314994 290516
rect 427814 290504 427820 290516
rect 427872 290504 427878 290556
rect 74534 290436 74540 290488
rect 74592 290476 74598 290488
rect 246114 290476 246120 290488
rect 74592 290448 246120 290476
rect 74592 290436 74598 290448
rect 246114 290436 246120 290448
rect 246172 290436 246178 290488
rect 316402 290436 316408 290488
rect 316460 290476 316466 290488
rect 438854 290476 438860 290488
rect 316460 290448 438860 290476
rect 316460 290436 316466 290448
rect 438854 290436 438860 290448
rect 438912 290436 438918 290488
rect 122834 289280 122840 289332
rect 122892 289320 122898 289332
rect 255590 289320 255596 289332
rect 122892 289292 255596 289320
rect 122892 289280 122898 289292
rect 255590 289280 255596 289292
rect 255648 289280 255654 289332
rect 309410 289280 309416 289332
rect 309468 289320 309474 289332
rect 402974 289320 402980 289332
rect 309468 289292 402980 289320
rect 309468 289280 309474 289292
rect 402974 289280 402980 289292
rect 403032 289280 403038 289332
rect 118694 289212 118700 289264
rect 118752 289252 118758 289264
rect 255498 289252 255504 289264
rect 118752 289224 255504 289252
rect 118752 289212 118758 289224
rect 255498 289212 255504 289224
rect 255556 289212 255562 289264
rect 310698 289212 310704 289264
rect 310756 289252 310762 289264
rect 407206 289252 407212 289264
rect 310756 289224 407212 289252
rect 310756 289212 310762 289224
rect 407206 289212 407212 289224
rect 407264 289212 407270 289264
rect 115934 289144 115940 289196
rect 115992 289184 115998 289196
rect 254210 289184 254216 289196
rect 115992 289156 254216 289184
rect 115992 289144 115998 289156
rect 254210 289144 254216 289156
rect 254268 289144 254274 289196
rect 310790 289144 310796 289196
rect 310848 289184 310854 289196
rect 409874 289184 409880 289196
rect 310848 289156 409880 289184
rect 310848 289144 310854 289156
rect 409874 289144 409880 289156
rect 409932 289144 409938 289196
rect 70394 289076 70400 289128
rect 70452 289116 70458 289128
rect 246022 289116 246028 289128
rect 70452 289088 246028 289116
rect 70452 289076 70458 289088
rect 246022 289076 246028 289088
rect 246080 289076 246086 289128
rect 313458 289076 313464 289128
rect 313516 289116 313522 289128
rect 420914 289116 420920 289128
rect 313516 289088 420920 289116
rect 313516 289076 313522 289088
rect 420914 289076 420920 289088
rect 420972 289076 420978 289128
rect 111794 287920 111800 287972
rect 111852 287960 111858 287972
rect 254118 287960 254124 287972
rect 111852 287932 254124 287960
rect 111852 287920 111858 287932
rect 254118 287920 254124 287932
rect 254176 287920 254182 287972
rect 109034 287852 109040 287904
rect 109092 287892 109098 287904
rect 252738 287892 252744 287904
rect 109092 287864 252744 287892
rect 109092 287852 109098 287864
rect 252738 287852 252744 287864
rect 252796 287852 252802 287904
rect 308030 287852 308036 287904
rect 308088 287892 308094 287904
rect 391934 287892 391940 287904
rect 308088 287864 391940 287892
rect 308088 287852 308094 287864
rect 391934 287852 391940 287864
rect 391992 287852 391998 287904
rect 104894 287784 104900 287836
rect 104952 287824 104958 287836
rect 252830 287824 252836 287836
rect 104952 287796 252836 287824
rect 104952 287784 104958 287796
rect 252830 287784 252836 287796
rect 252888 287784 252894 287836
rect 307938 287784 307944 287836
rect 307996 287824 308002 287836
rect 396074 287824 396080 287836
rect 307996 287796 396080 287824
rect 307996 287784 308002 287796
rect 396074 287784 396080 287796
rect 396132 287784 396138 287836
rect 63494 287716 63500 287768
rect 63552 287756 63558 287768
rect 244642 287756 244648 287768
rect 63552 287728 244648 287756
rect 63552 287716 63558 287728
rect 244642 287716 244648 287728
rect 244700 287716 244706 287768
rect 309318 287716 309324 287768
rect 309376 287756 309382 287768
rect 398834 287756 398840 287768
rect 309376 287728 398840 287756
rect 309376 287716 309382 287728
rect 398834 287716 398840 287728
rect 398892 287716 398898 287768
rect 38654 287648 38660 287700
rect 38712 287688 38718 287700
rect 239122 287688 239128 287700
rect 38712 287660 239128 287688
rect 38712 287648 38718 287660
rect 239122 287648 239128 287660
rect 239180 287648 239186 287700
rect 312078 287648 312084 287700
rect 312136 287688 312142 287700
rect 416774 287688 416780 287700
rect 312136 287660 416780 287688
rect 312136 287648 312142 287660
rect 416774 287648 416780 287660
rect 416832 287648 416838 287700
rect 102226 286492 102232 286544
rect 102284 286532 102290 286544
rect 251450 286532 251456 286544
rect 102284 286504 251456 286532
rect 102284 286492 102290 286504
rect 251450 286492 251456 286504
rect 251508 286492 251514 286544
rect 303890 286492 303896 286544
rect 303948 286532 303954 286544
rect 373994 286532 374000 286544
rect 303948 286504 374000 286532
rect 303948 286492 303954 286504
rect 373994 286492 374000 286504
rect 374052 286492 374058 286544
rect 97994 286424 98000 286476
rect 98052 286464 98058 286476
rect 251542 286464 251548 286476
rect 98052 286436 251548 286464
rect 98052 286424 98058 286436
rect 251542 286424 251548 286436
rect 251600 286424 251606 286476
rect 305270 286424 305276 286476
rect 305328 286464 305334 286476
rect 378134 286464 378140 286476
rect 305328 286436 378140 286464
rect 305328 286424 305334 286436
rect 378134 286424 378140 286436
rect 378192 286424 378198 286476
rect 93854 286356 93860 286408
rect 93912 286396 93918 286408
rect 250070 286396 250076 286408
rect 93912 286368 250076 286396
rect 93912 286356 93918 286368
rect 250070 286356 250076 286368
rect 250128 286356 250134 286408
rect 306650 286356 306656 286408
rect 306708 286396 306714 286408
rect 389174 286396 389180 286408
rect 306708 286368 389180 286396
rect 306708 286356 306714 286368
rect 389174 286356 389180 286368
rect 389232 286356 389238 286408
rect 54478 286288 54484 286340
rect 54536 286328 54542 286340
rect 241974 286328 241980 286340
rect 54536 286300 241980 286328
rect 54536 286288 54542 286300
rect 241974 286288 241980 286300
rect 242032 286288 242038 286340
rect 343910 286288 343916 286340
rect 343968 286328 343974 286340
rect 576854 286328 576860 286340
rect 343968 286300 576860 286328
rect 343968 286288 343974 286300
rect 576854 286288 576860 286300
rect 576912 286288 576918 286340
rect 118786 285200 118792 285252
rect 118844 285240 118850 285252
rect 255406 285240 255412 285252
rect 118844 285212 255412 285240
rect 118844 285200 118850 285212
rect 255406 285200 255412 285212
rect 255464 285200 255470 285252
rect 303798 285200 303804 285252
rect 303856 285240 303862 285252
rect 371234 285240 371240 285252
rect 303856 285212 371240 285240
rect 303856 285200 303862 285212
rect 371234 285200 371240 285212
rect 371292 285200 371298 285252
rect 114554 285132 114560 285184
rect 114612 285172 114618 285184
rect 254394 285172 254400 285184
rect 114612 285144 254400 285172
rect 114612 285132 114618 285144
rect 254394 285132 254400 285144
rect 254452 285132 254458 285184
rect 319254 285132 319260 285184
rect 319312 285172 319318 285184
rect 447134 285172 447140 285184
rect 319312 285144 447140 285172
rect 319312 285132 319318 285144
rect 447134 285132 447140 285144
rect 447192 285132 447198 285184
rect 110506 285064 110512 285116
rect 110564 285104 110570 285116
rect 254026 285104 254032 285116
rect 110564 285076 254032 285104
rect 110564 285064 110570 285076
rect 254026 285064 254032 285076
rect 254084 285064 254090 285116
rect 342714 285064 342720 285116
rect 342772 285104 342778 285116
rect 552658 285104 552664 285116
rect 342772 285076 552664 285104
rect 342772 285064 342778 285076
rect 552658 285064 552664 285076
rect 552716 285064 552722 285116
rect 91094 284996 91100 285048
rect 91152 285036 91158 285048
rect 249978 285036 249984 285048
rect 91152 285008 249984 285036
rect 91152 284996 91158 285008
rect 249978 284996 249984 285008
rect 250036 284996 250042 285048
rect 341150 284996 341156 285048
rect 341208 285036 341214 285048
rect 565814 285036 565820 285048
rect 341208 285008 565820 285036
rect 341208 284996 341214 285008
rect 565814 284996 565820 285008
rect 565872 284996 565878 285048
rect 49694 284928 49700 284980
rect 49752 284968 49758 284980
rect 241882 284968 241888 284980
rect 49752 284940 241888 284968
rect 49752 284928 49758 284940
rect 241882 284928 241888 284940
rect 241940 284928 241946 284980
rect 342622 284928 342628 284980
rect 342680 284968 342686 284980
rect 569954 284968 569960 284980
rect 342680 284940 569960 284968
rect 342680 284928 342686 284940
rect 569954 284928 569960 284940
rect 570012 284928 570018 284980
rect 107654 283840 107660 283892
rect 107712 283880 107718 283892
rect 253014 283880 253020 283892
rect 107712 283852 253020 283880
rect 107712 283840 107718 283852
rect 253014 283840 253020 283852
rect 253072 283840 253078 283892
rect 103514 283772 103520 283824
rect 103572 283812 103578 283824
rect 252646 283812 252652 283824
rect 103572 283784 252652 283812
rect 103572 283772 103578 283784
rect 252646 283772 252652 283784
rect 252704 283772 252710 283824
rect 334342 283772 334348 283824
rect 334400 283812 334406 283824
rect 528554 283812 528560 283824
rect 334400 283784 528560 283812
rect 334400 283772 334406 283784
rect 528554 283772 528560 283784
rect 528612 283772 528618 283824
rect 100754 283704 100760 283756
rect 100812 283744 100818 283756
rect 251358 283744 251364 283756
rect 100812 283716 251364 283744
rect 100812 283704 100818 283716
rect 251358 283704 251364 283716
rect 251416 283704 251422 283756
rect 339770 283704 339776 283756
rect 339828 283744 339834 283756
rect 538950 283744 538956 283756
rect 339828 283716 538956 283744
rect 339828 283704 339834 283716
rect 538950 283704 538956 283716
rect 539008 283704 539014 283756
rect 77386 283636 77392 283688
rect 77444 283676 77450 283688
rect 247310 283676 247316 283688
rect 77444 283648 247316 283676
rect 77444 283636 77450 283648
rect 247310 283636 247316 283648
rect 247368 283636 247374 283688
rect 338298 283636 338304 283688
rect 338356 283676 338362 283688
rect 547874 283676 547880 283688
rect 338356 283648 547880 283676
rect 338356 283636 338362 283648
rect 547874 283636 547880 283648
rect 547932 283636 547938 283688
rect 31754 283568 31760 283620
rect 31812 283608 31818 283620
rect 237742 283608 237748 283620
rect 31812 283580 237748 283608
rect 31812 283568 31818 283580
rect 237742 283568 237748 283580
rect 237800 283568 237806 283620
rect 338390 283568 338396 283620
rect 338448 283608 338454 283620
rect 552014 283608 552020 283620
rect 338448 283580 552020 283608
rect 338448 283568 338454 283580
rect 552014 283568 552020 283580
rect 552072 283568 552078 283620
rect 160094 282412 160100 282464
rect 160152 282452 160158 282464
rect 262490 282452 262496 282464
rect 160152 282424 262496 282452
rect 160152 282412 160158 282424
rect 262490 282412 262496 282424
rect 262548 282412 262554 282464
rect 155954 282344 155960 282396
rect 156012 282384 156018 282396
rect 262582 282384 262588 282396
rect 156012 282356 262588 282384
rect 156012 282344 156018 282356
rect 262582 282344 262588 282356
rect 262640 282344 262646 282396
rect 317782 282344 317788 282396
rect 317840 282384 317846 282396
rect 442994 282384 443000 282396
rect 317840 282356 443000 282384
rect 317840 282344 317846 282356
rect 442994 282344 443000 282356
rect 443052 282344 443058 282396
rect 96614 282276 96620 282328
rect 96672 282316 96678 282328
rect 251266 282316 251272 282328
rect 96672 282288 251272 282316
rect 96672 282276 96678 282288
rect 251266 282276 251272 282288
rect 251324 282276 251330 282328
rect 333054 282276 333060 282328
rect 333112 282316 333118 282328
rect 520274 282316 520280 282328
rect 333112 282288 520280 282316
rect 333112 282276 333118 282288
rect 520274 282276 520280 282288
rect 520332 282276 520338 282328
rect 73154 282208 73160 282260
rect 73212 282248 73218 282260
rect 245930 282248 245936 282260
rect 73212 282220 245936 282248
rect 73212 282208 73218 282220
rect 245930 282208 245936 282220
rect 245988 282208 245994 282260
rect 334250 282208 334256 282260
rect 334308 282248 334314 282260
rect 527174 282248 527180 282260
rect 334308 282220 527180 282248
rect 334308 282208 334314 282220
rect 527174 282208 527180 282220
rect 527232 282208 527238 282260
rect 43530 282140 43536 282192
rect 43588 282180 43594 282192
rect 240502 282180 240508 282192
rect 43588 282152 240508 282180
rect 43588 282140 43594 282152
rect 240502 282140 240508 282152
rect 240560 282140 240566 282192
rect 334158 282140 334164 282192
rect 334216 282180 334222 282192
rect 531406 282180 531412 282192
rect 334216 282152 531412 282180
rect 334216 282140 334222 282152
rect 531406 282140 531412 282152
rect 531464 282140 531470 282192
rect 218422 281120 218428 281172
rect 218480 281160 218486 281172
rect 273714 281160 273720 281172
rect 218480 281132 273720 281160
rect 218480 281120 218486 281132
rect 273714 281120 273720 281132
rect 273772 281120 273778 281172
rect 205634 281052 205640 281104
rect 205692 281092 205698 281104
rect 272242 281092 272248 281104
rect 205692 281064 272248 281092
rect 205692 281052 205698 281064
rect 272242 281052 272248 281064
rect 272300 281052 272306 281104
rect 198734 280984 198740 281036
rect 198792 281024 198798 281036
rect 270954 281024 270960 281036
rect 198792 280996 270960 281024
rect 198792 280984 198798 280996
rect 270954 280984 270960 280996
rect 271012 280984 271018 281036
rect 329926 280984 329932 281036
rect 329984 281024 329990 281036
rect 509234 281024 509240 281036
rect 329984 280996 509240 281024
rect 329984 280984 329990 280996
rect 509234 280984 509240 280996
rect 509292 280984 509298 281036
rect 151814 280916 151820 280968
rect 151872 280956 151878 280968
rect 261386 280956 261392 280968
rect 151872 280928 261392 280956
rect 151872 280916 151878 280928
rect 261386 280916 261392 280928
rect 261444 280916 261450 280968
rect 331490 280916 331496 280968
rect 331548 280956 331554 280968
rect 513374 280956 513380 280968
rect 331548 280928 513380 280956
rect 331548 280916 331554 280928
rect 513374 280916 513380 280928
rect 513432 280916 513438 280968
rect 149054 280848 149060 280900
rect 149112 280888 149118 280900
rect 261294 280888 261300 280900
rect 149112 280860 261300 280888
rect 149112 280848 149118 280860
rect 261294 280848 261300 280860
rect 261352 280848 261358 280900
rect 331582 280848 331588 280900
rect 331640 280888 331646 280900
rect 516134 280888 516140 280900
rect 331640 280860 516140 280888
rect 331640 280848 331646 280860
rect 516134 280848 516140 280860
rect 516192 280848 516198 280900
rect 36538 280780 36544 280832
rect 36596 280820 36602 280832
rect 239030 280820 239036 280832
rect 36596 280792 239036 280820
rect 36596 280780 36602 280792
rect 239030 280780 239036 280792
rect 239088 280780 239094 280832
rect 341058 280780 341064 280832
rect 341116 280820 341122 280832
rect 563054 280820 563060 280832
rect 341116 280792 563060 280820
rect 341116 280780 341122 280792
rect 563054 280780 563060 280792
rect 563112 280780 563118 280832
rect 196618 279692 196624 279744
rect 196676 279732 196682 279744
rect 269482 279732 269488 279744
rect 196676 279704 269488 279732
rect 196676 279692 196682 279704
rect 269482 279692 269488 279704
rect 269540 279692 269546 279744
rect 191834 279624 191840 279676
rect 191892 279664 191898 279676
rect 269574 279664 269580 279676
rect 191892 279636 269580 279664
rect 191892 279624 191898 279636
rect 269574 279624 269580 279636
rect 269632 279624 269638 279676
rect 328638 279624 328644 279676
rect 328696 279664 328702 279676
rect 498194 279664 498200 279676
rect 328696 279636 498200 279664
rect 328696 279624 328702 279636
rect 498194 279624 498200 279636
rect 498252 279624 498258 279676
rect 187694 279556 187700 279608
rect 187752 279596 187758 279608
rect 268194 279596 268200 279608
rect 187752 279568 268200 279596
rect 187752 279556 187758 279568
rect 268194 279556 268200 279568
rect 268252 279556 268258 279608
rect 328730 279556 328736 279608
rect 328788 279596 328794 279608
rect 502334 279596 502340 279608
rect 328788 279568 502340 279596
rect 328788 279556 328794 279568
rect 502334 279556 502340 279568
rect 502392 279556 502398 279608
rect 144914 279488 144920 279540
rect 144972 279528 144978 279540
rect 259914 279528 259920 279540
rect 144972 279500 259920 279528
rect 144972 279488 144978 279500
rect 259914 279488 259920 279500
rect 259972 279488 259978 279540
rect 329834 279488 329840 279540
rect 329892 279528 329898 279540
rect 506566 279528 506572 279540
rect 329892 279500 506572 279528
rect 329892 279488 329898 279500
rect 506566 279488 506572 279500
rect 506624 279488 506630 279540
rect 69014 279420 69020 279472
rect 69072 279460 69078 279472
rect 245838 279460 245844 279472
rect 69072 279432 245844 279460
rect 69072 279420 69078 279432
rect 245838 279420 245844 279432
rect 245896 279420 245902 279472
rect 339678 279420 339684 279472
rect 339736 279460 339742 279472
rect 556246 279460 556252 279472
rect 339736 279432 556252 279460
rect 339736 279420 339742 279432
rect 556246 279420 556252 279432
rect 556304 279420 556310 279472
rect 184934 278264 184940 278316
rect 184992 278304 184998 278316
rect 268102 278304 268108 278316
rect 184992 278276 268108 278304
rect 184992 278264 184998 278276
rect 268102 278264 268108 278276
rect 268160 278264 268166 278316
rect 180794 278196 180800 278248
rect 180852 278236 180858 278248
rect 266722 278236 266728 278248
rect 180852 278208 266728 278236
rect 180852 278196 180858 278208
rect 266722 278196 266728 278208
rect 266780 278196 266786 278248
rect 325786 278196 325792 278248
rect 325844 278236 325850 278248
rect 488534 278236 488540 278248
rect 325844 278208 488540 278236
rect 325844 278196 325850 278208
rect 488534 278196 488540 278208
rect 488592 278196 488598 278248
rect 176654 278128 176660 278180
rect 176712 278168 176718 278180
rect 266630 278168 266636 278180
rect 176712 278140 266636 278168
rect 176712 278128 176718 278140
rect 266630 278128 266636 278140
rect 266688 278128 266694 278180
rect 327350 278128 327356 278180
rect 327408 278168 327414 278180
rect 491294 278168 491300 278180
rect 327408 278140 491300 278168
rect 327408 278128 327414 278140
rect 491294 278128 491300 278140
rect 491352 278128 491358 278180
rect 142154 278060 142160 278112
rect 142212 278100 142218 278112
rect 259822 278100 259828 278112
rect 142212 278072 259828 278100
rect 142212 278060 142218 278072
rect 259822 278060 259828 278072
rect 259880 278060 259886 278112
rect 327258 278060 327264 278112
rect 327316 278100 327322 278112
rect 495434 278100 495440 278112
rect 327316 278072 495440 278100
rect 327316 278060 327322 278072
rect 495434 278060 495440 278072
rect 495492 278060 495498 278112
rect 66254 277992 66260 278044
rect 66312 278032 66318 278044
rect 244550 278032 244556 278044
rect 66312 278004 244556 278032
rect 66312 277992 66318 278004
rect 244550 277992 244556 278004
rect 244608 277992 244614 278044
rect 337102 277992 337108 278044
rect 337160 278032 337166 278044
rect 545114 278032 545120 278044
rect 337160 278004 545120 278032
rect 337160 277992 337166 278004
rect 545114 277992 545120 278004
rect 545172 277992 545178 278044
rect 173894 276904 173900 276956
rect 173952 276944 173958 276956
rect 265342 276944 265348 276956
rect 173952 276916 265348 276944
rect 173952 276904 173958 276916
rect 265342 276904 265348 276916
rect 265400 276904 265406 276956
rect 169754 276836 169760 276888
rect 169812 276876 169818 276888
rect 265434 276876 265440 276888
rect 169812 276848 265440 276876
rect 169812 276836 169818 276848
rect 265434 276836 265440 276848
rect 265492 276836 265498 276888
rect 316310 276836 316316 276888
rect 316368 276876 316374 276888
rect 437474 276876 437480 276888
rect 316368 276848 437480 276876
rect 316368 276836 316374 276848
rect 437474 276836 437480 276848
rect 437532 276836 437538 276888
rect 61378 276768 61384 276820
rect 61436 276808 61442 276820
rect 243354 276808 243360 276820
rect 61436 276780 243360 276808
rect 61436 276768 61442 276780
rect 243354 276768 243360 276780
rect 243412 276768 243418 276820
rect 319162 276768 319168 276820
rect 319220 276808 319226 276820
rect 451274 276808 451280 276820
rect 319220 276780 451280 276808
rect 319220 276768 319226 276780
rect 451274 276768 451280 276780
rect 451332 276768 451338 276820
rect 62114 276700 62120 276752
rect 62172 276740 62178 276752
rect 244458 276740 244464 276752
rect 62172 276712 244464 276740
rect 62172 276700 62178 276712
rect 244458 276700 244464 276712
rect 244516 276700 244522 276752
rect 320542 276700 320548 276752
rect 320600 276740 320606 276752
rect 455414 276740 455420 276752
rect 320600 276712 455420 276740
rect 320600 276700 320606 276712
rect 455414 276700 455420 276712
rect 455472 276700 455478 276752
rect 26878 276632 26884 276684
rect 26936 276672 26942 276684
rect 236270 276672 236276 276684
rect 26936 276644 236276 276672
rect 26936 276632 26942 276644
rect 236270 276632 236276 276644
rect 236328 276632 236334 276684
rect 321738 276632 321744 276684
rect 321796 276672 321802 276684
rect 462314 276672 462320 276684
rect 321796 276644 462320 276672
rect 321796 276632 321802 276644
rect 462314 276632 462320 276644
rect 462372 276632 462378 276684
rect 313366 275476 313372 275528
rect 313424 275516 313430 275528
rect 419534 275516 419540 275528
rect 313424 275488 419540 275516
rect 313424 275476 313430 275488
rect 419534 275476 419540 275488
rect 419592 275476 419598 275528
rect 166994 275408 167000 275460
rect 167052 275448 167058 275460
rect 264054 275448 264060 275460
rect 167052 275420 264060 275448
rect 167052 275408 167058 275420
rect 264054 275408 264060 275420
rect 264112 275408 264118 275460
rect 314838 275408 314844 275460
rect 314896 275448 314902 275460
rect 426434 275448 426440 275460
rect 314896 275420 426440 275448
rect 314896 275408 314902 275420
rect 426434 275408 426440 275420
rect 426492 275408 426498 275460
rect 162854 275340 162860 275392
rect 162912 275380 162918 275392
rect 263962 275380 263968 275392
rect 162912 275352 263968 275380
rect 162912 275340 162918 275352
rect 263962 275340 263968 275352
rect 264020 275340 264026 275392
rect 316218 275340 316224 275392
rect 316276 275380 316282 275392
rect 433334 275380 433340 275392
rect 316276 275352 433340 275380
rect 316276 275340 316282 275352
rect 433334 275340 433340 275352
rect 433392 275340 433398 275392
rect 57238 275272 57244 275324
rect 57296 275312 57302 275324
rect 243262 275312 243268 275324
rect 57296 275284 243268 275312
rect 57296 275272 57302 275284
rect 243262 275272 243268 275284
rect 243320 275272 243326 275324
rect 317690 275272 317696 275324
rect 317748 275312 317754 275324
rect 444374 275312 444380 275324
rect 317748 275284 444380 275312
rect 317748 275272 317754 275284
rect 444374 275272 444380 275284
rect 444432 275272 444438 275324
rect 206278 274184 206284 274236
rect 206336 274224 206342 274236
rect 272058 274224 272064 274236
rect 206336 274196 272064 274224
rect 206336 274184 206342 274196
rect 272058 274184 272064 274196
rect 272116 274184 272122 274236
rect 201494 274116 201500 274168
rect 201552 274156 201558 274168
rect 270862 274156 270868 274168
rect 201552 274128 270868 274156
rect 201552 274116 201558 274128
rect 270862 274116 270868 274128
rect 270920 274116 270926 274168
rect 309226 274116 309232 274168
rect 309284 274156 309290 274168
rect 401594 274156 401600 274168
rect 309284 274128 401600 274156
rect 309284 274116 309290 274128
rect 401594 274116 401600 274128
rect 401652 274116 401658 274168
rect 158714 274048 158720 274100
rect 158772 274088 158778 274100
rect 262398 274088 262404 274100
rect 158772 274060 262404 274088
rect 158772 274048 158778 274060
rect 262398 274048 262404 274060
rect 262456 274048 262462 274100
rect 310606 274048 310612 274100
rect 310664 274088 310670 274100
rect 408494 274088 408500 274100
rect 310664 274060 408500 274088
rect 310664 274048 310670 274060
rect 408494 274048 408500 274060
rect 408552 274048 408558 274100
rect 138014 273980 138020 274032
rect 138072 274020 138078 274032
rect 258350 274020 258356 274032
rect 138072 273992 258356 274020
rect 138072 273980 138078 273992
rect 258350 273980 258356 273992
rect 258408 273980 258414 274032
rect 311986 273980 311992 274032
rect 312044 274020 312050 274032
rect 415486 274020 415492 274032
rect 312044 273992 415492 274020
rect 312044 273980 312050 273992
rect 415486 273980 415492 273992
rect 415544 273980 415550 274032
rect 30374 273912 30380 273964
rect 30432 273952 30438 273964
rect 237650 273952 237656 273964
rect 30432 273924 237656 273952
rect 30432 273912 30438 273924
rect 237650 273912 237656 273924
rect 237708 273912 237714 273964
rect 313274 273912 313280 273964
rect 313332 273952 313338 273964
rect 423766 273952 423772 273964
rect 313332 273924 423772 273952
rect 313332 273912 313338 273924
rect 423766 273912 423772 273924
rect 423824 273912 423830 273964
rect 364978 273164 364984 273216
rect 365036 273204 365042 273216
rect 579614 273204 579620 273216
rect 365036 273176 579620 273204
rect 365036 273164 365042 273176
rect 579614 273164 579620 273176
rect 579672 273164 579678 273216
rect 197354 272824 197360 272876
rect 197412 272864 197418 272876
rect 270770 272864 270776 272876
rect 197412 272836 270776 272864
rect 197412 272824 197418 272836
rect 270770 272824 270776 272836
rect 270828 272824 270834 272876
rect 193214 272756 193220 272808
rect 193272 272796 193278 272808
rect 269298 272796 269304 272808
rect 193272 272768 269304 272796
rect 193272 272756 193278 272768
rect 269298 272756 269304 272768
rect 269356 272756 269362 272808
rect 192478 272688 192484 272740
rect 192536 272728 192542 272740
rect 269390 272728 269396 272740
rect 192536 272700 269396 272728
rect 192536 272688 192542 272700
rect 269390 272688 269396 272700
rect 269448 272688 269454 272740
rect 154574 272620 154580 272672
rect 154632 272660 154638 272672
rect 262306 272660 262312 272672
rect 154632 272632 262312 272660
rect 154632 272620 154638 272632
rect 262306 272620 262312 272632
rect 262364 272620 262370 272672
rect 307754 272620 307760 272672
rect 307812 272660 307818 272672
rect 390554 272660 390560 272672
rect 307812 272632 390560 272660
rect 307812 272620 307818 272632
rect 390554 272620 390560 272632
rect 390612 272620 390618 272672
rect 131114 272552 131120 272604
rect 131172 272592 131178 272604
rect 257154 272592 257160 272604
rect 131172 272564 257160 272592
rect 131172 272552 131178 272564
rect 257154 272552 257160 272564
rect 257212 272552 257218 272604
rect 307846 272552 307852 272604
rect 307904 272592 307910 272604
rect 394694 272592 394700 272604
rect 307904 272564 394700 272592
rect 307904 272552 307910 272564
rect 394694 272552 394700 272564
rect 394752 272552 394758 272604
rect 27614 272484 27620 272536
rect 27672 272524 27678 272536
rect 237558 272524 237564 272536
rect 27672 272496 237564 272524
rect 27672 272484 27678 272496
rect 237558 272484 237564 272496
rect 237616 272484 237622 272536
rect 309134 272484 309140 272536
rect 309192 272524 309198 272536
rect 398926 272524 398932 272536
rect 309192 272496 398932 272524
rect 309192 272484 309198 272496
rect 398926 272484 398932 272496
rect 398984 272484 398990 272536
rect 188338 271464 188344 271516
rect 188396 271504 188402 271516
rect 268010 271504 268016 271516
rect 188396 271476 268016 271504
rect 188396 271464 188402 271476
rect 268010 271464 268016 271476
rect 268068 271464 268074 271516
rect 183554 271396 183560 271448
rect 183612 271436 183618 271448
rect 267918 271436 267924 271448
rect 183612 271408 267924 271436
rect 183612 271396 183618 271408
rect 267918 271396 267924 271408
rect 267976 271396 267982 271448
rect 179414 271328 179420 271380
rect 179472 271368 179478 271380
rect 266538 271368 266544 271380
rect 179472 271340 266544 271368
rect 179472 271328 179478 271340
rect 266538 271328 266544 271340
rect 266596 271328 266602 271380
rect 305178 271328 305184 271380
rect 305236 271368 305242 271380
rect 380894 271368 380900 271380
rect 305236 271340 380900 271368
rect 305236 271328 305242 271340
rect 380894 271328 380900 271340
rect 380952 271328 380958 271380
rect 140774 271260 140780 271312
rect 140832 271300 140838 271312
rect 259730 271300 259736 271312
rect 140832 271272 259736 271300
rect 140832 271260 140838 271272
rect 259730 271260 259736 271272
rect 259788 271260 259794 271312
rect 306558 271260 306564 271312
rect 306616 271300 306622 271312
rect 383654 271300 383660 271312
rect 306616 271272 383660 271300
rect 306616 271260 306622 271272
rect 383654 271260 383660 271272
rect 383712 271260 383718 271312
rect 93946 271192 93952 271244
rect 94004 271232 94010 271244
rect 249886 271232 249892 271244
rect 94004 271204 249892 271232
rect 94004 271192 94010 271204
rect 249886 271192 249892 271204
rect 249944 271192 249950 271244
rect 306466 271192 306472 271244
rect 306524 271232 306530 271244
rect 387794 271232 387800 271244
rect 306524 271204 387800 271232
rect 306524 271192 306530 271204
rect 387794 271192 387800 271204
rect 387852 271192 387858 271244
rect 22094 271124 22100 271176
rect 22152 271164 22158 271176
rect 236178 271164 236184 271176
rect 22152 271136 236184 271164
rect 22152 271124 22158 271136
rect 236178 271124 236184 271136
rect 236236 271124 236242 271176
rect 320450 271124 320456 271176
rect 320508 271164 320514 271176
rect 458174 271164 458180 271176
rect 320508 271136 458180 271164
rect 320508 271124 320514 271136
rect 458174 271124 458180 271136
rect 458232 271124 458238 271176
rect 176746 270104 176752 270156
rect 176804 270144 176810 270156
rect 266446 270144 266452 270156
rect 176804 270116 266452 270144
rect 176804 270104 176810 270116
rect 266446 270104 266452 270116
rect 266504 270104 266510 270156
rect 172514 270036 172520 270088
rect 172572 270076 172578 270088
rect 265250 270076 265256 270088
rect 172572 270048 265256 270076
rect 172572 270036 172578 270048
rect 265250 270036 265256 270048
rect 265308 270036 265314 270088
rect 168374 269968 168380 270020
rect 168432 270008 168438 270020
rect 265158 270008 265164 270020
rect 168432 269980 265164 270008
rect 168432 269968 168438 269980
rect 265158 269968 265164 269980
rect 265216 269968 265222 270020
rect 136634 269900 136640 269952
rect 136692 269940 136698 269952
rect 258258 269940 258264 269952
rect 136692 269912 258264 269940
rect 136692 269900 136698 269912
rect 258258 269900 258264 269912
rect 258316 269900 258322 269952
rect 303614 269900 303620 269952
rect 303672 269940 303678 269952
rect 374086 269940 374092 269952
rect 303672 269912 374092 269940
rect 303672 269900 303678 269912
rect 374086 269900 374092 269912
rect 374144 269900 374150 269952
rect 89714 269832 89720 269884
rect 89772 269872 89778 269884
rect 250254 269872 250260 269884
rect 89772 269844 250260 269872
rect 89772 269832 89778 269844
rect 250254 269832 250260 269844
rect 250312 269832 250318 269884
rect 305086 269832 305092 269884
rect 305144 269872 305150 269884
rect 376754 269872 376760 269884
rect 305144 269844 376760 269872
rect 305144 269832 305150 269844
rect 376754 269832 376760 269844
rect 376812 269832 376818 269884
rect 13814 269764 13820 269816
rect 13872 269804 13878 269816
rect 235074 269804 235080 269816
rect 13872 269776 235080 269804
rect 13872 269764 13878 269776
rect 235074 269764 235080 269776
rect 235132 269764 235138 269816
rect 317598 269764 317604 269816
rect 317656 269804 317662 269816
rect 440326 269804 440332 269816
rect 317656 269776 440332 269804
rect 317656 269764 317662 269776
rect 440326 269764 440332 269776
rect 440384 269764 440390 269816
rect 165614 268608 165620 268660
rect 165672 268648 165678 268660
rect 263870 268648 263876 268660
rect 165672 268620 263876 268648
rect 165672 268608 165678 268620
rect 263870 268608 263876 268620
rect 263928 268608 263934 268660
rect 302510 268608 302516 268660
rect 302568 268648 302574 268660
rect 365714 268648 365720 268660
rect 302568 268620 365720 268648
rect 302568 268608 302574 268620
rect 365714 268608 365720 268620
rect 365772 268608 365778 268660
rect 161474 268540 161480 268592
rect 161532 268580 161538 268592
rect 263778 268580 263784 268592
rect 161532 268552 263784 268580
rect 161532 268540 161538 268552
rect 263778 268540 263784 268552
rect 263836 268540 263842 268592
rect 320358 268540 320364 268592
rect 320416 268580 320422 268592
rect 456794 268580 456800 268592
rect 320416 268552 456800 268580
rect 320416 268540 320422 268552
rect 456794 268540 456800 268552
rect 456852 268540 456858 268592
rect 157334 268472 157340 268524
rect 157392 268512 157398 268524
rect 262674 268512 262680 268524
rect 157392 268484 262680 268512
rect 157392 268472 157398 268484
rect 262674 268472 262680 268484
rect 262732 268472 262738 268524
rect 339586 268472 339592 268524
rect 339644 268512 339650 268524
rect 516778 268512 516784 268524
rect 339644 268484 516784 268512
rect 339644 268472 339650 268484
rect 516778 268472 516784 268484
rect 516836 268472 516842 268524
rect 133874 268404 133880 268456
rect 133932 268444 133938 268456
rect 258166 268444 258172 268456
rect 133932 268416 258172 268444
rect 133932 268404 133938 268416
rect 258166 268404 258172 268416
rect 258224 268404 258230 268456
rect 342530 268404 342536 268456
rect 342588 268444 342594 268456
rect 520918 268444 520924 268456
rect 342588 268416 520924 268444
rect 342588 268404 342594 268416
rect 520918 268404 520924 268416
rect 520976 268404 520982 268456
rect 52454 268336 52460 268388
rect 52512 268376 52518 268388
rect 241790 268376 241796 268388
rect 52512 268348 241796 268376
rect 52512 268336 52518 268348
rect 241790 268336 241796 268348
rect 241848 268336 241854 268388
rect 342438 268336 342444 268388
rect 342496 268376 342502 268388
rect 525058 268376 525064 268388
rect 342496 268348 525064 268376
rect 342496 268336 342502 268348
rect 525058 268336 525064 268348
rect 525116 268336 525122 268388
rect 3326 267656 3332 267708
rect 3384 267696 3390 267708
rect 174538 267696 174544 267708
rect 3384 267668 174544 267696
rect 3384 267656 3390 267668
rect 174538 267656 174544 267668
rect 174596 267656 174602 267708
rect 153194 267180 153200 267232
rect 153252 267220 153258 267232
rect 261202 267220 261208 267232
rect 153252 267192 261208 267220
rect 153252 267180 153258 267192
rect 261202 267180 261208 267192
rect 261260 267180 261266 267232
rect 319070 267180 319076 267232
rect 319128 267220 319134 267232
rect 448514 267220 448520 267232
rect 319128 267192 448520 267220
rect 319128 267180 319134 267192
rect 448514 267180 448520 267192
rect 448572 267180 448578 267232
rect 150434 267112 150440 267164
rect 150492 267152 150498 267164
rect 261110 267152 261116 267164
rect 150492 267124 261116 267152
rect 150492 267112 150498 267124
rect 261110 267112 261116 267124
rect 261168 267112 261174 267164
rect 338206 267112 338212 267164
rect 338264 267152 338270 267164
rect 508498 267152 508504 267164
rect 338264 267124 508504 267152
rect 338264 267112 338270 267124
rect 508498 267112 508504 267124
rect 508556 267112 508562 267164
rect 48314 267044 48320 267096
rect 48372 267084 48378 267096
rect 241698 267084 241704 267096
rect 48372 267056 241704 267084
rect 48372 267044 48378 267056
rect 241698 267044 241704 267056
rect 241756 267044 241762 267096
rect 337010 267044 337016 267096
rect 337068 267084 337074 267096
rect 543734 267084 543740 267096
rect 337068 267056 543740 267084
rect 337068 267044 337074 267056
rect 543734 267044 543740 267056
rect 543792 267044 543798 267096
rect 8294 266976 8300 267028
rect 8352 267016 8358 267028
rect 233510 267016 233516 267028
rect 8352 266988 233516 267016
rect 8352 266976 8358 266988
rect 233510 266976 233516 266988
rect 233568 266976 233574 267028
rect 338114 266976 338120 267028
rect 338172 267016 338178 267028
rect 547966 267016 547972 267028
rect 338172 266988 547972 267016
rect 338172 266976 338178 266988
rect 547966 266976 547972 266988
rect 548024 266976 548030 267028
rect 209774 265956 209780 266008
rect 209832 265996 209838 266008
rect 271966 265996 271972 266008
rect 209832 265968 271972 265996
rect 209832 265956 209838 265968
rect 271966 265956 271972 265968
rect 272024 265956 272030 266008
rect 202874 265888 202880 265940
rect 202932 265928 202938 265940
rect 270678 265928 270684 265940
rect 202932 265900 270684 265928
rect 202932 265888 202938 265900
rect 270678 265888 270684 265900
rect 270736 265888 270742 265940
rect 200114 265820 200120 265872
rect 200172 265860 200178 265872
rect 270586 265860 270592 265872
rect 200172 265832 270592 265860
rect 200172 265820 200178 265832
rect 270586 265820 270592 265832
rect 270644 265820 270650 265872
rect 318978 265820 318984 265872
rect 319036 265860 319042 265872
rect 449894 265860 449900 265872
rect 319036 265832 449900 265860
rect 319036 265820 319042 265832
rect 449894 265820 449900 265832
rect 449952 265820 449958 265872
rect 146294 265752 146300 265804
rect 146352 265792 146358 265804
rect 261018 265792 261024 265804
rect 146352 265764 261024 265792
rect 146352 265752 146358 265764
rect 261018 265752 261024 265764
rect 261076 265752 261082 265804
rect 335630 265752 335636 265804
rect 335688 265792 335694 265804
rect 496078 265792 496084 265804
rect 335688 265764 496084 265792
rect 335688 265752 335694 265764
rect 496078 265752 496084 265764
rect 496136 265752 496142 265804
rect 126974 265684 126980 265736
rect 127032 265724 127038 265736
rect 257062 265724 257068 265736
rect 127032 265696 257068 265724
rect 127032 265684 127038 265696
rect 257062 265684 257068 265696
rect 257120 265684 257126 265736
rect 335538 265684 335544 265736
rect 335596 265724 335602 265736
rect 502978 265724 502984 265736
rect 335596 265696 502984 265724
rect 335596 265684 335602 265696
rect 502978 265684 502984 265696
rect 503036 265684 503042 265736
rect 44174 265616 44180 265668
rect 44232 265656 44238 265668
rect 240410 265656 240416 265668
rect 44232 265628 240416 265656
rect 44232 265616 44238 265628
rect 240410 265616 240416 265628
rect 240468 265616 240474 265668
rect 334066 265616 334072 265668
rect 334124 265656 334130 265668
rect 529934 265656 529940 265668
rect 334124 265628 529940 265656
rect 334124 265616 334130 265628
rect 529934 265616 529940 265628
rect 529992 265616 529998 265668
rect 195974 264528 195980 264580
rect 196032 264568 196038 264580
rect 269114 264568 269120 264580
rect 196032 264540 269120 264568
rect 196032 264528 196038 264540
rect 269114 264528 269120 264540
rect 269172 264528 269178 264580
rect 193306 264460 193312 264512
rect 193364 264500 193370 264512
rect 269206 264500 269212 264512
rect 193364 264472 269212 264500
rect 193364 264460 193370 264472
rect 269206 264460 269212 264472
rect 269264 264460 269270 264512
rect 189074 264392 189080 264444
rect 189132 264432 189138 264444
rect 267826 264432 267832 264444
rect 189132 264404 267832 264432
rect 189132 264392 189138 264404
rect 267826 264392 267832 264404
rect 267884 264392 267890 264444
rect 316126 264392 316132 264444
rect 316184 264432 316190 264444
rect 436094 264432 436100 264444
rect 316184 264404 436100 264432
rect 316184 264392 316190 264404
rect 436094 264392 436100 264404
rect 436152 264392 436158 264444
rect 139394 264324 139400 264376
rect 139452 264364 139458 264376
rect 259638 264364 259644 264376
rect 139452 264336 259644 264364
rect 139452 264324 139458 264336
rect 259638 264324 259644 264336
rect 259696 264324 259702 264376
rect 331398 264324 331404 264376
rect 331456 264364 331462 264376
rect 457438 264364 457444 264376
rect 331456 264336 457444 264364
rect 331456 264324 331462 264336
rect 457438 264324 457444 264336
rect 457496 264324 457502 264376
rect 85574 264256 85580 264308
rect 85632 264296 85638 264308
rect 248690 264296 248696 264308
rect 85632 264268 248696 264296
rect 85632 264256 85638 264268
rect 248690 264256 248696 264268
rect 248748 264256 248754 264308
rect 332870 264256 332876 264308
rect 332928 264296 332934 264308
rect 467098 264296 467104 264308
rect 332928 264268 467104 264296
rect 332928 264256 332934 264268
rect 467098 264256 467104 264268
rect 467156 264256 467162 264308
rect 2774 264188 2780 264240
rect 2832 264228 2838 264240
rect 232130 264228 232136 264240
rect 2832 264200 232136 264228
rect 2832 264188 2838 264200
rect 232130 264188 232136 264200
rect 232188 264188 232194 264240
rect 332962 264188 332968 264240
rect 333020 264228 333026 264240
rect 476758 264228 476764 264240
rect 333020 264200 476764 264228
rect 333020 264188 333026 264200
rect 476758 264188 476764 264200
rect 476816 264188 476822 264240
rect 185026 263100 185032 263152
rect 185084 263140 185090 263152
rect 267734 263140 267740 263152
rect 185084 263112 267740 263140
rect 185084 263100 185090 263112
rect 267734 263100 267740 263112
rect 267792 263100 267798 263152
rect 175274 263032 175280 263084
rect 175332 263072 175338 263084
rect 264974 263072 264980 263084
rect 175332 263044 264980 263072
rect 175332 263032 175338 263044
rect 264974 263032 264980 263044
rect 265032 263032 265038 263084
rect 311894 263032 311900 263084
rect 311952 263072 311958 263084
rect 412634 263072 412640 263084
rect 311952 263044 412640 263072
rect 311952 263032 311958 263044
rect 412634 263032 412640 263044
rect 412692 263032 412698 263084
rect 171134 262964 171140 263016
rect 171192 263004 171198 263016
rect 265066 263004 265072 263016
rect 171192 262976 265072 263004
rect 171192 262964 171198 262976
rect 265066 262964 265072 262976
rect 265124 262964 265130 263016
rect 328546 262964 328552 263016
rect 328604 263004 328610 263016
rect 432598 263004 432604 263016
rect 328604 262976 432604 263004
rect 328604 262964 328610 262976
rect 432598 262964 432604 262976
rect 432656 262964 432662 263016
rect 132494 262896 132500 262948
rect 132552 262936 132558 262948
rect 253198 262936 253204 262948
rect 132552 262908 253204 262936
rect 132552 262896 132558 262908
rect 253198 262896 253204 262908
rect 253256 262896 253262 262948
rect 328454 262896 328460 262948
rect 328512 262936 328518 262948
rect 498286 262936 498292 262948
rect 328512 262908 498292 262936
rect 328512 262896 328518 262908
rect 498286 262896 498292 262908
rect 498344 262896 498350 262948
rect 40034 262828 40040 262880
rect 40092 262868 40098 262880
rect 240318 262868 240324 262880
rect 40092 262840 240324 262868
rect 40092 262828 40098 262840
rect 240318 262828 240324 262840
rect 240376 262828 240382 262880
rect 331306 262828 331312 262880
rect 331364 262868 331370 262880
rect 511994 262868 512000 262880
rect 331364 262840 512000 262868
rect 331364 262828 331370 262840
rect 511994 262828 512000 262840
rect 512052 262828 512058 262880
rect 168466 261740 168472 261792
rect 168524 261780 168530 261792
rect 263686 261780 263692 261792
rect 168524 261752 263692 261780
rect 168524 261740 168530 261752
rect 263686 261740 263692 261752
rect 263744 261740 263750 261792
rect 164234 261672 164240 261724
rect 164292 261712 164298 261724
rect 263594 261712 263600 261724
rect 164292 261684 263600 261712
rect 164292 261672 164298 261684
rect 263594 261672 263600 261684
rect 263652 261672 263658 261724
rect 325694 261672 325700 261724
rect 325752 261712 325758 261724
rect 487154 261712 487160 261724
rect 325752 261684 487160 261712
rect 325752 261672 325758 261684
rect 487154 261672 487160 261684
rect 487212 261672 487218 261724
rect 160186 261604 160192 261656
rect 160244 261644 160250 261656
rect 260098 261644 260104 261656
rect 160244 261616 260104 261644
rect 160244 261604 160250 261616
rect 260098 261604 260104 261616
rect 260156 261604 260162 261656
rect 327166 261604 327172 261656
rect 327224 261644 327230 261656
rect 490006 261644 490012 261656
rect 327224 261616 490012 261644
rect 327224 261604 327230 261616
rect 490006 261604 490012 261616
rect 490064 261604 490070 261656
rect 128354 261536 128360 261588
rect 128412 261576 128418 261588
rect 256970 261576 256976 261588
rect 128412 261548 256976 261576
rect 128412 261536 128418 261548
rect 256970 261536 256976 261548
rect 257028 261536 257034 261588
rect 327074 261536 327080 261588
rect 327132 261576 327138 261588
rect 494054 261576 494060 261588
rect 327132 261548 494060 261576
rect 327132 261536 327138 261548
rect 494054 261536 494060 261548
rect 494112 261536 494118 261588
rect 82814 261468 82820 261520
rect 82872 261508 82878 261520
rect 248598 261508 248604 261520
rect 82872 261480 248604 261508
rect 82872 261468 82878 261480
rect 248598 261468 248604 261480
rect 248656 261468 248662 261520
rect 336918 261468 336924 261520
rect 336976 261508 336982 261520
rect 539686 261508 539692 261520
rect 336976 261480 539692 261508
rect 336976 261468 336982 261480
rect 539686 261468 539692 261480
rect 539744 261468 539750 261520
rect 211798 260312 211804 260364
rect 211856 260352 211862 260364
rect 266814 260352 266820 260364
rect 211856 260324 266820 260352
rect 211856 260312 211862 260324
rect 266814 260312 266820 260324
rect 266872 260312 266878 260364
rect 125594 260244 125600 260296
rect 125652 260284 125658 260296
rect 256878 260284 256884 260296
rect 125652 260256 256884 260284
rect 125652 260244 125658 260256
rect 256878 260244 256884 260256
rect 256936 260244 256942 260296
rect 324590 260244 324596 260296
rect 324648 260284 324654 260296
rect 480254 260284 480260 260296
rect 324648 260256 480260 260284
rect 324648 260244 324654 260256
rect 480254 260244 480260 260256
rect 480312 260244 480318 260296
rect 64874 260176 64880 260228
rect 64932 260216 64938 260228
rect 244366 260216 244372 260228
rect 64932 260188 244372 260216
rect 64932 260176 64938 260188
rect 244366 260176 244372 260188
rect 244424 260176 244430 260228
rect 333974 260176 333980 260228
rect 334032 260216 334038 260228
rect 525794 260216 525800 260228
rect 334032 260188 525800 260216
rect 334032 260176 334038 260188
rect 525794 260176 525800 260188
rect 525852 260176 525858 260228
rect 35894 260108 35900 260160
rect 35952 260148 35958 260160
rect 238938 260148 238944 260160
rect 35952 260120 238944 260148
rect 35952 260108 35958 260120
rect 238938 260108 238944 260120
rect 238996 260108 239002 260160
rect 343818 260108 343824 260160
rect 343876 260148 343882 260160
rect 575474 260148 575480 260160
rect 343876 260120 575480 260148
rect 343876 260108 343882 260120
rect 575474 260108 575480 260120
rect 575532 260108 575538 260160
rect 217226 258952 217232 259004
rect 217284 258992 217290 259004
rect 344094 258992 344100 259004
rect 217284 258964 344100 258992
rect 217284 258952 217290 258964
rect 344094 258952 344100 258964
rect 344152 258952 344158 259004
rect 69106 258884 69112 258936
rect 69164 258924 69170 258936
rect 245746 258924 245752 258936
rect 69164 258896 245752 258924
rect 69164 258884 69170 258896
rect 245746 258884 245752 258896
rect 245804 258884 245810 258936
rect 60734 258816 60740 258868
rect 60792 258856 60798 258868
rect 244734 258856 244740 258868
rect 60792 258828 244740 258856
rect 60792 258816 60798 258828
rect 244734 258816 244740 258828
rect 244792 258816 244798 258868
rect 35250 258748 35256 258800
rect 35308 258788 35314 258800
rect 238846 258788 238852 258800
rect 35308 258760 238852 258788
rect 35308 258748 35314 258760
rect 238846 258748 238852 258760
rect 238904 258748 238910 258800
rect 4798 258680 4804 258732
rect 4856 258720 4862 258732
rect 231854 258720 231860 258732
rect 4856 258692 231860 258720
rect 4856 258680 4862 258692
rect 231854 258680 231860 258692
rect 231912 258680 231918 258732
rect 320266 256164 320272 256216
rect 320324 256204 320330 256216
rect 454034 256204 454040 256216
rect 320324 256176 454040 256204
rect 320324 256164 320330 256176
rect 454034 256164 454040 256176
rect 454092 256164 454098 256216
rect 24854 256096 24860 256148
rect 24912 256136 24918 256148
rect 236086 256136 236092 256148
rect 24912 256108 236092 256136
rect 24912 256096 24918 256108
rect 236086 256096 236092 256108
rect 236144 256096 236150 256148
rect 321646 256096 321652 256148
rect 321704 256136 321710 256148
rect 460934 256136 460940 256148
rect 321704 256108 460940 256136
rect 321704 256096 321710 256108
rect 460934 256096 460940 256108
rect 460992 256096 460998 256148
rect 17218 256028 17224 256080
rect 17276 256068 17282 256080
rect 234982 256068 234988 256080
rect 17276 256040 234988 256068
rect 17276 256028 17282 256040
rect 234982 256028 234988 256040
rect 235040 256028 235046 256080
rect 323026 256028 323032 256080
rect 323084 256068 323090 256080
rect 467834 256068 467840 256080
rect 323084 256040 467840 256068
rect 323084 256028 323090 256040
rect 467834 256028 467840 256040
rect 467892 256028 467898 256080
rect 8938 255960 8944 256012
rect 8996 256000 9002 256012
rect 233418 256000 233424 256012
rect 8996 255972 233424 256000
rect 8996 255960 9002 255972
rect 233418 255960 233424 255972
rect 233476 255960 233482 256012
rect 324498 255960 324504 256012
rect 324556 256000 324562 256012
rect 474734 256000 474740 256012
rect 324556 255972 474740 256000
rect 324556 255960 324562 255972
rect 474734 255960 474740 255972
rect 474792 255960 474798 256012
rect 116578 254804 116584 254856
rect 116636 254844 116642 254856
rect 240226 254844 240232 254856
rect 116636 254816 240232 254844
rect 116636 254804 116642 254816
rect 240226 254804 240232 254816
rect 240284 254804 240290 254856
rect 79318 254736 79324 254788
rect 79376 254776 79382 254788
rect 243078 254776 243084 254788
rect 79376 254748 243084 254776
rect 79376 254736 79382 254748
rect 243078 254736 243084 254748
rect 243136 254736 243142 254788
rect 56594 254668 56600 254720
rect 56652 254708 56658 254720
rect 243170 254708 243176 254720
rect 56652 254680 243176 254708
rect 56652 254668 56658 254680
rect 243170 254668 243176 254680
rect 243228 254668 243234 254720
rect 318058 254668 318064 254720
rect 318116 254708 318122 254720
rect 432046 254708 432052 254720
rect 318116 254680 432052 254708
rect 318116 254668 318122 254680
rect 432046 254668 432052 254680
rect 432104 254668 432110 254720
rect 44266 254600 44272 254652
rect 44324 254640 44330 254652
rect 240594 254640 240600 254652
rect 44324 254612 240600 254640
rect 44324 254600 44330 254612
rect 240594 254600 240600 254612
rect 240652 254600 240658 254652
rect 342346 254600 342352 254652
rect 342404 254640 342410 254652
rect 574094 254640 574100 254652
rect 342404 254612 574100 254640
rect 342404 254600 342410 254612
rect 574094 254600 574100 254612
rect 574152 254600 574158 254652
rect 39298 254532 39304 254584
rect 39356 254572 39362 254584
rect 239214 254572 239220 254584
rect 39356 254544 239220 254572
rect 39356 254532 39362 254544
rect 239214 254532 239220 254544
rect 239272 254532 239278 254584
rect 344002 254532 344008 254584
rect 344060 254572 344066 254584
rect 578234 254572 578240 254584
rect 344060 254544 578240 254572
rect 344060 254532 344066 254544
rect 578234 254532 578240 254544
rect 578292 254532 578298 254584
rect 2866 254192 2872 254244
rect 2924 254232 2930 254244
rect 4890 254232 4896 254244
rect 2924 254204 4896 254232
rect 2924 254192 2930 254204
rect 4890 254192 4896 254204
rect 4948 254192 4954 254244
rect 86954 253444 86960 253496
rect 87012 253484 87018 253496
rect 248874 253484 248880 253496
rect 87012 253456 248880 253484
rect 87012 253444 87018 253456
rect 248874 253444 248880 253456
rect 248932 253444 248938 253496
rect 294230 253444 294236 253496
rect 294288 253484 294294 253496
rect 365990 253484 365996 253496
rect 294288 253456 365996 253484
rect 294288 253444 294294 253456
rect 365990 253444 365996 253456
rect 366048 253444 366054 253496
rect 84194 253376 84200 253428
rect 84252 253416 84258 253428
rect 248506 253416 248512 253428
rect 84252 253388 248512 253416
rect 84252 253376 84258 253388
rect 248506 253376 248512 253388
rect 248564 253376 248570 253428
rect 331214 253376 331220 253428
rect 331272 253416 331278 253428
rect 514846 253416 514852 253428
rect 331272 253388 514852 253416
rect 331272 253376 331278 253388
rect 514846 253376 514852 253388
rect 514904 253376 514910 253428
rect 80054 253308 80060 253360
rect 80112 253348 80118 253360
rect 247218 253348 247224 253360
rect 80112 253320 247224 253348
rect 80112 253308 80118 253320
rect 247218 253308 247224 253320
rect 247276 253308 247282 253360
rect 332686 253308 332692 253360
rect 332744 253348 332750 253360
rect 517514 253348 517520 253360
rect 332744 253320 517520 253348
rect 332744 253308 332750 253320
rect 517514 253308 517520 253320
rect 517572 253308 517578 253360
rect 17954 253240 17960 253292
rect 18012 253280 18018 253292
rect 234890 253280 234896 253292
rect 18012 253252 234896 253280
rect 18012 253240 18018 253252
rect 234890 253240 234896 253252
rect 234948 253240 234954 253292
rect 332778 253240 332784 253292
rect 332836 253280 332842 253292
rect 521654 253280 521660 253292
rect 332836 253252 521660 253280
rect 332836 253240 332842 253252
rect 521654 253240 521660 253252
rect 521712 253240 521718 253292
rect 9674 253172 9680 253224
rect 9732 253212 9738 253224
rect 233326 253212 233332 253224
rect 9732 253184 233332 253212
rect 9732 253172 9738 253184
rect 233326 253172 233332 253184
rect 233384 253172 233390 253224
rect 342254 253172 342260 253224
rect 342312 253212 342318 253224
rect 571334 253212 571340 253224
rect 342312 253184 571340 253212
rect 342312 253172 342318 253184
rect 571334 253172 571340 253184
rect 571392 253172 571398 253224
rect 218514 252152 218520 252204
rect 218572 252192 218578 252204
rect 347774 252192 347780 252204
rect 218572 252164 347780 252192
rect 218572 252152 218578 252164
rect 347774 252152 347780 252164
rect 347832 252152 347838 252204
rect 121454 252084 121460 252136
rect 121512 252124 121518 252136
rect 255774 252124 255780 252136
rect 121512 252096 255780 252124
rect 121512 252084 121518 252096
rect 255774 252084 255780 252096
rect 255832 252084 255838 252136
rect 31018 252016 31024 252068
rect 31076 252056 31082 252068
rect 237834 252056 237840 252068
rect 31076 252028 237840 252056
rect 31076 252016 31082 252028
rect 237834 252016 237840 252028
rect 237892 252016 237898 252068
rect 317506 252016 317512 252068
rect 317564 252056 317570 252068
rect 445754 252056 445760 252068
rect 317564 252028 445760 252056
rect 317564 252016 317570 252028
rect 445754 252016 445760 252028
rect 445812 252016 445818 252068
rect 26234 251948 26240 252000
rect 26292 251988 26298 252000
rect 237466 251988 237472 252000
rect 26292 251960 237472 251988
rect 26292 251948 26298 251960
rect 237466 251948 237472 251960
rect 237524 251948 237530 252000
rect 318794 251948 318800 252000
rect 318852 251988 318858 252000
rect 448606 251988 448612 252000
rect 318852 251960 448612 251988
rect 318852 251948 318858 251960
rect 448606 251948 448612 251960
rect 448664 251948 448670 252000
rect 20714 251880 20720 251932
rect 20772 251920 20778 251932
rect 236362 251920 236368 251932
rect 20772 251892 236368 251920
rect 20772 251880 20778 251892
rect 236362 251880 236368 251892
rect 236420 251880 236426 251932
rect 318886 251880 318892 251932
rect 318944 251920 318950 251932
rect 452654 251920 452660 251932
rect 318944 251892 452660 251920
rect 318944 251880 318950 251892
rect 452654 251880 452660 251892
rect 452712 251880 452718 251932
rect 12434 251812 12440 251864
rect 12492 251852 12498 251864
rect 234798 251852 234804 251864
rect 12492 251824 234804 251852
rect 12492 251812 12498 251824
rect 234798 251812 234804 251824
rect 234856 251812 234862 251864
rect 320174 251812 320180 251864
rect 320232 251852 320238 251864
rect 456886 251852 456892 251864
rect 320232 251824 456892 251852
rect 320232 251812 320238 251824
rect 456886 251812 456892 251824
rect 456944 251812 456950 251864
rect 292850 251132 292856 251184
rect 292908 251172 292914 251184
rect 358814 251172 358820 251184
rect 292908 251144 358820 251172
rect 292908 251132 292914 251144
rect 358814 251132 358820 251144
rect 358872 251132 358878 251184
rect 298370 251064 298376 251116
rect 298428 251104 298434 251116
rect 364702 251104 364708 251116
rect 298428 251076 364708 251104
rect 298428 251064 298434 251076
rect 364702 251064 364708 251076
rect 364760 251064 364766 251116
rect 299934 250996 299940 251048
rect 299992 251036 299998 251048
rect 367186 251036 367192 251048
rect 299992 251008 367192 251036
rect 299992 250996 299998 251008
rect 367186 250996 367192 251008
rect 367244 250996 367250 251048
rect 292942 250928 292948 250980
rect 293000 250968 293006 250980
rect 360194 250968 360200 250980
rect 293000 250940 360200 250968
rect 293000 250928 293006 250940
rect 360194 250928 360200 250940
rect 360252 250928 360258 250980
rect 295794 250860 295800 250912
rect 295852 250900 295858 250912
rect 363138 250900 363144 250912
rect 295852 250872 363144 250900
rect 295852 250860 295858 250872
rect 363138 250860 363144 250872
rect 363196 250860 363202 250912
rect 297174 250792 297180 250844
rect 297232 250832 297238 250844
rect 364794 250832 364800 250844
rect 297232 250804 364800 250832
rect 297232 250792 297238 250804
rect 364794 250792 364800 250804
rect 364852 250792 364858 250844
rect 174538 250724 174544 250776
rect 174596 250764 174602 250776
rect 251634 250764 251640 250776
rect 174596 250736 251640 250764
rect 174596 250724 174602 250736
rect 251634 250724 251640 250736
rect 251692 250724 251698 250776
rect 298462 250724 298468 250776
rect 298520 250764 298526 250776
rect 367094 250764 367100 250776
rect 298520 250736 367100 250764
rect 298520 250724 298526 250736
rect 367094 250724 367100 250736
rect 367152 250724 367158 250776
rect 78674 250656 78680 250708
rect 78732 250696 78738 250708
rect 247126 250696 247132 250708
rect 78732 250668 247132 250696
rect 78732 250656 78738 250668
rect 247126 250656 247132 250668
rect 247184 250656 247190 250708
rect 293034 250656 293040 250708
rect 293092 250696 293098 250708
rect 364886 250696 364892 250708
rect 293092 250668 364892 250696
rect 293092 250656 293098 250668
rect 364886 250656 364892 250668
rect 364944 250656 364950 250708
rect 75914 250588 75920 250640
rect 75972 250628 75978 250640
rect 247034 250628 247040 250640
rect 75972 250600 247040 250628
rect 75972 250588 75978 250600
rect 247034 250588 247040 250600
rect 247092 250588 247098 250640
rect 291470 250588 291476 250640
rect 291528 250628 291534 250640
rect 368474 250628 368480 250640
rect 291528 250600 368480 250628
rect 291528 250588 291534 250600
rect 368474 250588 368480 250600
rect 368532 250588 368538 250640
rect 71774 250520 71780 250572
rect 71832 250560 71838 250572
rect 245654 250560 245660 250572
rect 71832 250532 245660 250560
rect 71832 250520 71838 250532
rect 245654 250520 245660 250532
rect 245712 250520 245718 250572
rect 304994 250520 305000 250572
rect 305052 250560 305058 250572
rect 382366 250560 382372 250572
rect 305052 250532 382372 250560
rect 305052 250520 305058 250532
rect 382366 250520 382372 250532
rect 382424 250520 382430 250572
rect 16574 250452 16580 250504
rect 16632 250492 16638 250504
rect 234706 250492 234712 250504
rect 16632 250464 234712 250492
rect 16632 250452 16638 250464
rect 234706 250452 234712 250464
rect 234764 250452 234770 250504
rect 291562 250452 291568 250504
rect 291620 250492 291626 250504
rect 369854 250492 369860 250504
rect 291620 250464 369860 250492
rect 291620 250452 291626 250464
rect 369854 250452 369860 250464
rect 369912 250452 369918 250504
rect 297266 250384 297272 250436
rect 297324 250424 297330 250436
rect 363230 250424 363236 250436
rect 297324 250396 363236 250424
rect 297324 250384 297330 250396
rect 363230 250384 363236 250396
rect 363288 250384 363294 250436
rect 301222 250316 301228 250368
rect 301280 250356 301286 250368
rect 365898 250356 365904 250368
rect 301280 250328 365904 250356
rect 301280 250316 301286 250328
rect 365898 250316 365904 250328
rect 365956 250316 365962 250368
rect 295702 250248 295708 250300
rect 295760 250288 295766 250300
rect 360286 250288 360292 250300
rect 295760 250260 360292 250288
rect 295760 250248 295766 250260
rect 360286 250248 360292 250260
rect 360344 250248 360350 250300
rect 209866 249228 209872 249280
rect 209924 249268 209930 249280
rect 272334 249268 272340 249280
rect 209924 249240 272340 249268
rect 209924 249228 209930 249240
rect 272334 249228 272340 249240
rect 272392 249228 272398 249280
rect 317414 249228 317420 249280
rect 317472 249268 317478 249280
rect 441614 249268 441620 249280
rect 317472 249240 441620 249268
rect 317472 249228 317478 249240
rect 441614 249228 441620 249240
rect 441672 249228 441678 249280
rect 201586 249160 201592 249212
rect 201644 249200 201650 249212
rect 270494 249200 270500 249212
rect 201644 249172 270500 249200
rect 201644 249160 201650 249172
rect 270494 249160 270500 249172
rect 270552 249160 270558 249212
rect 336734 249160 336740 249212
rect 336792 249200 336798 249212
rect 534718 249200 534724 249212
rect 336792 249172 534724 249200
rect 336792 249160 336798 249172
rect 534718 249160 534724 249172
rect 534776 249160 534782 249212
rect 135254 249092 135260 249144
rect 135312 249132 135318 249144
rect 258442 249132 258448 249144
rect 135312 249104 258448 249132
rect 135312 249092 135318 249104
rect 258442 249092 258448 249104
rect 258500 249092 258506 249144
rect 335446 249092 335452 249144
rect 335504 249132 335510 249144
rect 534074 249132 534080 249144
rect 335504 249104 534080 249132
rect 335504 249092 335510 249104
rect 534074 249092 534080 249104
rect 534132 249092 534138 249144
rect 57974 249024 57980 249076
rect 58032 249064 58038 249076
rect 242986 249064 242992 249076
rect 58032 249036 242992 249064
rect 58032 249024 58038 249036
rect 242986 249024 242992 249036
rect 243044 249024 243050 249076
rect 335354 249024 335360 249076
rect 335412 249064 335418 249076
rect 538214 249064 538220 249076
rect 335412 249036 538220 249064
rect 335412 249024 335418 249036
rect 538214 249024 538220 249036
rect 538272 249024 538278 249076
rect 299750 248344 299756 248396
rect 299808 248384 299814 248396
rect 363322 248384 363328 248396
rect 299808 248356 363328 248384
rect 299808 248344 299814 248356
rect 363322 248344 363328 248356
rect 363380 248344 363386 248396
rect 298278 248276 298284 248328
rect 298336 248316 298342 248328
rect 362954 248316 362960 248328
rect 298336 248288 362960 248316
rect 298336 248276 298342 248288
rect 362954 248276 362960 248288
rect 363012 248276 363018 248328
rect 295610 248208 295616 248260
rect 295668 248248 295674 248260
rect 361666 248248 361672 248260
rect 295668 248220 361672 248248
rect 295668 248208 295674 248220
rect 361666 248208 361672 248220
rect 361724 248208 361730 248260
rect 298186 248140 298192 248192
rect 298244 248180 298250 248192
rect 364610 248180 364616 248192
rect 298244 248152 364616 248180
rect 298244 248140 298250 248152
rect 364610 248140 364616 248152
rect 364668 248140 364674 248192
rect 296990 248072 296996 248124
rect 297048 248112 297054 248124
rect 364334 248112 364340 248124
rect 297048 248084 364340 248112
rect 297048 248072 297054 248084
rect 364334 248072 364340 248084
rect 364392 248072 364398 248124
rect 297082 248004 297088 248056
rect 297140 248044 297146 248056
rect 364518 248044 364524 248056
rect 297140 248016 364524 248044
rect 297140 248004 297146 248016
rect 364518 248004 364524 248016
rect 364576 248004 364582 248056
rect 151906 247936 151912 247988
rect 151964 247976 151970 247988
rect 260834 247976 260840 247988
rect 151964 247948 260840 247976
rect 151964 247936 151970 247948
rect 260834 247936 260840 247948
rect 260892 247936 260898 247988
rect 296806 247936 296812 247988
rect 296864 247976 296870 247988
rect 364426 247976 364432 247988
rect 296864 247948 364432 247976
rect 296864 247936 296870 247948
rect 364426 247936 364432 247948
rect 364484 247936 364490 247988
rect 147674 247868 147680 247920
rect 147732 247908 147738 247920
rect 260926 247908 260932 247920
rect 147732 247880 260932 247908
rect 147732 247868 147738 247880
rect 260926 247868 260932 247880
rect 260984 247868 260990 247920
rect 292666 247868 292672 247920
rect 292724 247908 292730 247920
rect 360838 247908 360844 247920
rect 292724 247880 360844 247908
rect 292724 247868 292730 247880
rect 360838 247868 360844 247880
rect 360896 247868 360902 247920
rect 143534 247800 143540 247852
rect 143592 247840 143598 247852
rect 259546 247840 259552 247852
rect 143592 247812 259552 247840
rect 143592 247800 143598 247812
rect 259546 247800 259552 247812
rect 259604 247800 259610 247852
rect 292758 247800 292764 247852
rect 292816 247840 292822 247852
rect 362126 247840 362132 247852
rect 292816 247812 362132 247840
rect 292816 247800 292822 247812
rect 362126 247800 362132 247812
rect 362184 247800 362190 247852
rect 127066 247732 127072 247784
rect 127124 247772 127130 247784
rect 256786 247772 256792 247784
rect 127124 247744 256792 247772
rect 127124 247732 127130 247744
rect 256786 247732 256792 247744
rect 256844 247732 256850 247784
rect 291378 247732 291384 247784
rect 291436 247772 291442 247784
rect 366082 247772 366088 247784
rect 291436 247744 366088 247772
rect 291436 247732 291442 247744
rect 366082 247732 366088 247744
rect 366140 247732 366146 247784
rect 53834 247664 53840 247716
rect 53892 247704 53898 247716
rect 242894 247704 242900 247716
rect 53892 247676 242900 247704
rect 53892 247664 53898 247676
rect 242894 247664 242900 247676
rect 242952 247664 242958 247716
rect 288710 247664 288716 247716
rect 288768 247704 288774 247716
rect 364978 247704 364984 247716
rect 288768 247676 364984 247704
rect 288768 247664 288774 247676
rect 364978 247664 364984 247676
rect 365036 247664 365042 247716
rect 294138 247596 294144 247648
rect 294196 247636 294202 247648
rect 356698 247636 356704 247648
rect 294196 247608 356704 247636
rect 294196 247596 294202 247608
rect 356698 247596 356704 247608
rect 356756 247596 356762 247648
rect 295426 247528 295432 247580
rect 295484 247568 295490 247580
rect 358354 247568 358360 247580
rect 295484 247540 358360 247568
rect 295484 247528 295490 247540
rect 358354 247528 358360 247540
rect 358412 247528 358418 247580
rect 301130 247460 301136 247512
rect 301188 247500 301194 247512
rect 363046 247500 363052 247512
rect 301188 247472 363052 247500
rect 301188 247460 301194 247472
rect 363046 247460 363052 247472
rect 363104 247460 363110 247512
rect 211154 246576 211160 246628
rect 211212 246616 211218 246628
rect 273254 246616 273260 246628
rect 211212 246588 273260 246616
rect 211212 246576 211218 246588
rect 273254 246576 273260 246588
rect 273312 246576 273318 246628
rect 314746 246576 314752 246628
rect 314804 246616 314810 246628
rect 387058 246616 387064 246628
rect 314804 246588 387064 246616
rect 314804 246576 314810 246588
rect 387058 246576 387064 246588
rect 387116 246576 387122 246628
rect 53098 246508 53104 246560
rect 53156 246548 53162 246560
rect 241514 246548 241520 246560
rect 53156 246520 241520 246548
rect 53156 246508 53162 246520
rect 241514 246508 241520 246520
rect 241572 246508 241578 246560
rect 289998 246508 290004 246560
rect 290056 246548 290062 246560
rect 367278 246548 367284 246560
rect 290056 246520 367284 246548
rect 290056 246508 290062 246520
rect 367278 246508 367284 246520
rect 367336 246508 367342 246560
rect 48958 246440 48964 246492
rect 49016 246480 49022 246492
rect 241606 246480 241612 246492
rect 49016 246452 241612 246480
rect 49016 246440 49022 246452
rect 241606 246440 241612 246452
rect 241664 246440 241670 246492
rect 310514 246440 310520 246492
rect 310572 246480 310578 246492
rect 405734 246480 405740 246492
rect 310572 246452 405740 246480
rect 310572 246440 310578 246452
rect 405734 246440 405740 246452
rect 405792 246440 405798 246492
rect 13078 246372 13084 246424
rect 13136 246412 13142 246424
rect 234614 246412 234620 246424
rect 13136 246384 234620 246412
rect 13136 246372 13142 246384
rect 234614 246372 234620 246384
rect 234672 246372 234678 246424
rect 314654 246372 314660 246424
rect 314712 246412 314718 246424
rect 430574 246412 430580 246424
rect 314712 246384 430580 246412
rect 314712 246372 314718 246384
rect 430574 246372 430580 246384
rect 430632 246372 430638 246424
rect 6914 246304 6920 246356
rect 6972 246344 6978 246356
rect 233694 246344 233700 246356
rect 6972 246316 233700 246344
rect 6972 246304 6978 246316
rect 233694 246304 233700 246316
rect 233752 246304 233758 246356
rect 324406 246304 324412 246356
rect 324464 246344 324470 246356
rect 481726 246344 481732 246356
rect 324464 246316 481732 246344
rect 324464 246304 324470 246316
rect 481726 246304 481732 246316
rect 481784 246304 481790 246356
rect 300854 245556 300860 245608
rect 300912 245596 300918 245608
rect 357434 245596 357440 245608
rect 300912 245568 357440 245596
rect 300912 245556 300918 245568
rect 357434 245556 357440 245568
rect 357492 245556 357498 245608
rect 300946 245488 300952 245540
rect 301004 245528 301010 245540
rect 358170 245528 358176 245540
rect 301004 245500 358176 245528
rect 301004 245488 301010 245500
rect 358170 245488 358176 245500
rect 358228 245488 358234 245540
rect 355778 245420 355784 245472
rect 355836 245460 355842 245472
rect 368566 245460 368572 245472
rect 355836 245432 368572 245460
rect 355836 245420 355842 245432
rect 368566 245420 368572 245432
rect 368624 245420 368630 245472
rect 219250 245352 219256 245404
rect 219308 245392 219314 245404
rect 287422 245392 287428 245404
rect 219308 245364 287428 245392
rect 219308 245352 219314 245364
rect 287422 245352 287428 245364
rect 287480 245352 287486 245404
rect 294046 245352 294052 245404
rect 294104 245392 294110 245404
rect 358078 245392 358084 245404
rect 294104 245364 358084 245392
rect 294104 245352 294110 245364
rect 358078 245352 358084 245364
rect 358136 245352 358142 245404
rect 213638 245284 213644 245336
rect 213696 245324 213702 245336
rect 288526 245324 288532 245336
rect 213696 245296 288532 245324
rect 213696 245284 213702 245296
rect 288526 245284 288532 245296
rect 288584 245284 288590 245336
rect 293954 245284 293960 245336
rect 294012 245324 294018 245336
rect 358170 245324 358176 245336
rect 294012 245296 358176 245324
rect 294012 245284 294018 245296
rect 358170 245284 358176 245296
rect 358228 245284 358234 245336
rect 358262 245284 358268 245336
rect 358320 245324 358326 245336
rect 367370 245324 367376 245336
rect 358320 245296 367376 245324
rect 358320 245284 358326 245296
rect 367370 245284 367376 245296
rect 367428 245284 367434 245336
rect 212994 245216 213000 245268
rect 213052 245256 213058 245268
rect 288618 245256 288624 245268
rect 213052 245228 288624 245256
rect 213052 245216 213058 245228
rect 288618 245216 288624 245228
rect 288676 245216 288682 245268
rect 292574 245216 292580 245268
rect 292632 245256 292638 245268
rect 359458 245256 359464 245268
rect 292632 245228 359464 245256
rect 292632 245216 292638 245228
rect 359458 245216 359464 245228
rect 359516 245216 359522 245268
rect 143626 245148 143632 245200
rect 143684 245188 143690 245200
rect 259454 245188 259460 245200
rect 143684 245160 259460 245188
rect 143684 245148 143690 245160
rect 259454 245148 259460 245160
rect 259512 245148 259518 245200
rect 291286 245148 291292 245200
rect 291344 245188 291350 245200
rect 368658 245188 368664 245200
rect 291344 245160 368664 245188
rect 291344 245148 291350 245160
rect 368658 245148 368664 245160
rect 368716 245148 368722 245200
rect 135346 245080 135352 245132
rect 135404 245120 135410 245132
rect 254578 245120 254584 245132
rect 135404 245092 254584 245120
rect 135404 245080 135410 245092
rect 254578 245080 254584 245092
rect 254636 245080 254642 245132
rect 324314 245080 324320 245132
rect 324372 245120 324378 245132
rect 476114 245120 476120 245132
rect 324372 245092 476120 245120
rect 324372 245080 324378 245092
rect 476114 245080 476120 245092
rect 476172 245080 476178 245132
rect 129734 245012 129740 245064
rect 129792 245052 129798 245064
rect 256694 245052 256700 245064
rect 129792 245024 256700 245052
rect 129792 245012 129798 245024
rect 256694 245012 256700 245024
rect 256752 245012 256758 245064
rect 339494 245012 339500 245064
rect 339552 245052 339558 245064
rect 557534 245052 557540 245064
rect 339552 245024 557540 245052
rect 339552 245012 339558 245024
rect 557534 245012 557540 245024
rect 557592 245012 557598 245064
rect 7650 244944 7656 244996
rect 7708 244984 7714 244996
rect 231946 244984 231952 244996
rect 7708 244956 231952 244984
rect 7708 244944 7714 244956
rect 231946 244944 231952 244956
rect 232004 244944 232010 244996
rect 340874 244944 340880 244996
rect 340932 244984 340938 244996
rect 561674 244984 561680 244996
rect 340932 244956 561680 244984
rect 340932 244944 340938 244956
rect 561674 244944 561680 244956
rect 561732 244944 561738 244996
rect 4890 244876 4896 244928
rect 4948 244916 4954 244928
rect 232038 244916 232044 244928
rect 4948 244888 232044 244916
rect 4948 244876 4954 244888
rect 232038 244876 232044 244888
rect 232096 244876 232102 244928
rect 340966 244876 340972 244928
rect 341024 244916 341030 244928
rect 564526 244916 564532 244928
rect 341024 244888 564532 244916
rect 341024 244876 341030 244888
rect 564526 244876 564532 244888
rect 564584 244876 564590 244928
rect 355594 244536 355600 244588
rect 355652 244576 355658 244588
rect 363506 244576 363512 244588
rect 355652 244548 363512 244576
rect 355652 244536 355658 244548
rect 363506 244536 363512 244548
rect 363564 244536 363570 244588
rect 355686 244264 355692 244316
rect 355744 244304 355750 244316
rect 362310 244304 362316 244316
rect 355744 244276 362316 244304
rect 355744 244264 355750 244276
rect 362310 244264 362316 244276
rect 362368 244264 362374 244316
rect 355318 244128 355324 244180
rect 355376 244168 355382 244180
rect 362218 244168 362224 244180
rect 355376 244140 362224 244168
rect 355376 244128 355382 244140
rect 362218 244128 362224 244140
rect 362276 244128 362282 244180
rect 355410 243788 355416 243840
rect 355468 243828 355474 243840
rect 369946 243828 369952 243840
rect 355468 243800 369952 243828
rect 355468 243788 355474 243800
rect 369946 243788 369952 243800
rect 370004 243788 370010 243840
rect 291194 243720 291200 243772
rect 291252 243760 291258 243772
rect 358262 243760 358268 243772
rect 291252 243732 358268 243760
rect 291252 243720 291258 243732
rect 358262 243720 358268 243732
rect 358320 243720 358326 243772
rect 219158 243652 219164 243704
rect 219216 243692 219222 243704
rect 286042 243692 286048 243704
rect 219216 243664 286048 243692
rect 219216 243652 219222 243664
rect 286042 243652 286048 243664
rect 286100 243652 286106 243704
rect 289906 243652 289912 243704
rect 289964 243692 289970 243704
rect 359550 243692 359556 243704
rect 289964 243664 359556 243692
rect 289964 243652 289970 243664
rect 359550 243652 359556 243664
rect 359608 243652 359614 243704
rect 218606 243584 218612 243636
rect 218664 243624 218670 243636
rect 285766 243624 285772 243636
rect 218664 243596 285772 243624
rect 218664 243584 218670 243596
rect 285766 243584 285772 243596
rect 285824 243584 285830 243636
rect 289814 243584 289820 243636
rect 289872 243624 289878 243636
rect 360930 243624 360936 243636
rect 289872 243596 360936 243624
rect 289872 243584 289878 243596
rect 360930 243584 360936 243596
rect 360988 243584 360994 243636
rect 217134 243516 217140 243568
rect 217192 243556 217198 243568
rect 287330 243556 287336 243568
rect 217192 243528 287336 243556
rect 217192 243516 217198 243528
rect 287330 243516 287336 243528
rect 287388 243516 287394 243568
rect 288434 243516 288440 243568
rect 288492 243556 288498 243568
rect 363598 243556 363604 243568
rect 288492 243528 363604 243556
rect 288492 243516 288498 243528
rect 363598 243516 363604 243528
rect 363656 243516 363662 243568
rect 215754 195780 215760 195832
rect 215812 195820 215818 195832
rect 217502 195820 217508 195832
rect 215812 195792 217508 195820
rect 215812 195780 215818 195792
rect 217502 195780 217508 195792
rect 217560 195780 217566 195832
rect 214374 195236 214380 195288
rect 214432 195276 214438 195288
rect 217318 195276 217324 195288
rect 214432 195248 217324 195276
rect 214432 195236 214438 195248
rect 217318 195236 217324 195248
rect 217376 195236 217382 195288
rect 210694 193128 210700 193180
rect 210752 193168 210758 193180
rect 216674 193168 216680 193180
rect 210752 193140 216680 193168
rect 210752 193128 210758 193140
rect 216674 193128 216680 193140
rect 216732 193128 216738 193180
rect 210878 189660 210884 189712
rect 210936 189700 210942 189712
rect 218054 189700 218060 189712
rect 210936 189672 218060 189700
rect 210936 189660 210942 189672
rect 218054 189660 218060 189672
rect 218112 189660 218118 189712
rect 210786 188980 210792 189032
rect 210844 189020 210850 189032
rect 216674 189020 216680 189032
rect 210844 188992 216680 189020
rect 210844 188980 210850 188992
rect 216674 188980 216680 188992
rect 216732 188980 216738 189032
rect 212994 168920 213000 168972
rect 213052 168960 213058 168972
rect 217410 168960 217416 168972
rect 213052 168932 217416 168960
rect 213052 168920 213058 168932
rect 217410 168920 217416 168932
rect 217468 168920 217474 168972
rect 218790 166268 218796 166320
rect 218848 166308 218854 166320
rect 218974 166308 218980 166320
rect 218848 166280 218980 166308
rect 218848 166268 218854 166280
rect 218974 166268 218980 166280
rect 219032 166268 219038 166320
rect 356238 159808 356244 159860
rect 356296 159848 356302 159860
rect 357986 159848 357992 159860
rect 356296 159820 357992 159848
rect 356296 159808 356302 159820
rect 357986 159808 357992 159820
rect 358044 159808 358050 159860
rect 214466 159604 214472 159656
rect 214524 159644 214530 159656
rect 256694 159644 256700 159656
rect 214524 159616 256700 159644
rect 214524 159604 214530 159616
rect 256694 159604 256700 159616
rect 256752 159604 256758 159656
rect 211706 159536 211712 159588
rect 211764 159576 211770 159588
rect 255314 159576 255320 159588
rect 211764 159548 255320 159576
rect 211764 159536 211770 159548
rect 255314 159536 255320 159548
rect 255372 159536 255378 159588
rect 317690 159536 317696 159588
rect 317748 159576 317754 159588
rect 356790 159576 356796 159588
rect 317748 159548 356796 159576
rect 317748 159536 317754 159548
rect 356790 159536 356796 159548
rect 356848 159536 356854 159588
rect 213178 159468 213184 159520
rect 213236 159508 213242 159520
rect 259546 159508 259552 159520
rect 213236 159480 259552 159508
rect 213236 159468 213242 159480
rect 259546 159468 259552 159480
rect 259604 159468 259610 159520
rect 314654 159468 314660 159520
rect 314712 159508 314718 159520
rect 357802 159508 357808 159520
rect 314712 159480 357808 159508
rect 314712 159468 314718 159480
rect 357802 159468 357808 159480
rect 357860 159468 357866 159520
rect 217870 159400 217876 159452
rect 217928 159440 217934 159452
rect 284386 159440 284392 159452
rect 217928 159412 284392 159440
rect 217928 159400 217934 159412
rect 284386 159400 284392 159412
rect 284444 159400 284450 159452
rect 307846 159400 307852 159452
rect 307904 159440 307910 159452
rect 359366 159440 359372 159452
rect 307904 159412 359372 159440
rect 307904 159400 307910 159412
rect 359366 159400 359372 159412
rect 359424 159400 359430 159452
rect 213546 159332 213552 159384
rect 213604 159372 213610 159384
rect 281534 159372 281540 159384
rect 213604 159344 281540 159372
rect 213604 159332 213610 159344
rect 281534 159332 281540 159344
rect 281592 159332 281598 159384
rect 292574 159332 292580 159384
rect 292632 159372 292638 159384
rect 359182 159372 359188 159384
rect 292632 159344 359188 159372
rect 292632 159332 292638 159344
rect 359182 159332 359188 159344
rect 359240 159332 359246 159384
rect 355318 159264 355324 159316
rect 355376 159304 355382 159316
rect 361942 159304 361948 159316
rect 355376 159276 361948 159304
rect 355376 159264 355382 159276
rect 361942 159264 361948 159276
rect 362000 159264 362006 159316
rect 285950 159196 285956 159248
rect 286008 159236 286014 159248
rect 365162 159236 365168 159248
rect 286008 159208 365168 159236
rect 286008 159196 286014 159208
rect 365162 159196 365168 159208
rect 365220 159196 365226 159248
rect 291010 159128 291016 159180
rect 291068 159168 291074 159180
rect 371878 159168 371884 159180
rect 291068 159140 371884 159168
rect 291068 159128 291074 159140
rect 371878 159128 371884 159140
rect 371936 159128 371942 159180
rect 279234 159060 279240 159112
rect 279292 159100 279298 159112
rect 362034 159100 362040 159112
rect 279292 159072 362040 159100
rect 279292 159060 279298 159072
rect 362034 159060 362040 159072
rect 362092 159060 362098 159112
rect 277026 158992 277032 159044
rect 277084 159032 277090 159044
rect 360562 159032 360568 159044
rect 277084 159004 360568 159032
rect 277084 158992 277090 159004
rect 360562 158992 360568 159004
rect 360620 158992 360626 159044
rect 278130 158924 278136 158976
rect 278188 158964 278194 158976
rect 355318 158964 355324 158976
rect 278188 158936 355324 158964
rect 278188 158924 278194 158936
rect 355318 158924 355324 158936
rect 355376 158924 355382 158976
rect 355410 158924 355416 158976
rect 355468 158964 355474 158976
rect 360654 158964 360660 158976
rect 355468 158936 360660 158964
rect 355468 158924 355474 158936
rect 360654 158924 360660 158936
rect 360712 158924 360718 158976
rect 273346 158856 273352 158908
rect 273404 158896 273410 158908
rect 359274 158896 359280 158908
rect 273404 158868 359280 158896
rect 273404 158856 273410 158868
rect 359274 158856 359280 158868
rect 359332 158856 359338 158908
rect 214466 158788 214472 158840
rect 214524 158828 214530 158840
rect 214650 158828 214656 158840
rect 214524 158800 214656 158828
rect 214524 158788 214530 158800
rect 214650 158788 214656 158800
rect 214708 158788 214714 158840
rect 275830 158788 275836 158840
rect 275888 158828 275894 158840
rect 360746 158828 360752 158840
rect 275888 158800 360752 158828
rect 275888 158788 275894 158800
rect 360746 158788 360752 158800
rect 360804 158788 360810 158840
rect 213086 158720 213092 158772
rect 213144 158760 213150 158772
rect 239582 158760 239588 158772
rect 213144 158732 239588 158760
rect 213144 158720 213150 158732
rect 239582 158720 239588 158732
rect 239640 158720 239646 158772
rect 274450 158720 274456 158772
rect 274508 158760 274514 158772
rect 355410 158760 355416 158772
rect 274508 158732 355416 158760
rect 274508 158720 274514 158732
rect 355410 158720 355416 158732
rect 355468 158720 355474 158772
rect 355502 158720 355508 158772
rect 355560 158760 355566 158772
rect 357894 158760 357900 158772
rect 355560 158732 357900 158760
rect 355560 158720 355566 158732
rect 357894 158720 357900 158732
rect 357952 158720 357958 158772
rect 211982 158652 211988 158704
rect 212040 158692 212046 158704
rect 238110 158692 238116 158704
rect 212040 158664 238116 158692
rect 212040 158652 212046 158664
rect 238110 158652 238116 158664
rect 238168 158652 238174 158704
rect 268378 158652 268384 158704
rect 268436 158692 268442 158704
rect 373074 158692 373080 158704
rect 268436 158664 373080 158692
rect 268436 158652 268442 158664
rect 373074 158652 373080 158664
rect 373132 158652 373138 158704
rect 218974 158584 218980 158636
rect 219032 158624 219038 158636
rect 220814 158624 220820 158636
rect 219032 158596 220820 158624
rect 219032 158584 219038 158596
rect 220814 158584 220820 158596
rect 220872 158584 220878 158636
rect 224218 158584 224224 158636
rect 224276 158624 224282 158636
rect 229094 158624 229100 158636
rect 224276 158596 229100 158624
rect 224276 158584 224282 158596
rect 229094 158584 229100 158596
rect 229152 158584 229158 158636
rect 268746 158584 268752 158636
rect 268804 158624 268810 158636
rect 357618 158624 357624 158636
rect 268804 158596 357624 158624
rect 268804 158584 268810 158596
rect 357618 158584 357624 158596
rect 357676 158584 357682 158636
rect 219066 158516 219072 158568
rect 219124 158556 219130 158568
rect 234614 158556 234620 158568
rect 219124 158528 234620 158556
rect 219124 158516 219130 158528
rect 234614 158516 234620 158528
rect 234672 158516 234678 158568
rect 272242 158516 272248 158568
rect 272300 158556 272306 158568
rect 292574 158556 292580 158568
rect 272300 158528 292580 158556
rect 272300 158516 272306 158528
rect 292574 158516 292580 158528
rect 292632 158516 292638 158568
rect 298554 158516 298560 158568
rect 298612 158556 298618 158568
rect 356238 158556 356244 158568
rect 298612 158528 356244 158556
rect 298612 158516 298618 158528
rect 356238 158516 356244 158528
rect 356296 158516 356302 158568
rect 211890 158448 211896 158500
rect 211948 158488 211954 158500
rect 230474 158488 230480 158500
rect 211948 158460 230480 158488
rect 211948 158448 211954 158460
rect 230474 158448 230480 158460
rect 230532 158448 230538 158500
rect 301038 158448 301044 158500
rect 301096 158488 301102 158500
rect 357526 158488 357532 158500
rect 301096 158460 357532 158488
rect 301096 158448 301102 158460
rect 357526 158448 357532 158460
rect 357584 158448 357590 158500
rect 216306 158380 216312 158432
rect 216364 158420 216370 158432
rect 238754 158420 238760 158432
rect 216364 158392 238760 158420
rect 216364 158380 216370 158392
rect 238754 158380 238760 158392
rect 238812 158380 238818 158432
rect 303522 158380 303528 158432
rect 303580 158420 303586 158432
rect 357710 158420 357716 158432
rect 303580 158392 357716 158420
rect 303580 158380 303586 158392
rect 357710 158380 357716 158392
rect 357768 158380 357774 158432
rect 212074 158312 212080 158364
rect 212132 158352 212138 158364
rect 234706 158352 234712 158364
rect 212132 158324 234712 158352
rect 212132 158312 212138 158324
rect 234706 158312 234712 158324
rect 234764 158312 234770 158364
rect 306098 158312 306104 158364
rect 306156 158352 306162 158364
rect 359090 158352 359096 158364
rect 306156 158324 359096 158352
rect 306156 158312 306162 158324
rect 359090 158312 359096 158324
rect 359148 158312 359154 158364
rect 216214 158244 216220 158296
rect 216272 158284 216278 158296
rect 242986 158284 242992 158296
rect 216272 158256 242992 158284
rect 216272 158244 216278 158256
rect 242986 158244 242992 158256
rect 243044 158244 243050 158296
rect 271138 158244 271144 158296
rect 271196 158284 271202 158296
rect 307846 158284 307852 158296
rect 271196 158256 307852 158284
rect 271196 158244 271202 158256
rect 307846 158244 307852 158256
rect 307904 158244 307910 158296
rect 308674 158244 308680 158296
rect 308732 158284 308738 158296
rect 358906 158284 358912 158296
rect 308732 158256 358912 158284
rect 308732 158244 308738 158256
rect 358906 158244 358912 158256
rect 358964 158244 358970 158296
rect 212258 158176 212264 158228
rect 212316 158216 212322 158228
rect 241514 158216 241520 158228
rect 212316 158188 241520 158216
rect 212316 158176 212322 158188
rect 241514 158176 241520 158188
rect 241572 158176 241578 158228
rect 311066 158176 311072 158228
rect 311124 158216 311130 158228
rect 358998 158216 359004 158228
rect 311124 158188 359004 158216
rect 311124 158176 311130 158188
rect 358998 158176 359004 158188
rect 359056 158176 359062 158228
rect 216122 158108 216128 158160
rect 216180 158148 216186 158160
rect 245654 158148 245660 158160
rect 216180 158120 245660 158148
rect 216180 158108 216186 158120
rect 245654 158108 245660 158120
rect 245712 158108 245718 158160
rect 313458 158108 313464 158160
rect 313516 158148 313522 158160
rect 359642 158148 359648 158160
rect 313516 158120 359648 158148
rect 313516 158108 313522 158120
rect 359642 158108 359648 158120
rect 359700 158108 359706 158160
rect 215938 158040 215944 158092
rect 215996 158080 216002 158092
rect 247034 158080 247040 158092
rect 215996 158052 247040 158080
rect 215996 158040 216002 158052
rect 247034 158040 247040 158052
rect 247092 158040 247098 158092
rect 269850 158040 269856 158092
rect 269908 158080 269914 158092
rect 314654 158080 314660 158092
rect 269908 158052 314660 158080
rect 269908 158040 269914 158052
rect 314654 158040 314660 158052
rect 314712 158040 314718 158092
rect 315850 158040 315856 158092
rect 315908 158080 315914 158092
rect 360470 158080 360476 158092
rect 315908 158052 360476 158080
rect 315908 158040 315914 158052
rect 360470 158040 360476 158052
rect 360528 158040 360534 158092
rect 218882 157972 218888 158024
rect 218940 158012 218946 158024
rect 252554 158012 252560 158024
rect 218940 157984 252560 158012
rect 218940 157972 218946 157984
rect 252554 157972 252560 157984
rect 252612 157972 252618 158024
rect 293586 157972 293592 158024
rect 293644 158012 293650 158024
rect 317690 158012 317696 158024
rect 293644 157984 317696 158012
rect 293644 157972 293650 157984
rect 317690 157972 317696 157984
rect 317748 157972 317754 158024
rect 318610 157972 318616 158024
rect 318668 158012 318674 158024
rect 360378 158012 360384 158024
rect 318668 157984 360384 158012
rect 318668 157972 318674 157984
rect 360378 157972 360384 157984
rect 360436 157972 360442 158024
rect 214558 157904 214564 157956
rect 214616 157944 214622 157956
rect 224218 157944 224224 157956
rect 214616 157916 224224 157944
rect 214616 157904 214622 157916
rect 224218 157904 224224 157916
rect 224276 157904 224282 157956
rect 321002 157904 321008 157956
rect 321060 157944 321066 157956
rect 361022 157944 361028 157956
rect 321060 157916 361028 157944
rect 321060 157904 321066 157916
rect 361022 157904 361028 157916
rect 361080 157904 361086 157956
rect 214650 157836 214656 157888
rect 214708 157876 214714 157888
rect 219434 157876 219440 157888
rect 214708 157848 219440 157876
rect 214708 157836 214714 157848
rect 219434 157836 219440 157848
rect 219492 157836 219498 157888
rect 323394 157836 323400 157888
rect 323452 157876 323458 157888
rect 361758 157876 361764 157888
rect 323452 157848 361764 157876
rect 323452 157836 323458 157848
rect 361758 157836 361764 157848
rect 361816 157836 361822 157888
rect 325970 157768 325976 157820
rect 326028 157808 326034 157820
rect 361850 157808 361856 157820
rect 326028 157780 361856 157808
rect 326028 157768 326034 157780
rect 361850 157768 361856 157780
rect 361908 157768 361914 157820
rect 216214 157360 216220 157412
rect 216272 157400 216278 157412
rect 223574 157400 223580 157412
rect 216272 157372 223580 157400
rect 216272 157360 216278 157372
rect 223574 157360 223580 157372
rect 223632 157360 223638 157412
rect 242434 157292 242440 157344
rect 242492 157332 242498 157344
rect 367922 157332 367928 157344
rect 242492 157304 367928 157332
rect 242492 157292 242498 157304
rect 367922 157292 367928 157304
rect 367980 157292 367986 157344
rect 244274 157224 244280 157276
rect 244332 157264 244338 157276
rect 368750 157264 368756 157276
rect 244332 157236 368756 157264
rect 244332 157224 244338 157236
rect 368750 157224 368756 157236
rect 368808 157224 368814 157276
rect 248322 157156 248328 157208
rect 248380 157196 248386 157208
rect 370222 157196 370228 157208
rect 248380 157168 370228 157196
rect 248380 157156 248386 157168
rect 370222 157156 370228 157168
rect 370280 157156 370286 157208
rect 250898 157088 250904 157140
rect 250956 157128 250962 157140
rect 370498 157128 370504 157140
rect 250956 157100 370504 157128
rect 250956 157088 250962 157100
rect 370498 157088 370504 157100
rect 370556 157088 370562 157140
rect 252094 157020 252100 157072
rect 252152 157060 252158 157072
rect 371602 157060 371608 157072
rect 252152 157032 371608 157060
rect 252152 157020 252158 157032
rect 371602 157020 371608 157032
rect 371660 157020 371666 157072
rect 257338 156952 257344 157004
rect 257396 156992 257402 157004
rect 366174 156992 366180 157004
rect 257396 156964 366180 156992
rect 257396 156952 257402 156964
rect 366174 156952 366180 156964
rect 366232 156952 366238 157004
rect 261754 156884 261760 156936
rect 261812 156924 261818 156936
rect 368934 156924 368940 156936
rect 261812 156896 368940 156924
rect 261812 156884 261818 156896
rect 368934 156884 368940 156896
rect 368992 156884 368998 156936
rect 259914 156816 259920 156868
rect 259972 156856 259978 156868
rect 365070 156856 365076 156868
rect 259972 156828 365076 156856
rect 259972 156816 259978 156828
rect 365070 156816 365076 156828
rect 365128 156816 365134 156868
rect 264330 156748 264336 156800
rect 264388 156788 264394 156800
rect 368842 156788 368848 156800
rect 264388 156760 368848 156788
rect 264388 156748 264394 156760
rect 368842 156748 368848 156760
rect 368900 156748 368906 156800
rect 265894 156680 265900 156732
rect 265952 156720 265958 156732
rect 367554 156720 367560 156732
rect 265952 156692 367560 156720
rect 265952 156680 265958 156692
rect 367554 156680 367560 156692
rect 367612 156680 367618 156732
rect 271046 156612 271052 156664
rect 271104 156652 271110 156664
rect 371786 156652 371792 156664
rect 271104 156624 371792 156652
rect 271104 156612 271110 156624
rect 371786 156612 371792 156624
rect 371844 156612 371850 156664
rect 276106 156544 276112 156596
rect 276164 156584 276170 156596
rect 370130 156584 370136 156596
rect 276164 156556 370136 156584
rect 276164 156544 276170 156556
rect 370130 156544 370136 156556
rect 370188 156544 370194 156596
rect 283650 156476 283656 156528
rect 283708 156516 283714 156528
rect 371694 156516 371700 156528
rect 283708 156488 371700 156516
rect 283708 156476 283714 156488
rect 371694 156476 371700 156488
rect 371752 156476 371758 156528
rect 295978 156408 295984 156460
rect 296036 156448 296042 156460
rect 370590 156448 370596 156460
rect 296036 156420 370596 156448
rect 296036 156408 296042 156420
rect 370590 156408 370596 156420
rect 370648 156408 370654 156460
rect 240594 155864 240600 155916
rect 240652 155904 240658 155916
rect 369302 155904 369308 155916
rect 240652 155876 369308 155904
rect 240652 155864 240658 155876
rect 369302 155864 369308 155876
rect 369360 155864 369366 155916
rect 246758 155796 246764 155848
rect 246816 155836 246822 155848
rect 369026 155836 369032 155848
rect 246816 155808 369032 155836
rect 246816 155796 246822 155808
rect 369026 155796 369032 155808
rect 369084 155796 369090 155848
rect 248690 155728 248696 155780
rect 248748 155768 248754 155780
rect 369118 155768 369124 155780
rect 248748 155740 369124 155768
rect 248748 155728 248754 155740
rect 369118 155728 369124 155740
rect 369176 155728 369182 155780
rect 247770 155660 247776 155712
rect 247828 155700 247834 155712
rect 367646 155700 367652 155712
rect 247828 155672 367652 155700
rect 247828 155660 247834 155672
rect 367646 155660 367652 155672
rect 367704 155660 367710 155712
rect 218790 155592 218796 155644
rect 218848 155632 218854 155644
rect 251266 155632 251272 155644
rect 218848 155604 251272 155632
rect 218848 155592 218854 155604
rect 251266 155592 251272 155604
rect 251324 155592 251330 155644
rect 253474 155592 253480 155644
rect 253532 155632 253538 155644
rect 371418 155632 371424 155644
rect 253532 155604 371424 155632
rect 253532 155592 253538 155604
rect 371418 155592 371424 155604
rect 371476 155592 371482 155644
rect 245562 155524 245568 155576
rect 245620 155564 245626 155576
rect 362402 155564 362408 155576
rect 245620 155536 362408 155564
rect 245620 155524 245626 155536
rect 362402 155524 362408 155536
rect 362460 155524 362466 155576
rect 215846 155456 215852 155508
rect 215904 155496 215910 155508
rect 248414 155496 248420 155508
rect 215904 155468 248420 155496
rect 215904 155456 215910 155468
rect 248414 155456 248420 155468
rect 248472 155456 248478 155508
rect 250714 155456 250720 155508
rect 250772 155496 250778 155508
rect 367738 155496 367744 155508
rect 250772 155468 367744 155496
rect 250772 155456 250778 155468
rect 367738 155456 367744 155468
rect 367796 155456 367802 155508
rect 212350 155388 212356 155440
rect 212408 155428 212414 155440
rect 253934 155428 253940 155440
rect 212408 155400 253940 155428
rect 212408 155388 212414 155400
rect 253934 155388 253940 155400
rect 253992 155388 253998 155440
rect 256050 155388 256056 155440
rect 256108 155428 256114 155440
rect 372982 155428 372988 155440
rect 256108 155400 372988 155428
rect 256108 155388 256114 155400
rect 372982 155388 372988 155400
rect 373040 155388 373046 155440
rect 218698 155320 218704 155372
rect 218756 155360 218762 155372
rect 266354 155360 266360 155372
rect 218756 155332 266360 155360
rect 218756 155320 218762 155332
rect 266354 155320 266360 155332
rect 266412 155320 266418 155372
rect 266630 155320 266636 155372
rect 266688 155360 266694 155372
rect 367462 155360 367468 155372
rect 266688 155332 367468 155360
rect 266688 155320 266694 155332
rect 367462 155320 367468 155332
rect 367520 155320 367526 155372
rect 212166 155252 212172 155304
rect 212224 155292 212230 155304
rect 270494 155292 270500 155304
rect 212224 155264 270500 155292
rect 212224 155252 212230 155264
rect 270494 155252 270500 155264
rect 270552 155252 270558 155304
rect 273714 155252 273720 155304
rect 273772 155292 273778 155304
rect 371326 155292 371332 155304
rect 273772 155264 371332 155292
rect 273772 155252 273778 155264
rect 371326 155252 371332 155264
rect 371384 155252 371390 155304
rect 217502 155184 217508 155236
rect 217560 155224 217566 155236
rect 277394 155224 277400 155236
rect 217560 155196 277400 155224
rect 217560 155184 217566 155196
rect 277394 155184 277400 155196
rect 277452 155184 277458 155236
rect 278498 155184 278504 155236
rect 278556 155224 278562 155236
rect 371510 155224 371516 155236
rect 278556 155196 371516 155224
rect 278556 155184 278562 155196
rect 371510 155184 371516 155196
rect 371568 155184 371574 155236
rect 218606 155116 218612 155168
rect 218664 155156 218670 155168
rect 278774 155156 278780 155168
rect 218664 155128 278780 155156
rect 218664 155116 218670 155128
rect 278774 155116 278780 155128
rect 278832 155116 278838 155168
rect 281074 155116 281080 155168
rect 281132 155156 281138 155168
rect 370038 155156 370044 155168
rect 281132 155128 370044 155156
rect 281132 155116 281138 155128
rect 370038 155116 370044 155128
rect 370096 155116 370102 155168
rect 217134 155048 217140 155100
rect 217192 155088 217198 155100
rect 285674 155088 285680 155100
rect 217192 155060 285680 155088
rect 217192 155048 217198 155060
rect 285674 155048 285680 155060
rect 285732 155048 285738 155100
rect 288250 155048 288256 155100
rect 288308 155088 288314 155100
rect 370314 155088 370320 155100
rect 288308 155060 370320 155088
rect 288308 155048 288314 155060
rect 370314 155048 370320 155060
rect 370372 155048 370378 155100
rect 214466 154980 214472 155032
rect 214524 155020 214530 155032
rect 282914 155020 282920 155032
rect 214524 154992 282920 155020
rect 214524 154980 214530 154992
rect 282914 154980 282920 154992
rect 282972 154980 282978 155032
rect 261202 154504 261208 154556
rect 261260 154544 261266 154556
rect 372798 154544 372804 154556
rect 261260 154516 372804 154544
rect 261260 154504 261266 154516
rect 372798 154504 372804 154516
rect 372856 154504 372862 154556
rect 263686 154436 263692 154488
rect 263744 154476 263750 154488
rect 372890 154476 372896 154488
rect 263744 154448 372896 154476
rect 263744 154436 263750 154448
rect 372890 154436 372896 154448
rect 372948 154436 372954 154488
rect 265986 154368 265992 154420
rect 266044 154408 266050 154420
rect 372706 154408 372712 154420
rect 266044 154380 372712 154408
rect 266044 154368 266050 154380
rect 372706 154368 372712 154380
rect 372764 154368 372770 154420
rect 209682 152532 209688 152584
rect 209740 152572 209746 152584
rect 269114 152572 269120 152584
rect 209740 152544 269120 152572
rect 209740 152532 209746 152544
rect 269114 152532 269120 152544
rect 269172 152532 269178 152584
rect 213454 152464 213460 152516
rect 213512 152504 213518 152516
rect 273254 152504 273260 152516
rect 213512 152476 273260 152504
rect 213512 152464 213518 152476
rect 273254 152464 273260 152476
rect 273312 152464 273318 152516
rect 3602 150356 3608 150408
rect 3660 150396 3666 150408
rect 178770 150396 178776 150408
rect 3660 150368 178776 150396
rect 3660 150356 3666 150368
rect 178770 150356 178776 150368
rect 178828 150356 178834 150408
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 209038 111772 209044 111784
rect 3200 111744 209044 111772
rect 3200 111732 3206 111744
rect 209038 111732 209044 111744
rect 209096 111732 209102 111784
rect 3510 97588 3516 97640
rect 3568 97628 3574 97640
rect 7558 97628 7564 97640
rect 3568 97600 7564 97628
rect 3568 97588 3574 97600
rect 7558 97588 7564 97600
rect 7616 97588 7622 97640
rect 143534 11704 143540 11756
rect 143592 11744 143598 11756
rect 144730 11744 144736 11756
rect 143592 11716 144736 11744
rect 143592 11704 143598 11716
rect 144730 11704 144736 11716
rect 144788 11704 144794 11756
rect 168374 11704 168380 11756
rect 168432 11744 168438 11756
rect 169570 11744 169576 11756
rect 168432 11716 169576 11744
rect 168432 11704 168438 11716
rect 169570 11704 169576 11716
rect 169628 11704 169634 11756
rect 176654 11704 176660 11756
rect 176712 11744 176718 11756
rect 177850 11744 177856 11756
rect 176712 11716 177856 11744
rect 176712 11704 176718 11716
rect 177850 11704 177856 11716
rect 177908 11704 177914 11756
rect 234614 11704 234620 11756
rect 234672 11744 234678 11756
rect 235810 11744 235816 11756
rect 234672 11716 235816 11744
rect 234672 11704 234678 11716
rect 235810 11704 235816 11716
rect 235868 11704 235874 11756
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 307938 9596 307944 9648
rect 307996 9636 308002 9648
rect 369854 9636 369860 9648
rect 307996 9608 369860 9636
rect 307996 9596 308002 9608
rect 369854 9596 369860 9608
rect 369912 9596 369918 9648
rect 306742 9528 306748 9580
rect 306800 9568 306806 9580
rect 368658 9568 368664 9580
rect 306800 9540 368664 9568
rect 306800 9528 306806 9540
rect 368658 9528 368664 9540
rect 368716 9528 368722 9580
rect 305546 9460 305552 9512
rect 305604 9500 305610 9512
rect 367370 9500 367376 9512
rect 305604 9472 367376 9500
rect 305604 9460 305610 9472
rect 367370 9460 367376 9472
rect 367428 9460 367434 9512
rect 304350 9392 304356 9444
rect 304408 9432 304414 9444
rect 366082 9432 366088 9444
rect 304408 9404 366088 9432
rect 304408 9392 304414 9404
rect 366082 9392 366088 9404
rect 366140 9392 366146 9444
rect 299658 9324 299664 9376
rect 299716 9364 299722 9376
rect 362310 9364 362316 9376
rect 299716 9336 362316 9364
rect 299716 9324 299722 9336
rect 362310 9324 362316 9336
rect 362368 9324 362374 9376
rect 297266 9256 297272 9308
rect 297324 9296 297330 9308
rect 359550 9296 359556 9308
rect 297324 9268 359556 9296
rect 297324 9256 297330 9268
rect 359550 9256 359556 9268
rect 359608 9256 359614 9308
rect 301958 9188 301964 9240
rect 302016 9228 302022 9240
rect 369946 9228 369952 9240
rect 302016 9200 369952 9228
rect 302016 9188 302022 9200
rect 369946 9188 369952 9200
rect 370004 9188 370010 9240
rect 298462 9120 298468 9172
rect 298520 9160 298526 9172
rect 367278 9160 367284 9172
rect 298520 9132 367284 9160
rect 298520 9120 298526 9132
rect 367278 9120 367284 9132
rect 367336 9120 367342 9172
rect 296070 9052 296076 9104
rect 296128 9092 296134 9104
rect 364978 9092 364984 9104
rect 296128 9064 364984 9092
rect 296128 9052 296134 9064
rect 364978 9052 364984 9064
rect 365036 9052 365042 9104
rect 294874 8984 294880 9036
rect 294932 9024 294938 9036
rect 363598 9024 363604 9036
rect 294932 8996 363604 9024
rect 294932 8984 294938 8996
rect 363598 8984 363604 8996
rect 363656 8984 363662 9036
rect 293678 8916 293684 8968
rect 293736 8956 293742 8968
rect 368566 8956 368572 8968
rect 293736 8928 368572 8956
rect 293736 8916 293742 8928
rect 368566 8916 368572 8928
rect 368624 8916 368630 8968
rect 300762 8848 300768 8900
rect 300820 8888 300826 8900
rect 360930 8888 360936 8900
rect 300820 8860 360936 8888
rect 300820 8848 300826 8860
rect 360930 8848 360936 8860
rect 360988 8848 360994 8900
rect 303154 8780 303160 8832
rect 303212 8820 303218 8832
rect 363506 8820 363512 8832
rect 303212 8792 363512 8820
rect 303212 8780 303218 8792
rect 363506 8780 363512 8792
rect 363564 8780 363570 8832
rect 316218 8712 316224 8764
rect 316276 8752 316282 8764
rect 364886 8752 364892 8764
rect 316276 8724 364892 8752
rect 316276 8712 316282 8724
rect 364886 8712 364892 8724
rect 364944 8712 364950 8764
rect 323302 6808 323308 6860
rect 323360 6848 323366 6860
rect 358170 6848 358176 6860
rect 323360 6820 358176 6848
rect 323360 6808 323366 6820
rect 358170 6808 358176 6820
rect 358228 6808 358234 6860
rect 317322 6740 317328 6792
rect 317380 6780 317386 6792
rect 360838 6780 360844 6792
rect 317380 6752 360844 6780
rect 317380 6740 317386 6752
rect 360838 6740 360844 6752
rect 360896 6740 360902 6792
rect 320910 6672 320916 6724
rect 320968 6712 320974 6724
rect 365806 6712 365812 6724
rect 320968 6684 365812 6712
rect 320968 6672 320974 6684
rect 365806 6672 365812 6684
rect 365864 6672 365870 6724
rect 318518 6604 318524 6656
rect 318576 6644 318582 6656
rect 363414 6644 363420 6656
rect 318576 6616 363420 6644
rect 318576 6604 318582 6616
rect 363414 6604 363420 6616
rect 363472 6604 363478 6656
rect 313826 6536 313832 6588
rect 313884 6576 313890 6588
rect 359458 6576 359464 6588
rect 313884 6548 359464 6576
rect 313884 6536 313890 6548
rect 359458 6536 359464 6548
rect 359516 6536 359522 6588
rect 315022 6468 315028 6520
rect 315080 6508 315086 6520
rect 362126 6508 362132 6520
rect 315080 6480 362132 6508
rect 315080 6468 315086 6480
rect 362126 6468 362132 6480
rect 362184 6468 362190 6520
rect 312630 6400 312636 6452
rect 312688 6440 312694 6452
rect 360194 6440 360200 6452
rect 312688 6412 360200 6440
rect 312688 6400 312694 6412
rect 360194 6400 360200 6412
rect 360252 6400 360258 6452
rect 311434 6332 311440 6384
rect 311492 6372 311498 6384
rect 358814 6372 358820 6384
rect 311492 6344 358820 6372
rect 311492 6332 311498 6344
rect 358814 6332 358820 6344
rect 358872 6332 358878 6384
rect 310238 6264 310244 6316
rect 310296 6304 310302 6316
rect 358262 6304 358268 6316
rect 310296 6276 358268 6304
rect 310296 6264 310302 6276
rect 358262 6264 358268 6276
rect 358320 6264 358326 6316
rect 309042 6196 309048 6248
rect 309100 6236 309106 6248
rect 368474 6236 368480 6248
rect 309100 6208 368480 6236
rect 309100 6196 309106 6208
rect 368474 6196 368480 6208
rect 368532 6196 368538 6248
rect 292574 6128 292580 6180
rect 292632 6168 292638 6180
rect 362218 6168 362224 6180
rect 292632 6140 362224 6168
rect 292632 6128 292638 6140
rect 362218 6128 362224 6140
rect 362276 6128 362282 6180
rect 326798 6060 326804 6112
rect 326856 6100 326862 6112
rect 360286 6100 360292 6112
rect 326856 6072 360292 6100
rect 326856 6060 326862 6072
rect 360286 6060 360292 6072
rect 360344 6060 360350 6112
rect 330386 5992 330392 6044
rect 330444 6032 330450 6044
rect 363138 6032 363144 6044
rect 330444 6004 363144 6032
rect 330444 5992 330450 6004
rect 363138 5992 363144 6004
rect 363196 5992 363202 6044
rect 333882 5924 333888 5976
rect 333940 5964 333946 5976
rect 364794 5964 364800 5976
rect 333940 5936 364800 5964
rect 333940 5924 333946 5936
rect 364794 5924 364800 5936
rect 364852 5924 364858 5976
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 7742 4128 7748 4140
rect 2924 4100 7748 4128
rect 2924 4088 2930 4100
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17218 4128 17224 4140
rect 15988 4100 17224 4128
rect 15988 4088 15994 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 24210 4088 24216 4140
rect 24268 4128 24274 4140
rect 26878 4128 26884 4140
rect 24268 4100 26884 4128
rect 24268 4088 24274 4100
rect 26878 4088 26884 4100
rect 26936 4088 26942 4140
rect 213730 4088 213736 4140
rect 213788 4128 213794 4140
rect 260650 4128 260656 4140
rect 213788 4100 260656 4128
rect 213788 4088 213794 4100
rect 260650 4088 260656 4100
rect 260708 4088 260714 4140
rect 354030 4088 354036 4140
rect 354088 4128 354094 4140
rect 365254 4128 365260 4140
rect 354088 4100 365260 4128
rect 354088 4088 354094 4100
rect 365254 4088 365260 4100
rect 365312 4088 365318 4140
rect 217318 4020 217324 4072
rect 217376 4060 217382 4072
rect 276014 4060 276020 4072
rect 217376 4032 276020 4060
rect 217376 4020 217382 4032
rect 276014 4020 276020 4032
rect 276072 4020 276078 4072
rect 346946 4020 346952 4072
rect 347004 4060 347010 4072
rect 364610 4060 364616 4072
rect 347004 4032 364616 4060
rect 347004 4020 347010 4032
rect 364610 4020 364616 4032
rect 364668 4020 364674 4072
rect 214742 3952 214748 4004
rect 214800 3992 214806 4004
rect 262950 3992 262956 4004
rect 214800 3964 262956 3992
rect 214800 3952 214806 3964
rect 262950 3952 262956 3964
rect 263008 3952 263014 4004
rect 342162 3952 342168 4004
rect 342220 3992 342226 4004
rect 362494 3992 362500 4004
rect 342220 3964 362500 3992
rect 342220 3952 342226 3964
rect 362494 3952 362500 3964
rect 362552 3952 362558 4004
rect 503070 3952 503076 4004
rect 503128 3992 503134 4004
rect 537202 3992 537208 4004
rect 503128 3964 537208 3992
rect 503128 3952 503134 3964
rect 537202 3952 537208 3964
rect 537260 3952 537266 4004
rect 216490 3884 216496 3936
rect 216548 3924 216554 3936
rect 277118 3924 277124 3936
rect 216548 3896 277124 3924
rect 216548 3884 216554 3896
rect 277118 3884 277124 3896
rect 277176 3884 277182 3936
rect 343358 3884 343364 3936
rect 343416 3924 343422 3936
rect 362954 3924 362960 3936
rect 343416 3896 362960 3924
rect 343416 3884 343422 3896
rect 362954 3884 362960 3896
rect 363012 3884 363018 3936
rect 496078 3884 496084 3936
rect 496136 3924 496142 3936
rect 533706 3924 533712 3936
rect 496136 3896 533712 3924
rect 496136 3884 496142 3896
rect 533706 3884 533712 3896
rect 533764 3884 533770 3936
rect 211062 3816 211068 3868
rect 211120 3856 211126 3868
rect 272426 3856 272432 3868
rect 211120 3828 272432 3856
rect 211120 3816 211126 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 339862 3816 339868 3868
rect 339920 3856 339926 3868
rect 364426 3856 364432 3868
rect 339920 3828 364432 3856
rect 339920 3816 339926 3828
rect 364426 3816 364432 3828
rect 364484 3816 364490 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 554958 3856 554964 3868
rect 516836 3828 554964 3856
rect 516836 3816 516842 3828
rect 554958 3816 554964 3828
rect 555016 3816 555022 3868
rect 219158 3748 219164 3800
rect 219216 3788 219222 3800
rect 280706 3788 280712 3800
rect 219216 3760 280712 3788
rect 219216 3748 219222 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 336274 3748 336280 3800
rect 336332 3788 336338 3800
rect 364518 3788 364524 3800
rect 336332 3760 364524 3788
rect 336332 3748 336338 3760
rect 364518 3748 364524 3760
rect 364576 3748 364582 3800
rect 476758 3748 476764 3800
rect 476816 3788 476822 3800
rect 523034 3788 523040 3800
rect 476816 3760 523040 3788
rect 476816 3748 476822 3760
rect 523034 3748 523040 3760
rect 523092 3748 523098 3800
rect 538950 3748 538956 3800
rect 539008 3788 539014 3800
rect 559742 3788 559748 3800
rect 539008 3760 559748 3788
rect 539008 3748 539014 3760
rect 559742 3748 559748 3760
rect 559800 3748 559806 3800
rect 35986 3680 35992 3732
rect 36044 3720 36050 3732
rect 46198 3720 46204 3732
rect 36044 3692 46204 3720
rect 36044 3680 36050 3692
rect 46198 3680 46204 3692
rect 46256 3680 46262 3732
rect 219342 3680 219348 3732
rect 219400 3720 219406 3732
rect 287790 3720 287796 3732
rect 219400 3692 287796 3720
rect 219400 3680 219406 3692
rect 287790 3680 287796 3692
rect 287848 3680 287854 3732
rect 332686 3680 332692 3732
rect 332744 3720 332750 3732
rect 364334 3720 364340 3732
rect 332744 3692 364340 3720
rect 332744 3680 332750 3692
rect 364334 3680 364340 3692
rect 364392 3680 364398 3732
rect 431218 3680 431224 3732
rect 431276 3720 431282 3732
rect 479334 3720 479340 3732
rect 431276 3692 479340 3720
rect 431276 3680 431282 3692
rect 479334 3680 479340 3692
rect 479392 3680 479398 3732
rect 508498 3680 508504 3732
rect 508556 3720 508562 3732
rect 551462 3720 551468 3732
rect 508556 3692 551468 3720
rect 508556 3680 508562 3692
rect 551462 3680 551468 3692
rect 551520 3680 551526 3732
rect 43438 3652 43444 3664
rect 26206 3624 43444 3652
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13078 3584 13084 3596
rect 12400 3556 13084 3584
rect 12400 3544 12406 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 26206 3584 26234 3624
rect 43438 3612 43444 3624
rect 43496 3612 43502 3664
rect 46658 3612 46664 3664
rect 46716 3652 46722 3664
rect 46716 3624 55214 3652
rect 46716 3612 46722 3624
rect 20680 3556 26234 3584
rect 20680 3544 20686 3556
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 32398 3584 32404 3596
rect 28960 3556 32404 3584
rect 28960 3544 28966 3556
rect 32398 3544 32404 3556
rect 32456 3544 32462 3596
rect 38378 3544 38384 3596
rect 38436 3584 38442 3596
rect 39298 3584 39304 3596
rect 38436 3556 39304 3584
rect 38436 3544 38442 3556
rect 39298 3544 39304 3556
rect 39356 3544 39362 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 53098 3584 53104 3596
rect 51408 3556 53104 3584
rect 51408 3544 51414 3556
rect 53098 3544 53104 3556
rect 53156 3544 53162 3596
rect 53742 3544 53748 3596
rect 53800 3584 53806 3596
rect 54478 3584 54484 3596
rect 53800 3556 54484 3584
rect 53800 3544 53806 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 55186 3584 55214 3624
rect 60826 3612 60832 3664
rect 60884 3652 60890 3664
rect 79318 3652 79324 3664
rect 60884 3624 79324 3652
rect 60884 3612 60890 3624
rect 79318 3612 79324 3624
rect 79376 3612 79382 3664
rect 85666 3612 85672 3664
rect 85724 3652 85730 3664
rect 106918 3652 106924 3664
rect 85724 3624 106924 3652
rect 85724 3612 85730 3624
rect 106918 3612 106924 3624
rect 106976 3612 106982 3664
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 182818 3652 182824 3664
rect 114060 3624 182824 3652
rect 114060 3612 114066 3624
rect 182818 3612 182824 3624
rect 182876 3612 182882 3664
rect 189718 3652 189724 3664
rect 184216 3624 189724 3652
rect 116578 3584 116584 3596
rect 55186 3556 116584 3584
rect 116578 3544 116584 3556
rect 116636 3544 116642 3596
rect 118694 3544 118700 3596
rect 118752 3584 118758 3596
rect 119890 3584 119896 3596
rect 118752 3556 119896 3584
rect 118752 3544 118758 3556
rect 119890 3544 119896 3556
rect 119948 3544 119954 3596
rect 121086 3544 121092 3596
rect 121144 3584 121150 3596
rect 184216 3584 184244 3624
rect 189718 3612 189724 3624
rect 189776 3612 189782 3664
rect 216398 3612 216404 3664
rect 216456 3652 216462 3664
rect 284294 3652 284300 3664
rect 216456 3624 284300 3652
rect 216456 3612 216462 3624
rect 284294 3612 284300 3624
rect 284352 3612 284358 3664
rect 325602 3612 325608 3664
rect 325660 3652 325666 3664
rect 358354 3652 358360 3664
rect 325660 3624 358360 3652
rect 325660 3612 325666 3624
rect 358354 3612 358360 3624
rect 358412 3612 358418 3664
rect 457438 3612 457444 3664
rect 457496 3652 457502 3664
rect 457496 3624 460934 3652
rect 457496 3612 457502 3624
rect 121144 3556 184244 3584
rect 121144 3544 121150 3556
rect 187326 3544 187332 3596
rect 187384 3584 187390 3596
rect 188338 3584 188344 3596
rect 187384 3556 188344 3584
rect 187384 3544 187390 3556
rect 188338 3544 188344 3556
rect 188396 3544 188402 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 194410 3584 194416 3596
rect 193272 3556 194416 3584
rect 193272 3544 193278 3556
rect 194410 3544 194416 3556
rect 194468 3544 194474 3596
rect 195606 3544 195612 3596
rect 195664 3584 195670 3596
rect 196618 3584 196624 3596
rect 195664 3556 196624 3584
rect 195664 3544 195670 3556
rect 196618 3544 196624 3556
rect 196676 3544 196682 3596
rect 219342 3544 219348 3596
rect 219400 3584 219406 3596
rect 288986 3584 288992 3596
rect 219400 3556 288992 3584
rect 219400 3544 219406 3556
rect 288986 3544 288992 3556
rect 289044 3544 289050 3596
rect 329190 3544 329196 3596
rect 329248 3584 329254 3596
rect 355502 3584 355508 3596
rect 329248 3556 355508 3584
rect 329248 3544 329254 3556
rect 355502 3544 355508 3556
rect 355560 3544 355566 3596
rect 358078 3584 358084 3596
rect 355612 3556 358084 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 75178 3516 75184 3528
rect 5316 3488 75184 3516
rect 5316 3476 5322 3488
rect 75178 3476 75184 3488
rect 75236 3476 75242 3528
rect 77294 3476 77300 3528
rect 77352 3516 77358 3528
rect 78214 3516 78220 3528
rect 77352 3488 78220 3516
rect 77352 3476 77358 3488
rect 78214 3476 78220 3488
rect 78272 3476 78278 3528
rect 93854 3476 93860 3528
rect 93912 3516 93918 3528
rect 94774 3516 94780 3528
rect 93912 3488 94780 3516
rect 93912 3476 93918 3488
rect 94774 3476 94780 3488
rect 94832 3476 94838 3528
rect 102134 3476 102140 3528
rect 102192 3516 102198 3528
rect 103330 3516 103336 3528
rect 102192 3488 103336 3516
rect 102192 3476 102198 3488
rect 103330 3476 103336 3488
rect 103388 3476 103394 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 178678 3516 178684 3528
rect 106976 3488 178684 3516
rect 106976 3476 106982 3488
rect 178678 3476 178684 3488
rect 178736 3476 178742 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 192478 3516 192484 3528
rect 190880 3488 192484 3516
rect 190880 3476 190886 3488
rect 192478 3476 192484 3488
rect 192536 3476 192542 3528
rect 217410 3476 217416 3528
rect 217468 3516 217474 3528
rect 291378 3516 291384 3528
rect 217468 3488 291384 3516
rect 217468 3476 217474 3488
rect 291378 3476 291384 3488
rect 291436 3476 291442 3528
rect 324406 3476 324412 3528
rect 324464 3516 324470 3528
rect 355612 3516 355640 3556
rect 358078 3544 358084 3556
rect 358136 3544 358142 3596
rect 377398 3544 377404 3596
rect 377456 3544 377462 3596
rect 411898 3584 411904 3596
rect 393286 3556 411904 3584
rect 356698 3516 356704 3528
rect 324464 3488 355640 3516
rect 355704 3488 356704 3516
rect 324464 3476 324470 3488
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 8938 3448 8944 3460
rect 6512 3420 8944 3448
rect 6512 3408 6518 3420
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11204 3420 26234 3448
rect 11204 3408 11210 3420
rect 26206 3312 26234 3420
rect 30098 3408 30104 3460
rect 30156 3448 30162 3460
rect 31018 3448 31024 3460
rect 30156 3420 31024 3448
rect 30156 3408 30162 3420
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 35250 3448 35256 3460
rect 33652 3420 35256 3448
rect 33652 3408 33658 3420
rect 35250 3408 35256 3420
rect 35308 3408 35314 3460
rect 43070 3408 43076 3460
rect 43128 3448 43134 3460
rect 68278 3448 68284 3460
rect 43128 3420 68284 3448
rect 43128 3408 43134 3420
rect 68278 3408 68284 3420
rect 68336 3408 68342 3460
rect 69014 3408 69020 3460
rect 69072 3448 69078 3460
rect 69934 3448 69940 3460
rect 69072 3420 69940 3448
rect 69072 3408 69078 3420
rect 69934 3408 69940 3420
rect 69992 3408 69998 3460
rect 99834 3408 99840 3460
rect 99892 3448 99898 3460
rect 174538 3448 174544 3460
rect 99892 3420 174544 3448
rect 99892 3408 99898 3420
rect 174538 3408 174544 3420
rect 174596 3408 174602 3460
rect 182542 3408 182548 3460
rect 182600 3448 182606 3460
rect 211798 3448 211804 3460
rect 182600 3420 211804 3448
rect 182600 3408 182606 3420
rect 211798 3408 211804 3420
rect 211856 3408 211862 3460
rect 213638 3408 213644 3460
rect 213696 3448 213702 3460
rect 290182 3448 290188 3460
rect 213696 3420 290188 3448
rect 213696 3408 213702 3420
rect 290182 3408 290188 3420
rect 290240 3408 290246 3460
rect 322106 3408 322112 3460
rect 322164 3448 322170 3460
rect 355704 3448 355732 3488
rect 356698 3476 356704 3488
rect 356756 3476 356762 3528
rect 373994 3476 374000 3528
rect 374052 3516 374058 3528
rect 375282 3516 375288 3528
rect 374052 3488 375288 3516
rect 374052 3476 374058 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 377416 3516 377444 3544
rect 393286 3516 393314 3556
rect 411898 3544 411904 3556
rect 411956 3544 411962 3596
rect 442258 3544 442264 3596
rect 442316 3584 442322 3596
rect 442316 3556 451274 3584
rect 442316 3544 442322 3556
rect 377416 3488 393314 3516
rect 398834 3476 398840 3528
rect 398892 3516 398898 3528
rect 400122 3516 400128 3528
rect 398892 3488 400128 3516
rect 398892 3476 398898 3488
rect 400122 3476 400128 3488
rect 400180 3476 400186 3528
rect 407114 3476 407120 3528
rect 407172 3516 407178 3528
rect 408402 3516 408408 3528
rect 407172 3488 408408 3516
rect 407172 3476 407178 3488
rect 408402 3476 408408 3488
rect 408460 3476 408466 3528
rect 415486 3476 415492 3528
rect 415544 3516 415550 3528
rect 416682 3516 416688 3528
rect 415544 3488 416688 3516
rect 415544 3476 415550 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 423674 3476 423680 3528
rect 423732 3516 423738 3528
rect 424962 3516 424968 3528
rect 423732 3488 424968 3516
rect 423732 3476 423738 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 432046 3476 432052 3528
rect 432104 3516 432110 3528
rect 433242 3516 433248 3528
rect 432104 3488 433248 3516
rect 432104 3476 432110 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 440326 3476 440332 3528
rect 440384 3516 440390 3528
rect 441522 3516 441528 3528
rect 440384 3488 441528 3516
rect 440384 3476 440390 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 448606 3476 448612 3528
rect 448664 3516 448670 3528
rect 449802 3516 449808 3528
rect 448664 3488 449808 3516
rect 448664 3476 448670 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 451246 3516 451274 3556
rect 456794 3544 456800 3596
rect 456852 3584 456858 3596
rect 458082 3584 458088 3596
rect 456852 3556 458088 3584
rect 456852 3544 456858 3556
rect 458082 3544 458088 3556
rect 458140 3544 458146 3596
rect 460906 3584 460934 3624
rect 467098 3612 467104 3664
rect 467156 3652 467162 3664
rect 519538 3652 519544 3664
rect 467156 3624 519544 3652
rect 467156 3612 467162 3624
rect 519538 3612 519544 3624
rect 519596 3612 519602 3664
rect 534718 3612 534724 3664
rect 534776 3652 534782 3664
rect 541986 3652 541992 3664
rect 534776 3624 541992 3652
rect 534776 3612 534782 3624
rect 541986 3612 541992 3624
rect 542044 3612 542050 3664
rect 552750 3612 552756 3664
rect 552808 3652 552814 3664
rect 573910 3652 573916 3664
rect 552808 3624 573916 3652
rect 552808 3612 552814 3624
rect 573910 3612 573916 3624
rect 573968 3612 573974 3664
rect 515950 3584 515956 3596
rect 460906 3556 515956 3584
rect 515950 3544 515956 3556
rect 516008 3544 516014 3596
rect 525058 3544 525064 3596
rect 525116 3544 525122 3596
rect 531314 3544 531320 3596
rect 531372 3584 531378 3596
rect 532142 3584 532148 3596
rect 531372 3556 532148 3584
rect 531372 3544 531378 3556
rect 532142 3544 532148 3556
rect 532200 3544 532206 3596
rect 538858 3544 538864 3596
rect 538916 3584 538922 3596
rect 583386 3584 583392 3596
rect 538916 3556 583392 3584
rect 538916 3544 538922 3556
rect 583386 3544 583392 3556
rect 583444 3544 583450 3596
rect 505370 3516 505376 3528
rect 451246 3488 505376 3516
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 525076 3516 525104 3544
rect 572714 3516 572720 3528
rect 525076 3488 572720 3516
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 322164 3420 355732 3448
rect 322164 3408 322170 3420
rect 356330 3408 356336 3460
rect 356388 3448 356394 3460
rect 363046 3448 363052 3460
rect 356388 3420 363052 3448
rect 356388 3408 356394 3420
rect 363046 3408 363052 3420
rect 363104 3408 363110 3460
rect 382274 3408 382280 3460
rect 382332 3448 382338 3460
rect 383562 3448 383568 3460
rect 382332 3420 383568 3448
rect 382332 3408 382338 3420
rect 383562 3408 383568 3420
rect 383620 3408 383626 3460
rect 390554 3408 390560 3460
rect 390612 3448 390618 3460
rect 391842 3448 391848 3460
rect 390612 3420 391848 3448
rect 390612 3408 390618 3420
rect 391842 3408 391848 3420
rect 391900 3408 391906 3460
rect 429654 3448 429660 3460
rect 393286 3420 429660 3448
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 36538 3380 36544 3392
rect 34848 3352 36544 3380
rect 34848 3340 34854 3352
rect 36538 3340 36544 3352
rect 36596 3340 36602 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 57238 3380 57244 3392
rect 56100 3352 57244 3380
rect 56100 3340 56106 3352
rect 57238 3340 57244 3352
rect 57296 3340 57302 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 61378 3380 61384 3392
rect 59688 3352 61384 3380
rect 59688 3340 59694 3352
rect 61378 3340 61384 3352
rect 61436 3340 61442 3392
rect 212442 3340 212448 3392
rect 212500 3380 212506 3392
rect 258258 3380 258264 3392
rect 212500 3352 258264 3380
rect 212500 3340 212506 3352
rect 258258 3340 258264 3352
rect 258316 3340 258322 3392
rect 355226 3340 355232 3392
rect 355284 3380 355290 3392
rect 365898 3380 365904 3392
rect 355284 3352 365904 3380
rect 355284 3340 355290 3352
rect 365898 3340 365904 3352
rect 365956 3340 365962 3392
rect 387058 3340 387064 3392
rect 387116 3380 387122 3392
rect 393286 3380 393314 3420
rect 429654 3408 429660 3420
rect 429712 3408 429718 3460
rect 432598 3408 432604 3460
rect 432656 3448 432662 3460
rect 501782 3448 501788 3460
rect 432656 3420 501788 3448
rect 432656 3408 432662 3420
rect 501782 3408 501788 3420
rect 501840 3408 501846 3460
rect 520918 3408 520924 3460
rect 520976 3448 520982 3460
rect 569126 3448 569132 3460
rect 520976 3420 569132 3448
rect 520976 3408 520982 3420
rect 569126 3408 569132 3420
rect 569184 3408 569190 3460
rect 387116 3352 393314 3380
rect 387116 3340 387122 3352
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474182 3380 474188 3392
rect 473412 3352 474188 3380
rect 473412 3340 473418 3352
rect 474182 3340 474188 3352
rect 474240 3340 474246 3392
rect 481634 3340 481640 3392
rect 481692 3380 481698 3392
rect 482462 3380 482468 3392
rect 481692 3352 482468 3380
rect 481692 3340 481698 3352
rect 482462 3340 482468 3352
rect 482520 3340 482526 3392
rect 498194 3340 498200 3392
rect 498252 3380 498258 3392
rect 499022 3380 499028 3392
rect 498252 3352 499028 3380
rect 498252 3340 498258 3352
rect 499022 3340 499028 3352
rect 499080 3340 499086 3392
rect 547874 3340 547880 3392
rect 547932 3380 547938 3392
rect 548702 3380 548708 3392
rect 547932 3352 548708 3380
rect 547932 3340 547938 3352
rect 548702 3340 548708 3352
rect 548760 3340 548766 3392
rect 556154 3340 556160 3392
rect 556212 3380 556218 3392
rect 556982 3380 556988 3392
rect 556212 3352 556988 3380
rect 556212 3340 556218 3352
rect 556982 3340 556988 3352
rect 557040 3340 557046 3392
rect 35158 3312 35164 3324
rect 26206 3284 35164 3312
rect 35158 3272 35164 3284
rect 35216 3272 35222 3324
rect 213822 3272 213828 3324
rect 213880 3312 213886 3324
rect 245194 3312 245200 3324
rect 213880 3284 245200 3312
rect 213880 3272 213886 3284
rect 245194 3272 245200 3284
rect 245252 3272 245258 3324
rect 355502 3272 355508 3324
rect 355560 3312 355566 3324
rect 361666 3312 361672 3324
rect 355560 3284 361672 3312
rect 355560 3272 355566 3284
rect 361666 3272 361672 3284
rect 361724 3272 361730 3324
rect 47854 3204 47860 3256
rect 47912 3244 47918 3256
rect 48958 3244 48964 3256
rect 47912 3216 48964 3244
rect 47912 3204 47918 3216
rect 48958 3204 48964 3216
rect 49016 3204 49022 3256
rect 215202 3204 215208 3256
rect 215260 3244 215266 3256
rect 244090 3244 244096 3256
rect 215260 3216 244096 3244
rect 215260 3204 215266 3216
rect 244090 3204 244096 3216
rect 244148 3204 244154 3256
rect 352834 3204 352840 3256
rect 352892 3244 352898 3256
rect 357434 3244 357440 3256
rect 352892 3216 357440 3244
rect 352892 3204 352898 3216
rect 357434 3204 357440 3216
rect 357492 3204 357498 3256
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 4890 3176 4896 3188
rect 1728 3148 4896 3176
rect 1728 3136 1734 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 205082 3136 205088 3188
rect 205140 3176 205146 3188
rect 206278 3176 206284 3188
rect 205140 3148 206284 3176
rect 205140 3136 205146 3148
rect 206278 3136 206284 3148
rect 206336 3136 206342 3188
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 25498 2972 25504 2984
rect 19484 2944 25504 2972
rect 19484 2932 19490 2944
rect 25498 2932 25504 2944
rect 25556 2932 25562 2984
rect 41874 2932 41880 2984
rect 41932 2972 41938 2984
rect 43530 2972 43536 2984
rect 41932 2944 43536 2972
rect 41932 2932 41938 2944
rect 43530 2932 43536 2944
rect 43588 2932 43594 2984
rect 365714 1232 365720 1284
rect 365772 1272 365778 1284
rect 367002 1272 367008 1284
rect 365772 1244 367008 1272
rect 365772 1232 365778 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 348792 700476 348844 700528
rect 357532 700476 357584 700528
rect 300124 700408 300176 700460
rect 358912 700408 358964 700460
rect 361028 700408 361080 700460
rect 397460 700408 397512 700460
rect 283840 700340 283892 700392
rect 357440 700340 357492 700392
rect 360936 700340 360988 700392
rect 429844 700340 429896 700392
rect 267648 700272 267700 700324
rect 358820 700272 358872 700324
rect 360844 700272 360896 700324
rect 559656 700272 559708 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 362224 696940 362276 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 359464 670692 359516 670744
rect 580172 670692 580224 670744
rect 2780 656956 2832 657008
rect 4896 656956 4948 657008
rect 361120 643084 361172 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4988 632068 5040 632120
rect 3516 618264 3568 618316
rect 32404 618264 32456 618316
rect 358084 616836 358136 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 10324 605820 10376 605872
rect 3516 579776 3568 579828
rect 8944 579776 8996 579828
rect 3240 565836 3292 565888
rect 84844 565836 84896 565888
rect 217968 565088 218020 565140
rect 234620 565088 234672 565140
rect 331220 565088 331272 565140
rect 359004 565088 359056 565140
rect 371884 563048 371936 563100
rect 579804 563048 579856 563100
rect 2780 553664 2832 553716
rect 5080 553664 5132 553716
rect 358176 536800 358228 536852
rect 579620 536800 579672 536852
rect 2964 527144 3016 527196
rect 10416 527144 10468 527196
rect 358268 484372 358320 484424
rect 580172 484372 580224 484424
rect 219072 478184 219124 478236
rect 248420 478184 248472 478236
rect 217692 478116 217744 478168
rect 251180 478116 251232 478168
rect 311900 478116 311952 478168
rect 357532 478116 357584 478168
rect 258356 476688 258408 476740
rect 256608 476620 256660 476672
rect 260104 476620 260156 476672
rect 241612 476552 241664 476604
rect 252560 476552 252612 476604
rect 252652 476552 252704 476604
rect 263600 476552 263652 476604
rect 236092 476416 236144 476468
rect 247040 476484 247092 476536
rect 238852 476416 238904 476468
rect 244280 476416 244332 476468
rect 249800 476484 249852 476536
rect 255320 476484 255372 476536
rect 264980 476484 265032 476536
rect 238760 476348 238812 476400
rect 253848 476416 253900 476468
rect 258080 476416 258132 476468
rect 259552 476416 259604 476468
rect 278780 476688 278832 476740
rect 302240 476688 302292 476740
rect 280344 476620 280396 476672
rect 305000 476620 305052 476672
rect 284300 476552 284352 476604
rect 310520 476552 310572 476604
rect 281540 476484 281592 476536
rect 307760 476484 307812 476536
rect 245752 476348 245804 476400
rect 255412 476348 255464 476400
rect 260932 476348 260984 476400
rect 267832 476416 267884 476468
rect 285680 476416 285732 476468
rect 313280 476416 313332 476468
rect 234620 476280 234672 476332
rect 242900 476280 242952 476332
rect 248512 476280 248564 476332
rect 258264 476280 258316 476332
rect 260748 476280 260800 476332
rect 265624 476280 265676 476332
rect 270500 476348 270552 476400
rect 287060 476348 287112 476400
rect 314660 476348 314712 476400
rect 273260 476280 273312 476332
rect 288440 476280 288492 476332
rect 317420 476280 317472 476332
rect 241520 476212 241572 476264
rect 244280 476212 244332 476264
rect 251272 476212 251324 476264
rect 260840 476212 260892 476264
rect 263692 476212 263744 476264
rect 277768 476212 277820 476264
rect 289912 476212 289964 476264
rect 320180 476212 320232 476264
rect 242808 476144 242860 476196
rect 244924 476144 244976 476196
rect 251088 476144 251140 476196
rect 252652 476144 252704 476196
rect 258172 476144 258224 476196
rect 261484 476144 261536 476196
rect 262220 476144 262272 476196
rect 234712 476076 234764 476128
rect 235908 476076 235960 476128
rect 241428 476076 241480 476128
rect 242900 476076 242952 476128
rect 244372 476076 244424 476128
rect 245660 476076 245712 476128
rect 252376 476076 252428 476128
rect 253940 476076 253992 476128
rect 260748 476076 260800 476128
rect 262864 476076 262916 476128
rect 265164 476144 265216 476196
rect 280160 476144 280212 476196
rect 291200 476144 291252 476196
rect 322940 476144 322992 476196
rect 276020 476076 276072 476128
rect 292580 476076 292632 476128
rect 325792 476076 325844 476128
rect 217324 475328 217376 475380
rect 231860 475328 231912 475380
rect 273168 475328 273220 475380
rect 282920 475328 282972 475380
rect 3056 474716 3108 474768
rect 332600 474716 332652 474768
rect 219164 474036 219216 474088
rect 240232 474036 240284 474088
rect 3608 473968 3660 474020
rect 353300 473968 353352 474020
rect 273260 471248 273312 471300
rect 292672 471248 292724 471300
rect 277308 469956 277360 470008
rect 290004 469956 290056 470008
rect 270408 469888 270460 469940
rect 280252 469888 280304 469940
rect 271880 469820 271932 469872
rect 289820 469820 289872 469872
rect 267648 468596 267700 468648
rect 274640 468596 274692 468648
rect 275928 468596 275980 468648
rect 287152 468596 287204 468648
rect 266268 468528 266320 468580
rect 273352 468528 273404 468580
rect 274456 468528 274508 468580
rect 285772 468528 285824 468580
rect 217784 468460 217836 468512
rect 254032 468460 254084 468512
rect 267556 468460 267608 468512
rect 277400 468460 277452 468512
rect 278688 468460 278740 468512
rect 291292 468460 291344 468512
rect 262128 467780 262180 467832
rect 269120 467780 269172 467832
rect 264888 467236 264940 467288
rect 271972 467236 272024 467288
rect 274548 467236 274600 467288
rect 284484 467236 284536 467288
rect 263508 467168 263560 467220
rect 270684 467168 270736 467220
rect 271788 467168 271840 467220
rect 281632 467168 281684 467220
rect 269028 467100 269080 467152
rect 278872 467100 278924 467152
rect 280068 467100 280120 467152
rect 292672 467100 292724 467152
rect 218060 465672 218112 465724
rect 316040 465672 316092 465724
rect 3332 462340 3384 462392
rect 333980 462340 334032 462392
rect 274732 456152 274784 456204
rect 295340 456152 295392 456204
rect 217600 456084 217652 456136
rect 233240 456084 233292 456136
rect 276296 456084 276348 456136
rect 298100 456084 298152 456136
rect 217508 456016 217560 456068
rect 233332 456016 233384 456068
rect 277768 456016 277820 456068
rect 300860 456016 300912 456068
rect 336832 454860 336884 454912
rect 361028 454860 361080 454912
rect 219256 454792 219308 454844
rect 244280 454792 244332 454844
rect 270592 454792 270644 454844
rect 287244 454792 287296 454844
rect 302424 454792 302476 454844
rect 580264 454792 580316 454844
rect 219348 454724 219400 454776
rect 247132 454724 247184 454776
rect 267096 454724 267148 454776
rect 283012 454724 283064 454776
rect 300216 454724 300268 454776
rect 580356 454724 580408 454776
rect 217876 454656 217928 454708
rect 255872 454656 255924 454708
rect 268568 454656 268620 454708
rect 285864 454656 285916 454708
rect 298100 454656 298152 454708
rect 580540 454656 580592 454708
rect 84844 453704 84896 453756
rect 330208 453704 330260 453756
rect 320272 453636 320324 453688
rect 358268 453636 358320 453688
rect 329932 453568 329984 453620
rect 362224 453568 362276 453620
rect 32404 453500 32456 453552
rect 327080 453500 327132 453552
rect 327172 453500 327224 453552
rect 361120 453500 361172 453552
rect 10324 453432 10376 453484
rect 351920 453432 351972 453484
rect 4896 453364 4948 453416
rect 352012 453364 352064 453416
rect 5080 453296 5132 453348
rect 353392 453296 353444 453348
rect 322940 452208 322992 452260
rect 358176 452208 358228 452260
rect 307944 452140 307996 452192
rect 360936 452140 360988 452192
rect 310520 452072 310572 452124
rect 364340 452072 364392 452124
rect 71780 452004 71832 452056
rect 347872 452004 347924 452056
rect 10416 451936 10468 451988
rect 331220 451936 331272 451988
rect 6920 451868 6972 451920
rect 350632 451868 350684 451920
rect 303620 450848 303672 450900
rect 360844 450848 360896 450900
rect 301320 450780 301372 450832
rect 359464 450780 359516 450832
rect 305920 450712 305972 450764
rect 494060 450712 494112 450764
rect 8944 450644 8996 450696
rect 329104 450644 329156 450696
rect 4804 450576 4856 450628
rect 324504 450576 324556 450628
rect 4988 450508 5040 450560
rect 326804 450508 326856 450560
rect 299020 449420 299072 449472
rect 358084 449420 358136 449472
rect 296720 449352 296772 449404
rect 371884 449352 371936 449404
rect 169760 449284 169812 449336
rect 317512 449284 317564 449336
rect 106924 449216 106976 449268
rect 319812 449216 319864 449268
rect 3424 449148 3476 449200
rect 325792 449148 325844 449200
rect 332140 449148 332192 449200
rect 527180 449148 527232 449200
rect 3148 448536 3200 448588
rect 233148 448536 233200 448588
rect 309784 448196 309836 448248
rect 412640 448196 412692 448248
rect 153200 448128 153252 448180
rect 319076 448128 319128 448180
rect 307484 448060 307536 448112
rect 477500 448060 477552 448112
rect 88340 447992 88392 448044
rect 321376 447992 321428 448044
rect 305184 447924 305236 447976
rect 542360 447924 542412 447976
rect 23480 447856 23532 447908
rect 323676 447856 323728 447908
rect 3516 447788 3568 447840
rect 332968 447788 333020 447840
rect 233148 446700 233200 446752
rect 233240 446632 233292 446684
rect 233884 446632 233936 446684
rect 234620 446632 234672 446684
rect 235540 446632 235592 446684
rect 248420 446700 248472 446752
rect 249340 446700 249392 446752
rect 251180 446700 251232 446752
rect 251732 446700 251784 446752
rect 252560 446700 252612 446752
rect 253204 446700 253256 446752
rect 253940 446700 253992 446752
rect 254676 446700 254728 446752
rect 258080 446700 258132 446752
rect 258540 446700 258592 446752
rect 274640 446700 274692 446752
rect 275652 446700 275704 446752
rect 278780 446700 278832 446752
rect 279516 446700 279568 446752
rect 281540 446700 281592 446752
rect 282460 446700 282512 446752
rect 289912 446700 289964 446752
rect 290188 446700 290240 446752
rect 291200 446700 291252 446752
rect 291844 446700 291896 446752
rect 292580 446700 292632 446752
rect 293316 446700 293368 446752
rect 327080 446700 327132 446752
rect 327908 446700 327960 446752
rect 351920 446700 351972 446752
rect 352748 446700 352800 446752
rect 353300 446700 353352 446752
rect 354220 446700 354272 446752
rect 355324 446632 355376 446684
rect 238760 446564 238812 446616
rect 239404 446564 239456 446616
rect 334440 446564 334492 446616
rect 462320 446564 462372 446616
rect 201500 446496 201552 446548
rect 343732 446496 343784 446548
rect 136640 446428 136692 446480
rect 346032 446428 346084 446480
rect 40040 446360 40092 446412
rect 322112 446360 322164 446412
rect 325240 446360 325292 446412
rect 580448 446360 580500 446412
rect 255964 445680 256016 445732
rect 260104 445680 260156 445732
rect 262036 445680 262088 445732
rect 262864 445680 262916 445732
rect 266636 445680 266688 445732
rect 260472 445612 260524 445664
rect 265624 445612 265676 445664
rect 268200 445680 268252 445732
rect 313648 445476 313700 445528
rect 340972 445476 341024 445528
rect 178776 445408 178828 445460
rect 349160 445408 349212 445460
rect 7564 445340 7616 445392
rect 351460 445340 351512 445392
rect 261484 445272 261536 445324
rect 265072 445272 265124 445324
rect 341432 445272 341484 445324
rect 358820 445272 358872 445324
rect 252468 445204 252520 445256
rect 257436 445204 257488 445256
rect 339132 445204 339184 445256
rect 359004 445204 359056 445256
rect 314476 445136 314528 445188
rect 357440 445136 357492 445188
rect 257988 445068 258040 445120
rect 263600 445068 263652 445120
rect 312912 445068 312964 445120
rect 358912 445068 358964 445120
rect 217968 445000 218020 445052
rect 315212 445000 315264 445052
rect 318800 445000 318852 445052
rect 356796 445000 356848 445052
rect 244924 444932 244976 444984
rect 246580 444932 246632 444984
rect 315856 444932 315908 444984
rect 358360 444932 358412 444984
rect 304172 444864 304224 444916
rect 359924 444864 359976 444916
rect 232412 444796 232464 444848
rect 337568 444796 337620 444848
rect 231216 444728 231268 444780
rect 339868 444728 339920 444780
rect 247040 444660 247092 444712
rect 360660 444660 360712 444712
rect 232228 444592 232280 444644
rect 346860 444592 346912 444644
rect 209044 444524 209096 444576
rect 349896 444524 349948 444576
rect 309048 444456 309100 444508
rect 321560 444456 321612 444508
rect 349804 444456 349856 444508
rect 359188 444456 359240 444508
rect 340880 444388 340932 444440
rect 357624 444388 357676 444440
rect 342260 443776 342312 443828
rect 581000 443776 581052 443828
rect 340972 443708 341024 443760
rect 580632 443708 580684 443760
rect 3424 443640 3476 443692
rect 247040 443640 247092 443692
rect 321560 443640 321612 443692
rect 580540 443640 580592 443692
rect 325976 443572 326028 443624
rect 336004 443572 336056 443624
rect 231124 443504 231176 443556
rect 342168 443504 342220 443556
rect 231308 443436 231360 443488
rect 356060 443436 356112 443488
rect 174544 443368 174596 443420
rect 342996 443368 343048 443420
rect 84844 443300 84896 443352
rect 340696 443300 340748 443352
rect 302148 443232 302200 443284
rect 580356 443232 580408 443284
rect 297456 443164 297508 443216
rect 580264 443164 580316 443216
rect 32404 443096 32456 443148
rect 338304 443096 338356 443148
rect 8944 443028 8996 443080
rect 325976 443028 326028 443080
rect 4896 442960 4948 443012
rect 344468 442960 344520 443012
rect 3516 442484 3568 442536
rect 304172 442484 304224 442536
rect 3792 442416 3844 442468
rect 315856 442484 315908 442536
rect 3976 442348 4028 442400
rect 318800 442416 318852 442468
rect 3884 442280 3936 442332
rect 311532 442280 311584 442332
rect 311716 442280 311768 442332
rect 3608 442212 3660 442264
rect 312084 442212 312136 442264
rect 316040 442212 316092 442264
rect 304448 442076 304500 442128
rect 318524 442212 318576 442264
rect 340880 442280 340932 442332
rect 349804 442212 349856 442264
rect 363696 441804 363748 441856
rect 363604 441736 363656 441788
rect 364984 441668 365036 441720
rect 580448 441600 580500 441652
rect 3700 439492 3752 439544
rect 232228 439492 232280 439544
rect 363696 431876 363748 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 8944 423580 8996 423632
rect 3332 411204 3384 411256
rect 232228 411204 232280 411256
rect 2872 398760 2924 398812
rect 231308 398760 231360 398812
rect 363604 379448 363656 379500
rect 579620 379448 579672 379500
rect 2872 372512 2924 372564
rect 32404 372512 32456 372564
rect 3332 358708 3384 358760
rect 231216 358708 231268 358760
rect 3332 320084 3384 320136
rect 84844 320084 84896 320136
rect 309416 310496 309468 310548
rect 309784 310496 309836 310548
rect 310796 310496 310848 310548
rect 311164 310496 311216 310548
rect 216128 309068 216180 309120
rect 279976 309068 280028 309120
rect 354956 309068 355008 309120
rect 369216 309068 369268 309120
rect 189724 309000 189776 309052
rect 255780 309000 255832 309052
rect 353116 309000 353168 309052
rect 366456 309000 366508 309052
rect 182824 308932 182876 308984
rect 254400 308932 254452 308984
rect 318800 308932 318852 308984
rect 319168 308932 319220 308984
rect 345388 308932 345440 308984
rect 366548 308932 366600 308984
rect 213552 308864 213604 308916
rect 286876 308864 286928 308916
rect 288900 308864 288952 308916
rect 297272 308864 297324 308916
rect 311992 308864 312044 308916
rect 312360 308864 312412 308916
rect 316132 308864 316184 308916
rect 317052 308864 317104 308916
rect 317420 308864 317472 308916
rect 317788 308864 317840 308916
rect 318984 308864 319036 308916
rect 319536 308864 319588 308916
rect 320180 308864 320232 308916
rect 320640 308864 320692 308916
rect 328460 308864 328512 308916
rect 328828 308864 328880 308916
rect 346308 308864 346360 308916
rect 368756 308864 368808 308916
rect 178684 308796 178736 308848
rect 253020 308796 253072 308848
rect 293960 308796 294012 308848
rect 354772 308796 354824 308848
rect 355416 308796 355468 308848
rect 361304 308796 361356 308848
rect 68284 308728 68336 308780
rect 240692 308728 240744 308780
rect 290740 308728 290792 308780
rect 43444 308660 43496 308712
rect 236368 308660 236420 308712
rect 290924 308660 290976 308712
rect 354680 308660 354732 308712
rect 355416 308660 355468 308712
rect 357256 308660 357308 308712
rect 46204 308592 46256 308644
rect 239312 308592 239364 308644
rect 290280 308592 290332 308644
rect 355692 308592 355744 308644
rect 367468 308592 367520 308644
rect 35164 308524 35216 308576
rect 234528 308524 234580 308576
rect 263692 308524 263744 308576
rect 264888 308524 264940 308576
rect 265072 308524 265124 308576
rect 265532 308524 265584 308576
rect 267832 308524 267884 308576
rect 268844 308524 268896 308576
rect 269120 308524 269172 308576
rect 270224 308524 270276 308576
rect 270500 308524 270552 308576
rect 271512 308524 271564 308576
rect 291384 308524 291436 308576
rect 32404 308456 32456 308508
rect 233148 308456 233200 308508
rect 233332 308456 233384 308508
rect 234252 308456 234304 308508
rect 263600 308456 263652 308508
rect 264060 308456 264112 308508
rect 265348 308456 265400 308508
rect 265900 308456 265952 308508
rect 267740 308456 267792 308508
rect 268200 308456 268252 308508
rect 269212 308456 269264 308508
rect 269672 308456 269724 308508
rect 270684 308456 270736 308508
rect 271604 308456 271656 308508
rect 271972 308456 272024 308508
rect 272984 308456 273036 308508
rect 297272 308524 297324 308576
rect 355324 308524 355376 308576
rect 355784 308524 355836 308576
rect 355968 308524 356020 308576
rect 356796 308524 356848 308576
rect 367560 308524 367612 308576
rect 25504 308388 25556 308440
rect 231768 308388 231820 308440
rect 231952 308388 232004 308440
rect 232872 308388 232924 308440
rect 233516 308388 233568 308440
rect 233884 308388 233936 308440
rect 263876 308388 263928 308440
rect 264428 308388 264480 308440
rect 265256 308388 265308 308440
rect 265808 308388 265860 308440
rect 266544 308388 266596 308440
rect 267188 308388 267240 308440
rect 268016 308388 268068 308440
rect 268568 308388 268620 308440
rect 269304 308388 269356 308440
rect 269764 308388 269816 308440
rect 270592 308388 270644 308440
rect 271052 308388 271104 308440
rect 272156 308388 272208 308440
rect 272524 308388 272576 308440
rect 354680 308456 354732 308508
rect 355600 308456 355652 308508
rect 355876 308456 355928 308508
rect 358084 308456 358136 308508
rect 216220 308320 216272 308372
rect 279332 308320 279384 308372
rect 289176 308320 289228 308372
rect 312084 308320 312136 308372
rect 313096 308320 313148 308372
rect 314660 308320 314712 308372
rect 315396 308320 315448 308372
rect 316132 308320 316184 308372
rect 316776 308320 316828 308372
rect 321560 308320 321612 308372
rect 322480 308320 322532 308372
rect 322940 308320 322992 308372
rect 323860 308320 323912 308372
rect 324320 308320 324372 308372
rect 324596 308320 324648 308372
rect 325792 308320 325844 308372
rect 326804 308320 326856 308372
rect 327080 308320 327132 308372
rect 327448 308320 327500 308372
rect 330116 308320 330168 308372
rect 330484 308320 330536 308372
rect 216312 308252 216364 308304
rect 278596 308252 278648 308304
rect 311992 308252 312044 308304
rect 312728 308252 312780 308304
rect 316040 308252 316092 308304
rect 316408 308252 316460 308304
rect 317512 308252 317564 308304
rect 317880 308252 317932 308304
rect 318892 308252 318944 308304
rect 319260 308252 319312 308304
rect 324412 308252 324464 308304
rect 325332 308252 325384 308304
rect 325700 308252 325752 308304
rect 326620 308252 326672 308304
rect 327264 308252 327316 308304
rect 328184 308252 328236 308304
rect 328552 308252 328604 308304
rect 329196 308252 329248 308304
rect 329840 308252 329892 308304
rect 330300 308252 330352 308304
rect 264980 308184 265032 308236
rect 266268 308184 266320 308236
rect 269488 308184 269540 308236
rect 270132 308184 270184 308236
rect 270868 308184 270920 308236
rect 271144 308184 271196 308236
rect 317696 308184 317748 308236
rect 318248 308184 318300 308236
rect 324596 308184 324648 308236
rect 325240 308184 325292 308236
rect 329932 308184 329984 308236
rect 330944 308184 330996 308236
rect 358268 308388 358320 308440
rect 359648 308388 359700 308440
rect 360200 308388 360252 308440
rect 356336 308320 356388 308372
rect 361028 308388 361080 308440
rect 361580 308388 361632 308440
rect 368848 308388 368900 308440
rect 360384 308320 360436 308372
rect 361120 308320 361172 308372
rect 361304 308320 361356 308372
rect 368940 308320 368992 308372
rect 353576 308252 353628 308304
rect 355784 308184 355836 308236
rect 219072 308116 219124 308168
rect 277952 308116 278004 308168
rect 313280 308116 313332 308168
rect 313648 308116 313700 308168
rect 315028 308116 315080 308168
rect 315856 308116 315908 308168
rect 317052 308116 317104 308168
rect 318064 308116 318116 308168
rect 318892 308116 318944 308168
rect 319812 308116 319864 308168
rect 320456 308116 320508 308168
rect 321100 308116 321152 308168
rect 328736 308116 328788 308168
rect 329564 308116 329616 308168
rect 354036 308116 354088 308168
rect 357532 308252 357584 308304
rect 366272 308252 366324 308304
rect 358084 308184 358136 308236
rect 367836 308184 367888 308236
rect 231768 308048 231820 308100
rect 236092 308048 236144 308100
rect 313556 308048 313608 308100
rect 314476 308048 314528 308100
rect 354772 308048 354824 308100
rect 355508 308048 355560 308100
rect 366180 308116 366232 308168
rect 366364 308048 366416 308100
rect 233148 307980 233200 308032
rect 237932 307980 237984 308032
rect 314752 307980 314804 308032
rect 315120 307980 315172 308032
rect 325884 307980 325936 308032
rect 326252 307980 326304 308032
rect 354496 307980 354548 308032
rect 365076 307980 365128 308032
rect 322296 307912 322348 307964
rect 323584 307912 323636 307964
rect 327080 307912 327132 307964
rect 327816 307912 327868 307964
rect 352656 307912 352708 307964
rect 357532 307912 357584 307964
rect 360568 307912 360620 307964
rect 361212 307912 361264 307964
rect 253204 307844 253256 307896
rect 258080 307844 258132 307896
rect 360292 307844 360344 307896
rect 360660 307844 360712 307896
rect 254768 307776 254820 307828
rect 258724 307776 258776 307828
rect 260656 307776 260708 307828
rect 263508 307776 263560 307828
rect 361672 307776 361724 307828
rect 361948 307776 362000 307828
rect 314660 307708 314712 307760
rect 315488 307708 315540 307760
rect 361856 307708 361908 307760
rect 362500 307708 362552 307760
rect 317512 307504 317564 307556
rect 318616 307504 318668 307556
rect 313280 307368 313332 307420
rect 314108 307368 314160 307420
rect 312360 307232 312412 307284
rect 377404 307232 377456 307284
rect 207020 307164 207072 307216
rect 272432 307164 272484 307216
rect 314016 307164 314068 307216
rect 422300 307164 422352 307216
rect 178040 307096 178092 307148
rect 267004 307096 267056 307148
rect 326160 307096 326212 307148
rect 484400 307096 484452 307148
rect 67640 307028 67692 307080
rect 245476 307028 245528 307080
rect 330760 307028 330812 307080
rect 507860 307028 507912 307080
rect 235172 306824 235224 306876
rect 307760 306824 307812 306876
rect 307944 306824 307996 306876
rect 235080 306620 235132 306672
rect 248604 306688 248656 306740
rect 285956 306688 286008 306740
rect 336924 306688 336976 306740
rect 249708 306620 249760 306672
rect 250260 306620 250312 306672
rect 249892 306552 249944 306604
rect 250352 306552 250404 306604
rect 297180 306552 297232 306604
rect 303804 306552 303856 306604
rect 304172 306552 304224 306604
rect 306380 306552 306432 306604
rect 306932 306552 306984 306604
rect 320364 306552 320416 306604
rect 320732 306552 320784 306604
rect 248604 306484 248656 306536
rect 285956 306484 286008 306536
rect 287152 306484 287204 306536
rect 287520 306484 287572 306536
rect 236092 306416 236144 306468
rect 237104 306416 237156 306468
rect 243268 306416 243320 306468
rect 243452 306416 243504 306468
rect 247224 306416 247276 306468
rect 247960 306416 248012 306468
rect 259552 306416 259604 306468
rect 260196 306416 260248 306468
rect 285680 306416 285732 306468
rect 286232 306416 286284 306468
rect 236276 306348 236328 306400
rect 237012 306348 237064 306400
rect 237748 306348 237800 306400
rect 238484 306348 238536 306400
rect 239128 306348 239180 306400
rect 239956 306348 240008 306400
rect 243084 306348 243136 306400
rect 244096 306348 244148 306400
rect 247132 306348 247184 306400
rect 247592 306348 247644 306400
rect 248512 306348 248564 306400
rect 248696 306348 248748 306400
rect 251180 306348 251232 306400
rect 252192 306348 252244 306400
rect 252744 306348 252796 306400
rect 253480 306348 253532 306400
rect 254216 306348 254268 306400
rect 254676 306348 254728 306400
rect 255688 306348 255740 306400
rect 256424 306348 256476 306400
rect 262404 306348 262456 306400
rect 263048 306348 263100 306400
rect 271696 306348 271748 306400
rect 276756 306348 276808 306400
rect 284300 306348 284352 306400
rect 285220 306348 285272 306400
rect 293960 306348 294012 306400
rect 294696 306348 294748 306400
rect 3332 306280 3384 306332
rect 231124 306280 231176 306332
rect 234896 306280 234948 306332
rect 235724 306280 235776 306332
rect 236184 306280 236236 306332
rect 236644 306280 236696 306332
rect 237656 306280 237708 306332
rect 238392 306280 238444 306332
rect 238944 306280 238996 306332
rect 239404 306280 239456 306332
rect 240416 306280 240468 306332
rect 240876 306280 240928 306332
rect 242992 306280 243044 306332
rect 243636 306280 243688 306332
rect 244372 306280 244424 306332
rect 244740 306280 244792 306332
rect 245660 306280 245712 306332
rect 246396 306280 246448 306332
rect 247408 306280 247460 306332
rect 248052 306280 248104 306332
rect 248420 306280 248472 306332
rect 249432 306280 249484 306332
rect 251364 306280 251416 306332
rect 251732 306280 251784 306332
rect 252928 306280 252980 306332
rect 253572 306280 253624 306332
rect 254308 306280 254360 306332
rect 255044 306280 255096 306332
rect 255596 306280 255648 306332
rect 256056 306280 256108 306332
rect 258356 306280 258408 306332
rect 259184 306280 259236 306332
rect 262496 306280 262548 306332
rect 263140 306280 263192 306332
rect 218888 306212 218940 306264
rect 281356 306280 281408 306332
rect 284392 306280 284444 306332
rect 284760 306280 284812 306332
rect 287244 306280 287296 306332
rect 287980 306280 288032 306332
rect 288440 306280 288492 306332
rect 289360 306280 289412 306332
rect 289820 306280 289872 306332
rect 290464 306280 290516 306332
rect 294144 306280 294196 306332
rect 294604 306280 294656 306332
rect 285772 306212 285824 306264
rect 286140 306212 286192 306264
rect 287336 306212 287388 306264
rect 287612 306212 287664 306264
rect 291200 306212 291252 306264
rect 292304 306212 292356 306264
rect 292764 306212 292816 306264
rect 293224 306212 293276 306264
rect 295340 306212 295392 306264
rect 295800 306212 295852 306264
rect 296720 306212 296772 306264
rect 357716 306552 357768 306604
rect 358084 306552 358136 306604
rect 358912 306484 358964 306536
rect 359280 306484 359332 306536
rect 299480 306416 299532 306468
rect 299848 306416 299900 306468
rect 336924 306416 336976 306468
rect 359096 306416 359148 306468
rect 359464 306416 359516 306468
rect 298192 306348 298244 306400
rect 299388 306348 299440 306400
rect 306656 306348 306708 306400
rect 307484 306348 307536 306400
rect 334164 306348 334216 306400
rect 334900 306348 334952 306400
rect 335452 306348 335504 306400
rect 335728 306348 335780 306400
rect 336832 306348 336884 306400
rect 338028 306348 338080 306400
rect 342260 306348 342312 306400
rect 342812 306348 342864 306400
rect 358728 306348 358780 306400
rect 298100 306280 298152 306332
rect 299020 306280 299072 306332
rect 299572 306280 299624 306332
rect 300768 306280 300820 306332
rect 300952 306280 301004 306332
rect 301320 306280 301372 306332
rect 303620 306280 303672 306332
rect 304540 306280 304592 306332
rect 306472 306280 306524 306332
rect 306748 306280 306800 306332
rect 309232 306280 309284 306332
rect 310152 306280 310204 306332
rect 310612 306280 310664 306332
rect 311532 306280 311584 306332
rect 331588 306280 331640 306332
rect 332324 306280 332376 306332
rect 332784 306280 332836 306332
rect 333244 306280 333296 306332
rect 334072 306280 334124 306332
rect 334808 306280 334860 306332
rect 335360 306280 335412 306332
rect 336280 306280 336332 306332
rect 337016 306280 337068 306332
rect 337568 306280 337620 306332
rect 338212 306280 338264 306332
rect 338948 306280 339000 306332
rect 339500 306280 339552 306332
rect 340328 306280 340380 306332
rect 340972 306280 341024 306332
rect 341524 306280 341576 306332
rect 342444 306280 342496 306332
rect 342904 306280 342956 306332
rect 347780 306280 347832 306332
rect 348608 306280 348660 306332
rect 354864 306280 354916 306332
rect 298284 306212 298336 306264
rect 298560 306212 298612 306264
rect 301044 306212 301096 306264
rect 301228 306212 301280 306264
rect 302516 306212 302568 306264
rect 303160 306212 303212 306264
rect 305000 306212 305052 306264
rect 305368 306212 305420 306264
rect 341156 306212 341208 306264
rect 341892 306212 341944 306264
rect 353392 306212 353444 306264
rect 358728 306212 358780 306264
rect 370136 306280 370188 306332
rect 371700 306212 371752 306264
rect 214564 306144 214616 306196
rect 271696 306144 271748 306196
rect 287428 306144 287480 306196
rect 288072 306144 288124 306196
rect 292580 306144 292632 306196
rect 293040 306144 293092 306196
rect 296904 306144 296956 306196
rect 297824 306144 297876 306196
rect 302424 306144 302476 306196
rect 303068 306144 303120 306196
rect 306472 306144 306524 306196
rect 307392 306144 307444 306196
rect 331404 306144 331456 306196
rect 331956 306144 332008 306196
rect 332600 306144 332652 306196
rect 333704 306144 333756 306196
rect 338396 306144 338448 306196
rect 339040 306144 339092 306196
rect 339776 306144 339828 306196
rect 340420 306144 340472 306196
rect 341248 306144 341300 306196
rect 341984 306144 342036 306196
rect 353852 306144 353904 306196
rect 216588 306076 216640 306128
rect 278872 306076 278924 306128
rect 284484 306076 284536 306128
rect 284852 306076 284904 306128
rect 292672 306076 292724 306128
rect 293684 306076 293736 306128
rect 296812 306076 296864 306128
rect 298008 306076 298060 306128
rect 299664 306076 299716 306128
rect 299940 306076 299992 306128
rect 301044 306076 301096 306128
rect 302148 306076 302200 306128
rect 303896 306076 303948 306128
rect 304908 306076 304960 306128
rect 305000 306076 305052 306128
rect 306104 306076 306156 306128
rect 331220 306076 331272 306128
rect 331680 306076 331732 306128
rect 350356 306076 350408 306128
rect 358636 306076 358688 306128
rect 371516 306144 371568 306196
rect 360108 306076 360160 306128
rect 367744 306076 367796 306128
rect 214840 306008 214892 306060
rect 278136 306008 278188 306060
rect 352196 306008 352248 306060
rect 215208 305940 215260 305992
rect 279516 305940 279568 305992
rect 299664 305940 299716 305992
rect 300400 305940 300452 305992
rect 331220 305940 331272 305992
rect 331864 305940 331916 305992
rect 335728 305940 335780 305992
rect 336648 305940 336700 305992
rect 359924 306008 359976 306060
rect 371332 306008 371384 306060
rect 371424 305940 371476 305992
rect 215944 305872 215996 305924
rect 280252 305872 280304 305924
rect 348976 305872 349028 305924
rect 367652 305872 367704 305924
rect 212448 305804 212500 305856
rect 282276 305804 282328 305856
rect 335544 305804 335596 305856
rect 336188 305804 336240 305856
rect 349712 305804 349764 305856
rect 369124 305804 369176 305856
rect 217876 305736 217928 305788
rect 287152 305736 287204 305788
rect 294052 305736 294104 305788
rect 295064 305736 295116 305788
rect 357716 305736 357768 305788
rect 358360 305736 358412 305788
rect 358452 305736 358504 305788
rect 370412 305736 370464 305788
rect 212356 305668 212408 305720
rect 281632 305668 281684 305720
rect 352932 305668 352984 305720
rect 359924 305668 359976 305720
rect 360016 305668 360068 305720
rect 371608 305668 371660 305720
rect 217692 305600 217744 305652
rect 344468 305600 344520 305652
rect 345572 305600 345624 305652
rect 370228 305600 370280 305652
rect 214932 305532 214984 305584
rect 276112 305532 276164 305584
rect 354312 305532 354364 305584
rect 370044 305532 370096 305584
rect 215116 305464 215168 305516
rect 276296 305464 276348 305516
rect 347228 305464 347280 305516
rect 362408 305464 362460 305516
rect 215024 305396 215076 305448
rect 275468 305396 275520 305448
rect 355232 305396 355284 305448
rect 365168 305396 365220 305448
rect 234712 305328 234764 305380
rect 235632 305328 235684 305380
rect 240232 305328 240284 305380
rect 241336 305328 241388 305380
rect 241796 305328 241848 305380
rect 242348 305328 242400 305380
rect 244556 305328 244608 305380
rect 245108 305328 245160 305380
rect 245936 305328 245988 305380
rect 246488 305328 246540 305380
rect 248696 305328 248748 305380
rect 248972 305328 249024 305380
rect 249800 305328 249852 305380
rect 250260 305328 250312 305380
rect 251456 305328 251508 305380
rect 252100 305328 252152 305380
rect 256700 305328 256752 305380
rect 257436 305328 257488 305380
rect 258264 305328 258316 305380
rect 258816 305328 258868 305380
rect 259460 305328 259512 305380
rect 260104 305328 260156 305380
rect 260840 305328 260892 305380
rect 261024 305328 261076 305380
rect 261208 305328 261260 305380
rect 262128 305328 262180 305380
rect 307944 305328 307996 305380
rect 308864 305328 308916 305380
rect 342352 305328 342404 305380
rect 343364 305328 343416 305380
rect 351736 305328 351788 305380
rect 358452 305328 358504 305380
rect 359280 305328 359332 305380
rect 359832 305328 359884 305380
rect 244372 305260 244424 305312
rect 245016 305260 245068 305312
rect 351092 305260 351144 305312
rect 360016 305260 360068 305312
rect 260840 305192 260892 305244
rect 261668 305192 261720 305244
rect 357808 305192 357860 305244
rect 358544 305192 358596 305244
rect 357440 305124 357492 305176
rect 357992 305124 358044 305176
rect 241520 305056 241572 305108
rect 242256 305056 242308 305108
rect 295524 304920 295576 304972
rect 296444 304920 296496 304972
rect 300860 304920 300912 304972
rect 301688 304920 301740 304972
rect 309968 304444 310020 304496
rect 400220 304444 400272 304496
rect 311164 304376 311216 304428
rect 404360 304376 404412 304428
rect 297088 304308 297140 304360
rect 297364 304308 297416 304360
rect 315120 304308 315172 304360
rect 425060 304308 425112 304360
rect 217508 304240 217560 304292
rect 351552 304240 351604 304292
rect 332968 304172 333020 304224
rect 333336 304172 333388 304224
rect 261116 303968 261168 304020
rect 261484 303968 261536 304020
rect 256792 303696 256844 303748
rect 257160 303696 257212 303748
rect 273444 303696 273496 303748
rect 274364 303696 274416 303748
rect 343640 303696 343692 303748
rect 344652 303696 344704 303748
rect 213828 303560 213880 303612
rect 279792 303560 279844 303612
rect 291292 303560 291344 303612
rect 291476 303560 291528 303612
rect 352472 303560 352524 303612
rect 371792 303560 371844 303612
rect 214472 303492 214524 303544
rect 282092 303492 282144 303544
rect 348516 303492 348568 303544
rect 367928 303492 367980 303544
rect 216036 303424 216088 303476
rect 283380 303424 283432 303476
rect 291476 303424 291528 303476
rect 291936 303424 291988 303476
rect 352012 303424 352064 303476
rect 373080 303424 373132 303476
rect 213736 303356 213788 303408
rect 282736 303356 282788 303408
rect 351276 303356 351328 303408
rect 372712 303356 372764 303408
rect 213184 303288 213236 303340
rect 282552 303288 282604 303340
rect 337108 303288 337160 303340
rect 337660 303288 337712 303340
rect 347688 303288 347740 303340
rect 369308 303288 369360 303340
rect 213368 303220 213420 303272
rect 283012 303220 283064 303272
rect 349896 303220 349948 303272
rect 372804 303220 372856 303272
rect 211712 303152 211764 303204
rect 281816 303152 281868 303204
rect 295616 303152 295668 303204
rect 295984 303152 296036 303204
rect 305184 303152 305236 303204
rect 306012 303152 306064 303204
rect 349252 303152 349304 303204
rect 373172 303152 373224 303204
rect 214656 303084 214708 303136
rect 287060 303084 287112 303136
rect 346492 303084 346544 303136
rect 370504 303084 370556 303136
rect 211988 303016 212040 303068
rect 345848 303016 345900 303068
rect 347412 303016 347464 303068
rect 370688 303016 370740 303068
rect 256976 302948 257028 303000
rect 257344 302948 257396 303000
rect 350632 302948 350684 303000
rect 372896 302948 372948 303000
rect 213092 302880 213144 302932
rect 346768 302880 346820 302932
rect 348332 302880 348384 302932
rect 372988 302880 373040 302932
rect 217968 302812 218020 302864
rect 283656 302812 283708 302864
rect 356060 302812 356112 302864
rect 371884 302812 371936 302864
rect 215852 302744 215904 302796
rect 280436 302744 280488 302796
rect 307852 302744 307904 302796
rect 308772 302744 308824 302796
rect 355968 302744 356020 302796
rect 370320 302744 370372 302796
rect 218980 302676 219032 302728
rect 281172 302676 281224 302728
rect 356980 302676 357032 302728
rect 370596 302676 370648 302728
rect 217416 302608 217468 302660
rect 350816 302608 350868 302660
rect 359004 302608 359056 302660
rect 359740 302608 359792 302660
rect 234988 302200 235040 302252
rect 235264 302200 235316 302252
rect 306748 301656 306800 301708
rect 382280 301656 382332 301708
rect 317880 301588 317932 301640
rect 440240 301588 440292 301640
rect 340788 301520 340840 301572
rect 560300 301520 560352 301572
rect 341432 301452 341484 301504
rect 564440 301452 564492 301504
rect 213276 300772 213328 300824
rect 283932 300772 283984 300824
rect 215760 300704 215812 300756
rect 285864 300704 285916 300756
rect 216404 300636 216456 300688
rect 287520 300636 287572 300688
rect 213460 300568 213512 300620
rect 284300 300568 284352 300620
rect 214380 300500 214432 300552
rect 286140 300500 286192 300552
rect 305368 300500 305420 300552
rect 375380 300500 375432 300552
rect 217048 300432 217100 300484
rect 349252 300432 349304 300484
rect 210792 300364 210844 300416
rect 346952 300364 347004 300416
rect 210700 300296 210752 300348
rect 349160 300296 349212 300348
rect 212172 300228 212224 300280
rect 284392 300228 284444 300280
rect 337200 300228 337252 300280
rect 542360 300228 542412 300280
rect 211068 300160 211120 300212
rect 284484 300160 284536 300212
rect 339408 300160 339460 300212
rect 553400 300160 553452 300212
rect 209688 300092 209740 300144
rect 284668 300092 284720 300144
rect 339868 300092 339920 300144
rect 556160 300092 556212 300144
rect 216496 300024 216548 300076
rect 285956 300024 286008 300076
rect 219348 299956 219400 300008
rect 287244 299956 287296 300008
rect 217784 299888 217836 299940
rect 285312 299888 285364 299940
rect 304448 298936 304500 298988
rect 372620 298936 372672 298988
rect 335268 298868 335320 298920
rect 531320 298868 531372 298920
rect 335820 298800 335872 298852
rect 535460 298800 535512 298852
rect 335728 298732 335780 298784
rect 539600 298732 539652 298784
rect 323584 297576 323636 297628
rect 465080 297576 465132 297628
rect 330116 297508 330168 297560
rect 506480 297508 506532 297560
rect 331680 297440 331732 297492
rect 510620 297440 510672 297492
rect 333888 297372 333940 297424
rect 524420 297372 524472 297424
rect 217600 296284 217652 296336
rect 343640 296284 343692 296336
rect 218704 296216 218756 296268
rect 347872 296216 347924 296268
rect 327540 296148 327592 296200
rect 492680 296148 492732 296200
rect 328920 296080 328972 296132
rect 499580 296080 499632 296132
rect 330024 296012 330076 296064
rect 503720 296012 503772 296064
rect 341248 295944 341300 295996
rect 567200 295944 567252 295996
rect 325976 294788 326028 294840
rect 481640 294788 481692 294840
rect 325884 294720 325936 294772
rect 485780 294720 485832 294772
rect 327448 294652 327500 294704
rect 489920 294652 489972 294704
rect 124220 294584 124272 294636
rect 255688 294584 255740 294636
rect 338488 294584 338540 294636
rect 549260 294584 549312 294636
rect 321928 293428 321980 293480
rect 466460 293428 466512 293480
rect 117320 293360 117372 293412
rect 254308 293360 254360 293412
rect 323308 293360 323360 293412
rect 473360 293360 473412 293412
rect 110420 293292 110472 293344
rect 252928 293292 252980 293344
rect 324688 293292 324740 293344
rect 477500 293292 477552 293344
rect 102140 293224 102192 293276
rect 251180 293224 251232 293276
rect 328828 293224 328880 293276
rect 496820 293224 496872 293276
rect 315028 292000 315080 292052
rect 431960 292000 432012 292052
rect 95240 291932 95292 291984
rect 250168 291932 250220 291984
rect 320640 291932 320692 291984
rect 459560 291932 459612 291984
rect 92480 291864 92532 291916
rect 249800 291864 249852 291916
rect 321836 291864 321888 291916
rect 463700 291864 463752 291916
rect 88340 291796 88392 291848
rect 248420 291796 248472 291848
rect 323216 291796 323268 291848
rect 470600 291796 470652 291848
rect 106924 290640 106976 290692
rect 248788 290640 248840 290692
rect 312176 290640 312228 290692
rect 414020 290640 414072 290692
rect 81440 290572 81492 290624
rect 247408 290572 247460 290624
rect 313556 290572 313608 290624
rect 423680 290572 423732 290624
rect 77300 290504 77352 290556
rect 247500 290504 247552 290556
rect 314936 290504 314988 290556
rect 427820 290504 427872 290556
rect 74540 290436 74592 290488
rect 246120 290436 246172 290488
rect 316408 290436 316460 290488
rect 438860 290436 438912 290488
rect 122840 289280 122892 289332
rect 255596 289280 255648 289332
rect 309416 289280 309468 289332
rect 402980 289280 403032 289332
rect 118700 289212 118752 289264
rect 255504 289212 255556 289264
rect 310704 289212 310756 289264
rect 407212 289212 407264 289264
rect 115940 289144 115992 289196
rect 254216 289144 254268 289196
rect 310796 289144 310848 289196
rect 409880 289144 409932 289196
rect 70400 289076 70452 289128
rect 246028 289076 246080 289128
rect 313464 289076 313516 289128
rect 420920 289076 420972 289128
rect 111800 287920 111852 287972
rect 254124 287920 254176 287972
rect 109040 287852 109092 287904
rect 252744 287852 252796 287904
rect 308036 287852 308088 287904
rect 391940 287852 391992 287904
rect 104900 287784 104952 287836
rect 252836 287784 252888 287836
rect 307944 287784 307996 287836
rect 396080 287784 396132 287836
rect 63500 287716 63552 287768
rect 244648 287716 244700 287768
rect 309324 287716 309376 287768
rect 398840 287716 398892 287768
rect 38660 287648 38712 287700
rect 239128 287648 239180 287700
rect 312084 287648 312136 287700
rect 416780 287648 416832 287700
rect 102232 286492 102284 286544
rect 251456 286492 251508 286544
rect 303896 286492 303948 286544
rect 374000 286492 374052 286544
rect 98000 286424 98052 286476
rect 251548 286424 251600 286476
rect 305276 286424 305328 286476
rect 378140 286424 378192 286476
rect 93860 286356 93912 286408
rect 250076 286356 250128 286408
rect 306656 286356 306708 286408
rect 389180 286356 389232 286408
rect 54484 286288 54536 286340
rect 241980 286288 242032 286340
rect 343916 286288 343968 286340
rect 576860 286288 576912 286340
rect 118792 285200 118844 285252
rect 255412 285200 255464 285252
rect 303804 285200 303856 285252
rect 371240 285200 371292 285252
rect 114560 285132 114612 285184
rect 254400 285132 254452 285184
rect 319260 285132 319312 285184
rect 447140 285132 447192 285184
rect 110512 285064 110564 285116
rect 254032 285064 254084 285116
rect 342720 285064 342772 285116
rect 552664 285064 552716 285116
rect 91100 284996 91152 285048
rect 249984 284996 250036 285048
rect 341156 284996 341208 285048
rect 565820 284996 565872 285048
rect 49700 284928 49752 284980
rect 241888 284928 241940 284980
rect 342628 284928 342680 284980
rect 569960 284928 570012 284980
rect 107660 283840 107712 283892
rect 253020 283840 253072 283892
rect 103520 283772 103572 283824
rect 252652 283772 252704 283824
rect 334348 283772 334400 283824
rect 528560 283772 528612 283824
rect 100760 283704 100812 283756
rect 251364 283704 251416 283756
rect 339776 283704 339828 283756
rect 538956 283704 539008 283756
rect 77392 283636 77444 283688
rect 247316 283636 247368 283688
rect 338304 283636 338356 283688
rect 547880 283636 547932 283688
rect 31760 283568 31812 283620
rect 237748 283568 237800 283620
rect 338396 283568 338448 283620
rect 552020 283568 552072 283620
rect 160100 282412 160152 282464
rect 262496 282412 262548 282464
rect 155960 282344 156012 282396
rect 262588 282344 262640 282396
rect 317788 282344 317840 282396
rect 443000 282344 443052 282396
rect 96620 282276 96672 282328
rect 251272 282276 251324 282328
rect 333060 282276 333112 282328
rect 520280 282276 520332 282328
rect 73160 282208 73212 282260
rect 245936 282208 245988 282260
rect 334256 282208 334308 282260
rect 527180 282208 527232 282260
rect 43536 282140 43588 282192
rect 240508 282140 240560 282192
rect 334164 282140 334216 282192
rect 531412 282140 531464 282192
rect 218428 281120 218480 281172
rect 273720 281120 273772 281172
rect 205640 281052 205692 281104
rect 272248 281052 272300 281104
rect 198740 280984 198792 281036
rect 270960 280984 271012 281036
rect 329932 280984 329984 281036
rect 509240 280984 509292 281036
rect 151820 280916 151872 280968
rect 261392 280916 261444 280968
rect 331496 280916 331548 280968
rect 513380 280916 513432 280968
rect 149060 280848 149112 280900
rect 261300 280848 261352 280900
rect 331588 280848 331640 280900
rect 516140 280848 516192 280900
rect 36544 280780 36596 280832
rect 239036 280780 239088 280832
rect 341064 280780 341116 280832
rect 563060 280780 563112 280832
rect 196624 279692 196676 279744
rect 269488 279692 269540 279744
rect 191840 279624 191892 279676
rect 269580 279624 269632 279676
rect 328644 279624 328696 279676
rect 498200 279624 498252 279676
rect 187700 279556 187752 279608
rect 268200 279556 268252 279608
rect 328736 279556 328788 279608
rect 502340 279556 502392 279608
rect 144920 279488 144972 279540
rect 259920 279488 259972 279540
rect 329840 279488 329892 279540
rect 506572 279488 506624 279540
rect 69020 279420 69072 279472
rect 245844 279420 245896 279472
rect 339684 279420 339736 279472
rect 556252 279420 556304 279472
rect 184940 278264 184992 278316
rect 268108 278264 268160 278316
rect 180800 278196 180852 278248
rect 266728 278196 266780 278248
rect 325792 278196 325844 278248
rect 488540 278196 488592 278248
rect 176660 278128 176712 278180
rect 266636 278128 266688 278180
rect 327356 278128 327408 278180
rect 491300 278128 491352 278180
rect 142160 278060 142212 278112
rect 259828 278060 259880 278112
rect 327264 278060 327316 278112
rect 495440 278060 495492 278112
rect 66260 277992 66312 278044
rect 244556 277992 244608 278044
rect 337108 277992 337160 278044
rect 545120 277992 545172 278044
rect 173900 276904 173952 276956
rect 265348 276904 265400 276956
rect 169760 276836 169812 276888
rect 265440 276836 265492 276888
rect 316316 276836 316368 276888
rect 437480 276836 437532 276888
rect 61384 276768 61436 276820
rect 243360 276768 243412 276820
rect 319168 276768 319220 276820
rect 451280 276768 451332 276820
rect 62120 276700 62172 276752
rect 244464 276700 244516 276752
rect 320548 276700 320600 276752
rect 455420 276700 455472 276752
rect 26884 276632 26936 276684
rect 236276 276632 236328 276684
rect 321744 276632 321796 276684
rect 462320 276632 462372 276684
rect 313372 275476 313424 275528
rect 419540 275476 419592 275528
rect 167000 275408 167052 275460
rect 264060 275408 264112 275460
rect 314844 275408 314896 275460
rect 426440 275408 426492 275460
rect 162860 275340 162912 275392
rect 263968 275340 264020 275392
rect 316224 275340 316276 275392
rect 433340 275340 433392 275392
rect 57244 275272 57296 275324
rect 243268 275272 243320 275324
rect 317696 275272 317748 275324
rect 444380 275272 444432 275324
rect 206284 274184 206336 274236
rect 272064 274184 272116 274236
rect 201500 274116 201552 274168
rect 270868 274116 270920 274168
rect 309232 274116 309284 274168
rect 401600 274116 401652 274168
rect 158720 274048 158772 274100
rect 262404 274048 262456 274100
rect 310612 274048 310664 274100
rect 408500 274048 408552 274100
rect 138020 273980 138072 274032
rect 258356 273980 258408 274032
rect 311992 273980 312044 274032
rect 415492 273980 415544 274032
rect 30380 273912 30432 273964
rect 237656 273912 237708 273964
rect 313280 273912 313332 273964
rect 423772 273912 423824 273964
rect 364984 273164 365036 273216
rect 579620 273164 579672 273216
rect 197360 272824 197412 272876
rect 270776 272824 270828 272876
rect 193220 272756 193272 272808
rect 269304 272756 269356 272808
rect 192484 272688 192536 272740
rect 269396 272688 269448 272740
rect 154580 272620 154632 272672
rect 262312 272620 262364 272672
rect 307760 272620 307812 272672
rect 390560 272620 390612 272672
rect 131120 272552 131172 272604
rect 257160 272552 257212 272604
rect 307852 272552 307904 272604
rect 394700 272552 394752 272604
rect 27620 272484 27672 272536
rect 237564 272484 237616 272536
rect 309140 272484 309192 272536
rect 398932 272484 398984 272536
rect 188344 271464 188396 271516
rect 268016 271464 268068 271516
rect 183560 271396 183612 271448
rect 267924 271396 267976 271448
rect 179420 271328 179472 271380
rect 266544 271328 266596 271380
rect 305184 271328 305236 271380
rect 380900 271328 380952 271380
rect 140780 271260 140832 271312
rect 259736 271260 259788 271312
rect 306564 271260 306616 271312
rect 383660 271260 383712 271312
rect 93952 271192 94004 271244
rect 249892 271192 249944 271244
rect 306472 271192 306524 271244
rect 387800 271192 387852 271244
rect 22100 271124 22152 271176
rect 236184 271124 236236 271176
rect 320456 271124 320508 271176
rect 458180 271124 458232 271176
rect 176752 270104 176804 270156
rect 266452 270104 266504 270156
rect 172520 270036 172572 270088
rect 265256 270036 265308 270088
rect 168380 269968 168432 270020
rect 265164 269968 265216 270020
rect 136640 269900 136692 269952
rect 258264 269900 258316 269952
rect 303620 269900 303672 269952
rect 374092 269900 374144 269952
rect 89720 269832 89772 269884
rect 250260 269832 250312 269884
rect 305092 269832 305144 269884
rect 376760 269832 376812 269884
rect 13820 269764 13872 269816
rect 235080 269764 235132 269816
rect 317604 269764 317656 269816
rect 440332 269764 440384 269816
rect 165620 268608 165672 268660
rect 263876 268608 263928 268660
rect 302516 268608 302568 268660
rect 365720 268608 365772 268660
rect 161480 268540 161532 268592
rect 263784 268540 263836 268592
rect 320364 268540 320416 268592
rect 456800 268540 456852 268592
rect 157340 268472 157392 268524
rect 262680 268472 262732 268524
rect 339592 268472 339644 268524
rect 516784 268472 516836 268524
rect 133880 268404 133932 268456
rect 258172 268404 258224 268456
rect 342536 268404 342588 268456
rect 520924 268404 520976 268456
rect 52460 268336 52512 268388
rect 241796 268336 241848 268388
rect 342444 268336 342496 268388
rect 525064 268336 525116 268388
rect 3332 267656 3384 267708
rect 174544 267656 174596 267708
rect 153200 267180 153252 267232
rect 261208 267180 261260 267232
rect 319076 267180 319128 267232
rect 448520 267180 448572 267232
rect 150440 267112 150492 267164
rect 261116 267112 261168 267164
rect 338212 267112 338264 267164
rect 508504 267112 508556 267164
rect 48320 267044 48372 267096
rect 241704 267044 241756 267096
rect 337016 267044 337068 267096
rect 543740 267044 543792 267096
rect 8300 266976 8352 267028
rect 233516 266976 233568 267028
rect 338120 266976 338172 267028
rect 547972 266976 548024 267028
rect 209780 265956 209832 266008
rect 271972 265956 272024 266008
rect 202880 265888 202932 265940
rect 270684 265888 270736 265940
rect 200120 265820 200172 265872
rect 270592 265820 270644 265872
rect 318984 265820 319036 265872
rect 449900 265820 449952 265872
rect 146300 265752 146352 265804
rect 261024 265752 261076 265804
rect 335636 265752 335688 265804
rect 496084 265752 496136 265804
rect 126980 265684 127032 265736
rect 257068 265684 257120 265736
rect 335544 265684 335596 265736
rect 502984 265684 503036 265736
rect 44180 265616 44232 265668
rect 240416 265616 240468 265668
rect 334072 265616 334124 265668
rect 529940 265616 529992 265668
rect 195980 264528 196032 264580
rect 269120 264528 269172 264580
rect 193312 264460 193364 264512
rect 269212 264460 269264 264512
rect 189080 264392 189132 264444
rect 267832 264392 267884 264444
rect 316132 264392 316184 264444
rect 436100 264392 436152 264444
rect 139400 264324 139452 264376
rect 259644 264324 259696 264376
rect 331404 264324 331456 264376
rect 457444 264324 457496 264376
rect 85580 264256 85632 264308
rect 248696 264256 248748 264308
rect 332876 264256 332928 264308
rect 467104 264256 467156 264308
rect 2780 264188 2832 264240
rect 232136 264188 232188 264240
rect 332968 264188 333020 264240
rect 476764 264188 476816 264240
rect 185032 263100 185084 263152
rect 267740 263100 267792 263152
rect 175280 263032 175332 263084
rect 264980 263032 265032 263084
rect 311900 263032 311952 263084
rect 412640 263032 412692 263084
rect 171140 262964 171192 263016
rect 265072 262964 265124 263016
rect 328552 262964 328604 263016
rect 432604 262964 432656 263016
rect 132500 262896 132552 262948
rect 253204 262896 253256 262948
rect 328460 262896 328512 262948
rect 498292 262896 498344 262948
rect 40040 262828 40092 262880
rect 240324 262828 240376 262880
rect 331312 262828 331364 262880
rect 512000 262828 512052 262880
rect 168472 261740 168524 261792
rect 263692 261740 263744 261792
rect 164240 261672 164292 261724
rect 263600 261672 263652 261724
rect 325700 261672 325752 261724
rect 487160 261672 487212 261724
rect 160192 261604 160244 261656
rect 260104 261604 260156 261656
rect 327172 261604 327224 261656
rect 490012 261604 490064 261656
rect 128360 261536 128412 261588
rect 256976 261536 257028 261588
rect 327080 261536 327132 261588
rect 494060 261536 494112 261588
rect 82820 261468 82872 261520
rect 248604 261468 248656 261520
rect 336924 261468 336976 261520
rect 539692 261468 539744 261520
rect 211804 260312 211856 260364
rect 266820 260312 266872 260364
rect 125600 260244 125652 260296
rect 256884 260244 256936 260296
rect 324596 260244 324648 260296
rect 480260 260244 480312 260296
rect 64880 260176 64932 260228
rect 244372 260176 244424 260228
rect 333980 260176 334032 260228
rect 525800 260176 525852 260228
rect 35900 260108 35952 260160
rect 238944 260108 238996 260160
rect 343824 260108 343876 260160
rect 575480 260108 575532 260160
rect 217232 258952 217284 259004
rect 344100 258952 344152 259004
rect 69112 258884 69164 258936
rect 245752 258884 245804 258936
rect 60740 258816 60792 258868
rect 244740 258816 244792 258868
rect 35256 258748 35308 258800
rect 238852 258748 238904 258800
rect 4804 258680 4856 258732
rect 231860 258680 231912 258732
rect 320272 256164 320324 256216
rect 454040 256164 454092 256216
rect 24860 256096 24912 256148
rect 236092 256096 236144 256148
rect 321652 256096 321704 256148
rect 460940 256096 460992 256148
rect 17224 256028 17276 256080
rect 234988 256028 235040 256080
rect 323032 256028 323084 256080
rect 467840 256028 467892 256080
rect 8944 255960 8996 256012
rect 233424 255960 233476 256012
rect 324504 255960 324556 256012
rect 474740 255960 474792 256012
rect 116584 254804 116636 254856
rect 240232 254804 240284 254856
rect 79324 254736 79376 254788
rect 243084 254736 243136 254788
rect 56600 254668 56652 254720
rect 243176 254668 243228 254720
rect 318064 254668 318116 254720
rect 432052 254668 432104 254720
rect 44272 254600 44324 254652
rect 240600 254600 240652 254652
rect 342352 254600 342404 254652
rect 574100 254600 574152 254652
rect 39304 254532 39356 254584
rect 239220 254532 239272 254584
rect 344008 254532 344060 254584
rect 578240 254532 578292 254584
rect 2872 254192 2924 254244
rect 4896 254192 4948 254244
rect 86960 253444 87012 253496
rect 248880 253444 248932 253496
rect 294236 253444 294288 253496
rect 365996 253444 366048 253496
rect 84200 253376 84252 253428
rect 248512 253376 248564 253428
rect 331220 253376 331272 253428
rect 514852 253376 514904 253428
rect 80060 253308 80112 253360
rect 247224 253308 247276 253360
rect 332692 253308 332744 253360
rect 517520 253308 517572 253360
rect 17960 253240 18012 253292
rect 234896 253240 234948 253292
rect 332784 253240 332836 253292
rect 521660 253240 521712 253292
rect 9680 253172 9732 253224
rect 233332 253172 233384 253224
rect 342260 253172 342312 253224
rect 571340 253172 571392 253224
rect 218520 252152 218572 252204
rect 347780 252152 347832 252204
rect 121460 252084 121512 252136
rect 255780 252084 255832 252136
rect 31024 252016 31076 252068
rect 237840 252016 237892 252068
rect 317512 252016 317564 252068
rect 445760 252016 445812 252068
rect 26240 251948 26292 252000
rect 237472 251948 237524 252000
rect 318800 251948 318852 252000
rect 448612 251948 448664 252000
rect 20720 251880 20772 251932
rect 236368 251880 236420 251932
rect 318892 251880 318944 251932
rect 452660 251880 452712 251932
rect 12440 251812 12492 251864
rect 234804 251812 234856 251864
rect 320180 251812 320232 251864
rect 456892 251812 456944 251864
rect 292856 251132 292908 251184
rect 358820 251132 358872 251184
rect 298376 251064 298428 251116
rect 364708 251064 364760 251116
rect 299940 250996 299992 251048
rect 367192 250996 367244 251048
rect 292948 250928 293000 250980
rect 360200 250928 360252 250980
rect 295800 250860 295852 250912
rect 363144 250860 363196 250912
rect 297180 250792 297232 250844
rect 364800 250792 364852 250844
rect 174544 250724 174596 250776
rect 251640 250724 251692 250776
rect 298468 250724 298520 250776
rect 367100 250724 367152 250776
rect 78680 250656 78732 250708
rect 247132 250656 247184 250708
rect 293040 250656 293092 250708
rect 364892 250656 364944 250708
rect 75920 250588 75972 250640
rect 247040 250588 247092 250640
rect 291476 250588 291528 250640
rect 368480 250588 368532 250640
rect 71780 250520 71832 250572
rect 245660 250520 245712 250572
rect 305000 250520 305052 250572
rect 382372 250520 382424 250572
rect 16580 250452 16632 250504
rect 234712 250452 234764 250504
rect 291568 250452 291620 250504
rect 369860 250452 369912 250504
rect 297272 250384 297324 250436
rect 363236 250384 363288 250436
rect 301228 250316 301280 250368
rect 365904 250316 365956 250368
rect 295708 250248 295760 250300
rect 360292 250248 360344 250300
rect 209872 249228 209924 249280
rect 272340 249228 272392 249280
rect 317420 249228 317472 249280
rect 441620 249228 441672 249280
rect 201592 249160 201644 249212
rect 270500 249160 270552 249212
rect 336740 249160 336792 249212
rect 534724 249160 534776 249212
rect 135260 249092 135312 249144
rect 258448 249092 258500 249144
rect 335452 249092 335504 249144
rect 534080 249092 534132 249144
rect 57980 249024 58032 249076
rect 242992 249024 243044 249076
rect 335360 249024 335412 249076
rect 538220 249024 538272 249076
rect 299756 248344 299808 248396
rect 363328 248344 363380 248396
rect 298284 248276 298336 248328
rect 362960 248276 363012 248328
rect 295616 248208 295668 248260
rect 361672 248208 361724 248260
rect 298192 248140 298244 248192
rect 364616 248140 364668 248192
rect 296996 248072 297048 248124
rect 364340 248072 364392 248124
rect 297088 248004 297140 248056
rect 364524 248004 364576 248056
rect 151912 247936 151964 247988
rect 260840 247936 260892 247988
rect 296812 247936 296864 247988
rect 364432 247936 364484 247988
rect 147680 247868 147732 247920
rect 260932 247868 260984 247920
rect 292672 247868 292724 247920
rect 360844 247868 360896 247920
rect 143540 247800 143592 247852
rect 259552 247800 259604 247852
rect 292764 247800 292816 247852
rect 362132 247800 362184 247852
rect 127072 247732 127124 247784
rect 256792 247732 256844 247784
rect 291384 247732 291436 247784
rect 366088 247732 366140 247784
rect 53840 247664 53892 247716
rect 242900 247664 242952 247716
rect 288716 247664 288768 247716
rect 364984 247664 365036 247716
rect 294144 247596 294196 247648
rect 356704 247596 356756 247648
rect 295432 247528 295484 247580
rect 358360 247528 358412 247580
rect 301136 247460 301188 247512
rect 363052 247460 363104 247512
rect 211160 246576 211212 246628
rect 273260 246576 273312 246628
rect 314752 246576 314804 246628
rect 387064 246576 387116 246628
rect 53104 246508 53156 246560
rect 241520 246508 241572 246560
rect 290004 246508 290056 246560
rect 367284 246508 367336 246560
rect 48964 246440 49016 246492
rect 241612 246440 241664 246492
rect 310520 246440 310572 246492
rect 405740 246440 405792 246492
rect 13084 246372 13136 246424
rect 234620 246372 234672 246424
rect 314660 246372 314712 246424
rect 430580 246372 430632 246424
rect 6920 246304 6972 246356
rect 233700 246304 233752 246356
rect 324412 246304 324464 246356
rect 481732 246304 481784 246356
rect 300860 245556 300912 245608
rect 357440 245556 357492 245608
rect 300952 245488 301004 245540
rect 358176 245488 358228 245540
rect 355784 245420 355836 245472
rect 368572 245420 368624 245472
rect 219256 245352 219308 245404
rect 287428 245352 287480 245404
rect 294052 245352 294104 245404
rect 358084 245352 358136 245404
rect 213644 245284 213696 245336
rect 288532 245284 288584 245336
rect 293960 245284 294012 245336
rect 358176 245284 358228 245336
rect 358268 245284 358320 245336
rect 367376 245284 367428 245336
rect 213000 245216 213052 245268
rect 288624 245216 288676 245268
rect 292580 245216 292632 245268
rect 359464 245216 359516 245268
rect 143632 245148 143684 245200
rect 259460 245148 259512 245200
rect 291292 245148 291344 245200
rect 368664 245148 368716 245200
rect 135352 245080 135404 245132
rect 254584 245080 254636 245132
rect 324320 245080 324372 245132
rect 476120 245080 476172 245132
rect 129740 245012 129792 245064
rect 256700 245012 256752 245064
rect 339500 245012 339552 245064
rect 557540 245012 557592 245064
rect 7656 244944 7708 244996
rect 231952 244944 232004 244996
rect 340880 244944 340932 244996
rect 561680 244944 561732 244996
rect 4896 244876 4948 244928
rect 232044 244876 232096 244928
rect 340972 244876 341024 244928
rect 564532 244876 564584 244928
rect 355600 244536 355652 244588
rect 363512 244536 363564 244588
rect 355692 244264 355744 244316
rect 362316 244264 362368 244316
rect 355324 244128 355376 244180
rect 362224 244128 362276 244180
rect 355416 243788 355468 243840
rect 369952 243788 370004 243840
rect 291200 243720 291252 243772
rect 358268 243720 358320 243772
rect 219164 243652 219216 243704
rect 286048 243652 286100 243704
rect 289912 243652 289964 243704
rect 359556 243652 359608 243704
rect 218612 243584 218664 243636
rect 285772 243584 285824 243636
rect 289820 243584 289872 243636
rect 360936 243584 360988 243636
rect 217140 243516 217192 243568
rect 287336 243516 287388 243568
rect 288440 243516 288492 243568
rect 363604 243516 363656 243568
rect 215760 195780 215812 195832
rect 217508 195780 217560 195832
rect 214380 195236 214432 195288
rect 217324 195236 217376 195288
rect 210700 193128 210752 193180
rect 216680 193128 216732 193180
rect 210884 189660 210936 189712
rect 218060 189660 218112 189712
rect 210792 188980 210844 189032
rect 216680 188980 216732 189032
rect 213000 168920 213052 168972
rect 217416 168920 217468 168972
rect 218796 166268 218848 166320
rect 218980 166268 219032 166320
rect 356244 159808 356296 159860
rect 357992 159808 358044 159860
rect 214472 159604 214524 159656
rect 256700 159604 256752 159656
rect 211712 159536 211764 159588
rect 255320 159536 255372 159588
rect 317696 159536 317748 159588
rect 356796 159536 356848 159588
rect 213184 159468 213236 159520
rect 259552 159468 259604 159520
rect 314660 159468 314712 159520
rect 357808 159468 357860 159520
rect 217876 159400 217928 159452
rect 284392 159400 284444 159452
rect 307852 159400 307904 159452
rect 359372 159400 359424 159452
rect 213552 159332 213604 159384
rect 281540 159332 281592 159384
rect 292580 159332 292632 159384
rect 359188 159332 359240 159384
rect 355324 159264 355376 159316
rect 361948 159264 362000 159316
rect 285956 159196 286008 159248
rect 365168 159196 365220 159248
rect 291016 159128 291068 159180
rect 371884 159128 371936 159180
rect 279240 159060 279292 159112
rect 362040 159060 362092 159112
rect 277032 158992 277084 159044
rect 360568 158992 360620 159044
rect 278136 158924 278188 158976
rect 355324 158924 355376 158976
rect 355416 158924 355468 158976
rect 360660 158924 360712 158976
rect 273352 158856 273404 158908
rect 359280 158856 359332 158908
rect 214472 158788 214524 158840
rect 214656 158788 214708 158840
rect 275836 158788 275888 158840
rect 360752 158788 360804 158840
rect 213092 158720 213144 158772
rect 239588 158720 239640 158772
rect 274456 158720 274508 158772
rect 355416 158720 355468 158772
rect 355508 158720 355560 158772
rect 357900 158720 357952 158772
rect 211988 158652 212040 158704
rect 238116 158652 238168 158704
rect 268384 158652 268436 158704
rect 373080 158652 373132 158704
rect 218980 158584 219032 158636
rect 220820 158584 220872 158636
rect 224224 158584 224276 158636
rect 229100 158584 229152 158636
rect 268752 158584 268804 158636
rect 357624 158584 357676 158636
rect 219072 158516 219124 158568
rect 234620 158516 234672 158568
rect 272248 158516 272300 158568
rect 292580 158516 292632 158568
rect 298560 158516 298612 158568
rect 356244 158516 356296 158568
rect 211896 158448 211948 158500
rect 230480 158448 230532 158500
rect 301044 158448 301096 158500
rect 357532 158448 357584 158500
rect 216312 158380 216364 158432
rect 238760 158380 238812 158432
rect 303528 158380 303580 158432
rect 357716 158380 357768 158432
rect 212080 158312 212132 158364
rect 234712 158312 234764 158364
rect 306104 158312 306156 158364
rect 359096 158312 359148 158364
rect 216220 158244 216272 158296
rect 242992 158244 243044 158296
rect 271144 158244 271196 158296
rect 307852 158244 307904 158296
rect 308680 158244 308732 158296
rect 358912 158244 358964 158296
rect 212264 158176 212316 158228
rect 241520 158176 241572 158228
rect 311072 158176 311124 158228
rect 359004 158176 359056 158228
rect 216128 158108 216180 158160
rect 245660 158108 245712 158160
rect 313464 158108 313516 158160
rect 359648 158108 359700 158160
rect 215944 158040 215996 158092
rect 247040 158040 247092 158092
rect 269856 158040 269908 158092
rect 314660 158040 314712 158092
rect 315856 158040 315908 158092
rect 360476 158040 360528 158092
rect 218888 157972 218940 158024
rect 252560 157972 252612 158024
rect 293592 157972 293644 158024
rect 317696 157972 317748 158024
rect 318616 157972 318668 158024
rect 360384 157972 360436 158024
rect 214564 157904 214616 157956
rect 224224 157904 224276 157956
rect 321008 157904 321060 157956
rect 361028 157904 361080 157956
rect 214656 157836 214708 157888
rect 219440 157836 219492 157888
rect 323400 157836 323452 157888
rect 361764 157836 361816 157888
rect 325976 157768 326028 157820
rect 361856 157768 361908 157820
rect 216220 157360 216272 157412
rect 223580 157360 223632 157412
rect 242440 157292 242492 157344
rect 367928 157292 367980 157344
rect 244280 157224 244332 157276
rect 368756 157224 368808 157276
rect 248328 157156 248380 157208
rect 370228 157156 370280 157208
rect 250904 157088 250956 157140
rect 370504 157088 370556 157140
rect 252100 157020 252152 157072
rect 371608 157020 371660 157072
rect 257344 156952 257396 157004
rect 366180 156952 366232 157004
rect 261760 156884 261812 156936
rect 368940 156884 368992 156936
rect 259920 156816 259972 156868
rect 365076 156816 365128 156868
rect 264336 156748 264388 156800
rect 368848 156748 368900 156800
rect 265900 156680 265952 156732
rect 367560 156680 367612 156732
rect 271052 156612 271104 156664
rect 371792 156612 371844 156664
rect 276112 156544 276164 156596
rect 370136 156544 370188 156596
rect 283656 156476 283708 156528
rect 371700 156476 371752 156528
rect 295984 156408 296036 156460
rect 370596 156408 370648 156460
rect 240600 155864 240652 155916
rect 369308 155864 369360 155916
rect 246764 155796 246816 155848
rect 369032 155796 369084 155848
rect 248696 155728 248748 155780
rect 369124 155728 369176 155780
rect 247776 155660 247828 155712
rect 367652 155660 367704 155712
rect 218796 155592 218848 155644
rect 251272 155592 251324 155644
rect 253480 155592 253532 155644
rect 371424 155592 371476 155644
rect 245568 155524 245620 155576
rect 362408 155524 362460 155576
rect 215852 155456 215904 155508
rect 248420 155456 248472 155508
rect 250720 155456 250772 155508
rect 367744 155456 367796 155508
rect 212356 155388 212408 155440
rect 253940 155388 253992 155440
rect 256056 155388 256108 155440
rect 372988 155388 373040 155440
rect 218704 155320 218756 155372
rect 266360 155320 266412 155372
rect 266636 155320 266688 155372
rect 367468 155320 367520 155372
rect 212172 155252 212224 155304
rect 270500 155252 270552 155304
rect 273720 155252 273772 155304
rect 371332 155252 371384 155304
rect 217508 155184 217560 155236
rect 277400 155184 277452 155236
rect 278504 155184 278556 155236
rect 371516 155184 371568 155236
rect 218612 155116 218664 155168
rect 278780 155116 278832 155168
rect 281080 155116 281132 155168
rect 370044 155116 370096 155168
rect 217140 155048 217192 155100
rect 285680 155048 285732 155100
rect 288256 155048 288308 155100
rect 370320 155048 370372 155100
rect 214472 154980 214524 155032
rect 282920 154980 282972 155032
rect 261208 154504 261260 154556
rect 372804 154504 372856 154556
rect 263692 154436 263744 154488
rect 372896 154436 372948 154488
rect 265992 154368 266044 154420
rect 372712 154368 372764 154420
rect 209688 152532 209740 152584
rect 269120 152532 269172 152584
rect 213460 152464 213512 152516
rect 273260 152464 273312 152516
rect 3608 150356 3660 150408
rect 178776 150356 178828 150408
rect 3148 111732 3200 111784
rect 209044 111732 209096 111784
rect 3516 97588 3568 97640
rect 7564 97588 7616 97640
rect 143540 11704 143592 11756
rect 144736 11704 144788 11756
rect 168380 11704 168432 11756
rect 169576 11704 169628 11756
rect 176660 11704 176712 11756
rect 177856 11704 177908 11756
rect 234620 11704 234672 11756
rect 235816 11704 235868 11756
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 307944 9596 307996 9648
rect 369860 9596 369912 9648
rect 306748 9528 306800 9580
rect 368664 9528 368716 9580
rect 305552 9460 305604 9512
rect 367376 9460 367428 9512
rect 304356 9392 304408 9444
rect 366088 9392 366140 9444
rect 299664 9324 299716 9376
rect 362316 9324 362368 9376
rect 297272 9256 297324 9308
rect 359556 9256 359608 9308
rect 301964 9188 302016 9240
rect 369952 9188 370004 9240
rect 298468 9120 298520 9172
rect 367284 9120 367336 9172
rect 296076 9052 296128 9104
rect 364984 9052 365036 9104
rect 294880 8984 294932 9036
rect 363604 8984 363656 9036
rect 293684 8916 293736 8968
rect 368572 8916 368624 8968
rect 300768 8848 300820 8900
rect 360936 8848 360988 8900
rect 303160 8780 303212 8832
rect 363512 8780 363564 8832
rect 316224 8712 316276 8764
rect 364892 8712 364944 8764
rect 323308 6808 323360 6860
rect 358176 6808 358228 6860
rect 317328 6740 317380 6792
rect 360844 6740 360896 6792
rect 320916 6672 320968 6724
rect 365812 6672 365864 6724
rect 318524 6604 318576 6656
rect 363420 6604 363472 6656
rect 313832 6536 313884 6588
rect 359464 6536 359516 6588
rect 315028 6468 315080 6520
rect 362132 6468 362184 6520
rect 312636 6400 312688 6452
rect 360200 6400 360252 6452
rect 311440 6332 311492 6384
rect 358820 6332 358872 6384
rect 310244 6264 310296 6316
rect 358268 6264 358320 6316
rect 309048 6196 309100 6248
rect 368480 6196 368532 6248
rect 292580 6128 292632 6180
rect 362224 6128 362276 6180
rect 326804 6060 326856 6112
rect 360292 6060 360344 6112
rect 330392 5992 330444 6044
rect 363144 5992 363196 6044
rect 333888 5924 333940 5976
rect 364800 5924 364852 5976
rect 2872 4088 2924 4140
rect 7748 4088 7800 4140
rect 15936 4088 15988 4140
rect 17224 4088 17276 4140
rect 24216 4088 24268 4140
rect 26884 4088 26936 4140
rect 213736 4088 213788 4140
rect 260656 4088 260708 4140
rect 354036 4088 354088 4140
rect 365260 4088 365312 4140
rect 217324 4020 217376 4072
rect 276020 4020 276072 4072
rect 346952 4020 347004 4072
rect 364616 4020 364668 4072
rect 214748 3952 214800 4004
rect 262956 3952 263008 4004
rect 342168 3952 342220 4004
rect 362500 3952 362552 4004
rect 503076 3952 503128 4004
rect 537208 3952 537260 4004
rect 216496 3884 216548 3936
rect 277124 3884 277176 3936
rect 343364 3884 343416 3936
rect 362960 3884 363012 3936
rect 496084 3884 496136 3936
rect 533712 3884 533764 3936
rect 211068 3816 211120 3868
rect 272432 3816 272484 3868
rect 339868 3816 339920 3868
rect 364432 3816 364484 3868
rect 516784 3816 516836 3868
rect 554964 3816 555016 3868
rect 219164 3748 219216 3800
rect 280712 3748 280764 3800
rect 336280 3748 336332 3800
rect 364524 3748 364576 3800
rect 476764 3748 476816 3800
rect 523040 3748 523092 3800
rect 538956 3748 539008 3800
rect 559748 3748 559800 3800
rect 35992 3680 36044 3732
rect 46204 3680 46256 3732
rect 219348 3680 219400 3732
rect 287796 3680 287848 3732
rect 332692 3680 332744 3732
rect 364340 3680 364392 3732
rect 431224 3680 431276 3732
rect 479340 3680 479392 3732
rect 508504 3680 508556 3732
rect 551468 3680 551520 3732
rect 12348 3544 12400 3596
rect 13084 3544 13136 3596
rect 20628 3544 20680 3596
rect 43444 3612 43496 3664
rect 46664 3612 46716 3664
rect 28908 3544 28960 3596
rect 32404 3544 32456 3596
rect 38384 3544 38436 3596
rect 39304 3544 39356 3596
rect 51356 3544 51408 3596
rect 53104 3544 53156 3596
rect 53748 3544 53800 3596
rect 54484 3544 54536 3596
rect 60832 3612 60884 3664
rect 79324 3612 79376 3664
rect 85672 3612 85724 3664
rect 106924 3612 106976 3664
rect 114008 3612 114060 3664
rect 182824 3612 182876 3664
rect 116584 3544 116636 3596
rect 118700 3544 118752 3596
rect 119896 3544 119948 3596
rect 121092 3544 121144 3596
rect 189724 3612 189776 3664
rect 216404 3612 216456 3664
rect 284300 3612 284352 3664
rect 325608 3612 325660 3664
rect 358360 3612 358412 3664
rect 457444 3612 457496 3664
rect 187332 3544 187384 3596
rect 188344 3544 188396 3596
rect 193220 3544 193272 3596
rect 194416 3544 194468 3596
rect 195612 3544 195664 3596
rect 196624 3544 196676 3596
rect 219348 3544 219400 3596
rect 288992 3544 289044 3596
rect 329196 3544 329248 3596
rect 355508 3544 355560 3596
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 5264 3476 5316 3528
rect 75184 3476 75236 3528
rect 77300 3476 77352 3528
rect 78220 3476 78272 3528
rect 93860 3476 93912 3528
rect 94780 3476 94832 3528
rect 102140 3476 102192 3528
rect 103336 3476 103388 3528
rect 106924 3476 106976 3528
rect 178684 3476 178736 3528
rect 190828 3476 190880 3528
rect 192484 3476 192536 3528
rect 217416 3476 217468 3528
rect 291384 3476 291436 3528
rect 324412 3476 324464 3528
rect 358084 3544 358136 3596
rect 377404 3544 377456 3596
rect 6460 3408 6512 3460
rect 8944 3408 8996 3460
rect 11152 3408 11204 3460
rect 30104 3408 30156 3460
rect 31024 3408 31076 3460
rect 33600 3408 33652 3460
rect 35256 3408 35308 3460
rect 43076 3408 43128 3460
rect 68284 3408 68336 3460
rect 69020 3408 69072 3460
rect 69940 3408 69992 3460
rect 99840 3408 99892 3460
rect 174544 3408 174596 3460
rect 182548 3408 182600 3460
rect 211804 3408 211856 3460
rect 213644 3408 213696 3460
rect 290188 3408 290240 3460
rect 322112 3408 322164 3460
rect 356704 3476 356756 3528
rect 374000 3476 374052 3528
rect 375288 3476 375340 3528
rect 411904 3544 411956 3596
rect 442264 3544 442316 3596
rect 398840 3476 398892 3528
rect 400128 3476 400180 3528
rect 407120 3476 407172 3528
rect 408408 3476 408460 3528
rect 415492 3476 415544 3528
rect 416688 3476 416740 3528
rect 423680 3476 423732 3528
rect 424968 3476 425020 3528
rect 432052 3476 432104 3528
rect 433248 3476 433300 3528
rect 440332 3476 440384 3528
rect 441528 3476 441580 3528
rect 448612 3476 448664 3528
rect 449808 3476 449860 3528
rect 456800 3544 456852 3596
rect 458088 3544 458140 3596
rect 467104 3612 467156 3664
rect 519544 3612 519596 3664
rect 534724 3612 534776 3664
rect 541992 3612 542044 3664
rect 552756 3612 552808 3664
rect 573916 3612 573968 3664
rect 515956 3544 516008 3596
rect 525064 3544 525116 3596
rect 531320 3544 531372 3596
rect 532148 3544 532200 3596
rect 538864 3544 538916 3596
rect 583392 3544 583444 3596
rect 505376 3476 505428 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 572720 3476 572772 3528
rect 356336 3408 356388 3460
rect 363052 3408 363104 3460
rect 382280 3408 382332 3460
rect 383568 3408 383620 3460
rect 390560 3408 390612 3460
rect 391848 3408 391900 3460
rect 34796 3340 34848 3392
rect 36544 3340 36596 3392
rect 56048 3340 56100 3392
rect 57244 3340 57296 3392
rect 59636 3340 59688 3392
rect 61384 3340 61436 3392
rect 212448 3340 212500 3392
rect 258264 3340 258316 3392
rect 355232 3340 355284 3392
rect 365904 3340 365956 3392
rect 387064 3340 387116 3392
rect 429660 3408 429712 3460
rect 432604 3408 432656 3460
rect 501788 3408 501840 3460
rect 520924 3408 520976 3460
rect 569132 3408 569184 3460
rect 473360 3340 473412 3392
rect 474188 3340 474240 3392
rect 481640 3340 481692 3392
rect 482468 3340 482520 3392
rect 498200 3340 498252 3392
rect 499028 3340 499080 3392
rect 547880 3340 547932 3392
rect 548708 3340 548760 3392
rect 556160 3340 556212 3392
rect 556988 3340 557040 3392
rect 35164 3272 35216 3324
rect 213828 3272 213880 3324
rect 245200 3272 245252 3324
rect 355508 3272 355560 3324
rect 361672 3272 361724 3324
rect 47860 3204 47912 3256
rect 48964 3204 49016 3256
rect 215208 3204 215260 3256
rect 244096 3204 244148 3256
rect 352840 3204 352892 3256
rect 357440 3204 357492 3256
rect 1676 3136 1728 3188
rect 4896 3136 4948 3188
rect 205088 3136 205140 3188
rect 206284 3136 206336 3188
rect 19432 2932 19484 2984
rect 25504 2932 25556 2984
rect 41880 2932 41932 2984
rect 43536 2932 43588 2984
rect 365720 1232 365772 1284
rect 367008 1232 367060 1284
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657014 2820 658135
rect 2780 657008 2832 657014
rect 2780 656950 2832 656956
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 2792 553722 2820 553823
rect 2780 553716 2832 553722
rect 2780 553658 2832 553664
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3436 449206 3464 671191
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3528 579834 3556 579935
rect 3516 579828 3568 579834
rect 3516 579770 3568 579776
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 449200 3476 449206
rect 3424 449142 3476 449148
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3528 447846 3556 514791
rect 3606 501800 3662 501809
rect 3606 501735 3662 501744
rect 3620 474026 3648 501735
rect 3608 474020 3660 474026
rect 3608 473962 3660 473968
rect 4816 450634 4844 683674
rect 4896 657008 4948 657014
rect 4896 656950 4948 656956
rect 4908 453422 4936 656950
rect 4988 632120 5040 632126
rect 4988 632062 5040 632068
rect 4896 453416 4948 453422
rect 4896 453358 4948 453364
rect 4804 450628 4856 450634
rect 4804 450570 4856 450576
rect 5000 450566 5028 632062
rect 5080 553716 5132 553722
rect 5080 553658 5132 553664
rect 5092 453354 5120 553658
rect 5080 453348 5132 453354
rect 5080 453290 5132 453296
rect 6932 451926 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 10324 605872 10376 605878
rect 10324 605814 10376 605820
rect 8944 579828 8996 579834
rect 8944 579770 8996 579776
rect 6920 451920 6972 451926
rect 6920 451862 6972 451868
rect 8956 450702 8984 579770
rect 10336 453490 10364 605814
rect 10416 527196 10468 527202
rect 10416 527138 10468 527144
rect 10324 453484 10376 453490
rect 10324 453426 10376 453432
rect 10428 451994 10456 527138
rect 10416 451988 10468 451994
rect 10416 451930 10468 451936
rect 8944 450696 8996 450702
rect 8944 450638 8996 450644
rect 4988 450560 5040 450566
rect 4988 450502 5040 450508
rect 23492 447914 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 32404 618316 32456 618322
rect 32404 618258 32456 618264
rect 32416 453558 32444 618258
rect 32404 453552 32456 453558
rect 32404 453494 32456 453500
rect 23480 447908 23532 447914
rect 23480 447850 23532 447856
rect 3516 447840 3568 447846
rect 3516 447782 3568 447788
rect 40052 446418 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 452062 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 84844 565888 84896 565894
rect 84844 565830 84896 565836
rect 84856 453762 84884 565830
rect 84844 453756 84896 453762
rect 84844 453698 84896 453704
rect 71780 452056 71832 452062
rect 71780 451998 71832 452004
rect 88352 448050 88380 702406
rect 105464 699718 105492 703520
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 106936 449274 106964 699654
rect 106924 449268 106976 449274
rect 106924 449210 106976 449216
rect 88340 448044 88392 448050
rect 88340 447986 88392 447992
rect 136652 446486 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 448186 153240 702406
rect 169772 449342 169800 702406
rect 169760 449336 169812 449342
rect 169760 449278 169812 449284
rect 153200 448180 153252 448186
rect 153200 448122 153252 448128
rect 201512 446554 201540 702986
rect 217968 565140 218020 565146
rect 217968 565082 218020 565088
rect 217874 516896 217930 516905
rect 217874 516831 217930 516840
rect 217782 515944 217838 515953
rect 217782 515879 217838 515888
rect 217690 513768 217746 513777
rect 217690 513703 217746 513712
rect 217598 489968 217654 489977
rect 217598 489903 217654 489912
rect 217322 488336 217378 488345
rect 217322 488271 217378 488280
rect 217336 475386 217364 488271
rect 217506 488064 217562 488073
rect 217506 487999 217562 488008
rect 217324 475380 217376 475386
rect 217324 475322 217376 475328
rect 217520 456074 217548 487999
rect 217612 456142 217640 489903
rect 217704 478174 217732 513703
rect 217692 478168 217744 478174
rect 217692 478110 217744 478116
rect 217796 468518 217824 515879
rect 217784 468512 217836 468518
rect 217784 468454 217836 468460
rect 217600 456136 217652 456142
rect 217600 456078 217652 456084
rect 217508 456068 217560 456074
rect 217508 456010 217560 456016
rect 217888 454714 217916 516831
rect 217876 454708 217928 454714
rect 217876 454650 217928 454656
rect 201500 446548 201552 446554
rect 201500 446490 201552 446496
rect 136640 446480 136692 446486
rect 136640 446422 136692 446428
rect 40040 446412 40092 446418
rect 40040 446354 40092 446360
rect 178776 445460 178828 445466
rect 178776 445402 178828 445408
rect 7564 445392 7616 445398
rect 7564 445334 7616 445340
rect 3424 443692 3476 443698
rect 3424 443634 3476 443640
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 2872 398812 2924 398818
rect 2872 398754 2924 398760
rect 2884 397497 2912 398754
rect 2870 397488 2926 397497
rect 2870 397423 2926 397432
rect 2872 372564 2924 372570
rect 2872 372506 2924 372512
rect 2884 371385 2912 372506
rect 2870 371376 2926 371385
rect 2870 371311 2926 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 267708 3384 267714
rect 3332 267650 3384 267656
rect 3344 267209 3372 267650
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 2780 264240 2832 264246
rect 2780 264182 2832 264188
rect 2792 16574 2820 264182
rect 2872 254244 2924 254250
rect 2872 254186 2924 254192
rect 2884 254153 2912 254186
rect 2870 254144 2926 254153
rect 2870 254079 2926 254088
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 84697 3464 443634
rect 4896 443012 4948 443018
rect 4896 442954 4948 442960
rect 3516 442536 3568 442542
rect 3516 442478 3568 442484
rect 3528 136785 3556 442478
rect 3792 442468 3844 442474
rect 3792 442410 3844 442416
rect 3608 442264 3660 442270
rect 3608 442206 3660 442212
rect 3620 188873 3648 442206
rect 3700 439544 3752 439550
rect 3700 439486 3752 439492
rect 3712 201929 3740 439486
rect 3804 241097 3832 442410
rect 3976 442400 4028 442406
rect 3976 442342 4028 442348
rect 3884 442332 3936 442338
rect 3884 442274 3936 442280
rect 3896 293185 3924 442274
rect 3988 345409 4016 442342
rect 3974 345400 4030 345409
rect 3974 345335 4030 345344
rect 3882 293176 3938 293185
rect 3882 293111 3938 293120
rect 4804 258732 4856 258738
rect 4804 258674 4856 258680
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3608 150408 3660 150414
rect 3608 150350 3660 150356
rect 3620 149841 3648 150350
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97640 3568 97646
rect 3514 97608 3516 97617
rect 3568 97608 3570 97617
rect 3514 97543 3570 97552
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 2792 16546 3648 16574
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1688 480 1716 3130
rect 2884 480 2912 4082
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 4816 3534 4844 258674
rect 4908 254250 4936 442954
rect 4896 254244 4948 254250
rect 4896 254186 4948 254192
rect 6920 246356 6972 246362
rect 6920 246298 6972 246304
rect 4896 244928 4948 244934
rect 4896 244870 4948 244876
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4908 3194 4936 244870
rect 6932 6914 6960 246298
rect 7576 97646 7604 445334
rect 174544 443420 174596 443426
rect 174544 443362 174596 443368
rect 84844 443352 84896 443358
rect 84844 443294 84896 443300
rect 32404 443148 32456 443154
rect 32404 443090 32456 443096
rect 8944 443080 8996 443086
rect 8944 443022 8996 443028
rect 8956 423638 8984 443022
rect 8944 423632 8996 423638
rect 8944 423574 8996 423580
rect 32416 372570 32444 443090
rect 32404 372564 32456 372570
rect 32404 372506 32456 372512
rect 84856 320142 84884 443294
rect 84844 320136 84896 320142
rect 84844 320078 84896 320084
rect 68284 308780 68336 308786
rect 68284 308722 68336 308728
rect 43444 308712 43496 308718
rect 43444 308654 43496 308660
rect 35164 308576 35216 308582
rect 35164 308518 35216 308524
rect 32404 308508 32456 308514
rect 32404 308450 32456 308456
rect 25504 308440 25556 308446
rect 25504 308382 25556 308388
rect 22100 271176 22152 271182
rect 22100 271118 22152 271124
rect 13820 269816 13872 269822
rect 13820 269758 13872 269764
rect 8300 267028 8352 267034
rect 8300 266970 8352 266976
rect 7656 244996 7708 245002
rect 7656 244938 7708 244944
rect 7564 97640 7616 97646
rect 7564 97582 7616 97588
rect 7668 16574 7696 244938
rect 8312 16574 8340 266970
rect 8944 256012 8996 256018
rect 8944 255954 8996 255960
rect 7668 16546 7788 16574
rect 8312 16546 8800 16574
rect 6932 6886 7696 6914
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5276 480 5304 3470
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 6886
rect 7760 4146 7788 16546
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8772 480 8800 16546
rect 8956 3466 8984 255954
rect 9680 253224 9732 253230
rect 9680 253166 9732 253172
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 253166
rect 12440 251864 12492 251870
rect 12440 251806 12492 251812
rect 12452 16574 12480 251806
rect 13084 246424 13136 246430
rect 13084 246366 13136 246372
rect 12452 16546 13032 16574
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 12360 480 12388 3538
rect 13004 3482 13032 16546
rect 13096 3602 13124 246366
rect 13832 16574 13860 269758
rect 17224 256080 17276 256086
rect 17224 256022 17276 256028
rect 16580 250504 16632 250510
rect 16580 250446 16632 250452
rect 16592 16574 16620 250446
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13004 3454 13584 3482
rect 13556 480 13584 3454
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 480 15976 4082
rect 17052 480 17080 16546
rect 17236 4146 17264 256022
rect 17960 253292 18012 253298
rect 17960 253234 18012 253240
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 253234
rect 20720 251932 20772 251938
rect 20720 251874 20772 251880
rect 20732 16574 20760 251874
rect 22112 16574 22140 271118
rect 24860 256148 24912 256154
rect 24860 256090 24912 256096
rect 24872 16574 24900 256090
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 24872 16546 25360 16574
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 480 19472 2926
rect 20640 480 20668 3538
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24228 480 24256 4082
rect 25332 480 25360 16546
rect 25516 2990 25544 308382
rect 31760 283620 31812 283626
rect 31760 283562 31812 283568
rect 26884 276684 26936 276690
rect 26884 276626 26936 276632
rect 26240 252000 26292 252006
rect 26240 251942 26292 251948
rect 25504 2984 25556 2990
rect 25504 2926 25556 2932
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 251942
rect 26896 4146 26924 276626
rect 30380 273964 30432 273970
rect 30380 273906 30432 273912
rect 27620 272536 27672 272542
rect 27620 272478 27672 272484
rect 27632 16574 27660 272478
rect 30392 16574 30420 273906
rect 31024 252068 31076 252074
rect 31024 252010 31076 252016
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 27724 480 27752 16546
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28920 480 28948 3538
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 30116 480 30144 3402
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31036 3466 31064 252010
rect 31772 16574 31800 283562
rect 31772 16546 31984 16574
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3602 32444 308450
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 480 33640 3402
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 34808 480 34836 3334
rect 35176 3330 35204 308518
rect 38660 287700 38712 287706
rect 38660 287642 38712 287648
rect 36544 280832 36596 280838
rect 36544 280774 36596 280780
rect 35900 260160 35952 260166
rect 35900 260102 35952 260108
rect 35256 258800 35308 258806
rect 35256 258742 35308 258748
rect 35268 3466 35296 258742
rect 35912 16574 35940 260102
rect 35912 16546 36492 16574
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 35256 3460 35308 3466
rect 35256 3402 35308 3408
rect 35164 3324 35216 3330
rect 35164 3266 35216 3272
rect 36004 480 36032 3674
rect 36464 490 36492 16546
rect 36556 3398 36584 280774
rect 38672 16574 38700 287642
rect 40040 262880 40092 262886
rect 40040 262822 40092 262828
rect 39304 254584 39356 254590
rect 39304 254526 39356 254532
rect 38672 16546 39160 16574
rect 38384 3596 38436 3602
rect 38384 3538 38436 3544
rect 36544 3392 36596 3398
rect 36544 3334 36596 3340
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36464 462 36860 490
rect 38396 480 38424 3538
rect 36832 354 36860 462
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3602 39344 254526
rect 40052 16574 40080 262822
rect 40052 16546 40264 16574
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 43456 3670 43484 308654
rect 46204 308644 46256 308650
rect 46204 308586 46256 308592
rect 43536 282192 43588 282198
rect 43536 282134 43588 282140
rect 43444 3664 43496 3670
rect 43444 3606 43496 3612
rect 43076 3460 43128 3466
rect 43076 3402 43128 3408
rect 41880 2984 41932 2990
rect 41880 2926 41932 2932
rect 41892 480 41920 2926
rect 43088 480 43116 3402
rect 43548 2990 43576 282134
rect 44180 265668 44232 265674
rect 44180 265610 44232 265616
rect 44192 6914 44220 265610
rect 44272 254652 44324 254658
rect 44272 254594 44324 254600
rect 44284 16574 44312 254594
rect 44284 16546 45048 16574
rect 44192 6886 44312 6914
rect 43536 2984 43588 2990
rect 43536 2926 43588 2932
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46216 3738 46244 308586
rect 67640 307080 67692 307086
rect 67640 307022 67692 307028
rect 63500 287768 63552 287774
rect 63500 287710 63552 287716
rect 54484 286340 54536 286346
rect 54484 286282 54536 286288
rect 49700 284980 49752 284986
rect 49700 284922 49752 284928
rect 48320 267096 48372 267102
rect 48320 267038 48372 267044
rect 48332 16574 48360 267038
rect 48964 246492 49016 246498
rect 48964 246434 49016 246440
rect 48332 16546 48544 16574
rect 46204 3732 46256 3738
rect 46204 3674 46256 3680
rect 46664 3664 46716 3670
rect 46664 3606 46716 3612
rect 46676 480 46704 3606
rect 47860 3256 47912 3262
rect 47860 3198 47912 3204
rect 47872 480 47900 3198
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 48976 3262 49004 246434
rect 49712 16574 49740 284922
rect 52460 268388 52512 268394
rect 52460 268330 52512 268336
rect 52472 16574 52500 268330
rect 53840 247716 53892 247722
rect 53840 247658 53892 247664
rect 53104 246560 53156 246566
rect 53104 246502 53156 246508
rect 49712 16546 50200 16574
rect 52472 16546 52592 16574
rect 48964 3256 49016 3262
rect 48964 3198 49016 3204
rect 50172 480 50200 16546
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 51368 480 51396 3538
rect 52564 480 52592 16546
rect 53116 3602 53144 246502
rect 53852 16574 53880 247658
rect 53852 16546 54432 16574
rect 53104 3596 53156 3602
rect 53104 3538 53156 3544
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 53760 480 53788 3538
rect 54404 3482 54432 16546
rect 54496 3602 54524 286282
rect 61384 276820 61436 276826
rect 61384 276762 61436 276768
rect 57244 275324 57296 275330
rect 57244 275266 57296 275272
rect 56600 254720 56652 254726
rect 56600 254662 56652 254668
rect 56612 16574 56640 254662
rect 56612 16546 56824 16574
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 54404 3454 54984 3482
rect 54956 480 54984 3454
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56060 480 56088 3334
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3398 57284 275266
rect 60740 258868 60792 258874
rect 60740 258810 60792 258816
rect 57980 249076 58032 249082
rect 57980 249018 58032 249024
rect 57992 16574 58020 249018
rect 60752 16574 60780 258810
rect 57992 16546 58480 16574
rect 60752 16546 61332 16574
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 58452 480 58480 16546
rect 60832 3664 60884 3670
rect 60832 3606 60884 3612
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 59648 480 59676 3334
rect 60844 480 60872 3606
rect 61304 490 61332 16546
rect 61396 3398 61424 276762
rect 62120 276752 62172 276758
rect 62120 276694 62172 276700
rect 62132 16574 62160 276694
rect 63512 16574 63540 287710
rect 66260 278044 66312 278050
rect 66260 277986 66312 277992
rect 64880 260228 64932 260234
rect 64880 260170 64932 260176
rect 64892 16574 64920 260170
rect 66272 16574 66300 277986
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61384 3392 61436 3398
rect 61384 3334 61436 3340
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61304 462 61700 490
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61672 354 61700 462
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 307022
rect 68296 3466 68324 308722
rect 75182 308408 75238 308417
rect 75182 308343 75238 308352
rect 74540 290488 74592 290494
rect 74540 290430 74592 290436
rect 70400 289128 70452 289134
rect 70400 289070 70452 289076
rect 69020 279472 69072 279478
rect 69020 279414 69072 279420
rect 69032 3466 69060 279414
rect 69112 258936 69164 258942
rect 69112 258878 69164 258884
rect 68284 3460 68336 3466
rect 68284 3402 68336 3408
rect 69020 3460 69072 3466
rect 69020 3402 69072 3408
rect 69124 480 69152 258878
rect 70412 16574 70440 289070
rect 73160 282260 73212 282266
rect 73160 282202 73212 282208
rect 71780 250572 71832 250578
rect 71780 250514 71832 250520
rect 71792 16574 71820 250514
rect 73172 16574 73200 282202
rect 74552 16574 74580 290430
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69940 3460 69992 3466
rect 69940 3402 69992 3408
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3402
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 75196 3534 75224 308343
rect 124220 294636 124272 294642
rect 124220 294578 124272 294584
rect 117320 293412 117372 293418
rect 117320 293354 117372 293360
rect 110420 293344 110472 293350
rect 110420 293286 110472 293292
rect 102140 293276 102192 293282
rect 102140 293218 102192 293224
rect 95240 291984 95292 291990
rect 95240 291926 95292 291932
rect 92480 291916 92532 291922
rect 92480 291858 92532 291864
rect 88340 291848 88392 291854
rect 88340 291790 88392 291796
rect 81440 290624 81492 290630
rect 81440 290566 81492 290572
rect 77300 290556 77352 290562
rect 77300 290498 77352 290504
rect 75920 250640 75972 250646
rect 75920 250582 75972 250588
rect 75184 3528 75236 3534
rect 75184 3470 75236 3476
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 250582
rect 77312 3534 77340 290498
rect 77392 283688 77444 283694
rect 77392 283630 77444 283636
rect 77300 3528 77352 3534
rect 77300 3470 77352 3476
rect 77404 480 77432 283630
rect 79324 254788 79376 254794
rect 79324 254730 79376 254736
rect 78680 250708 78732 250714
rect 78680 250650 78732 250656
rect 78692 16574 78720 250650
rect 78692 16546 79272 16574
rect 78220 3528 78272 3534
rect 78220 3470 78272 3476
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3470
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 79336 3670 79364 254730
rect 80060 253360 80112 253366
rect 80060 253302 80112 253308
rect 80072 16574 80100 253302
rect 81452 16574 81480 290566
rect 85580 264308 85632 264314
rect 85580 264250 85632 264256
rect 82820 261520 82872 261526
rect 82820 261462 82872 261468
rect 82832 16574 82860 261462
rect 84200 253428 84252 253434
rect 84200 253370 84252 253376
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 79324 3664 79376 3670
rect 79324 3606 79376 3612
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 253370
rect 85592 16574 85620 264250
rect 86960 253496 87012 253502
rect 86960 253438 87012 253444
rect 86972 16574 87000 253438
rect 88352 16574 88380 291790
rect 91100 285048 91152 285054
rect 91100 284990 91152 284996
rect 89720 269884 89772 269890
rect 89720 269826 89772 269832
rect 89732 16574 89760 269826
rect 91112 16574 91140 284990
rect 85592 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85672 3664 85724 3670
rect 85672 3606 85724 3612
rect 85684 480 85712 3606
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 291858
rect 93860 286408 93912 286414
rect 93860 286350 93912 286356
rect 93872 3534 93900 286350
rect 93952 271244 94004 271250
rect 93952 271186 94004 271192
rect 93860 3528 93912 3534
rect 93860 3470 93912 3476
rect 93964 480 93992 271186
rect 95252 16574 95280 291926
rect 98000 286476 98052 286482
rect 98000 286418 98052 286424
rect 96620 282328 96672 282334
rect 96620 282270 96672 282276
rect 96632 16574 96660 282270
rect 98012 16574 98040 286418
rect 100760 283756 100812 283762
rect 100760 283698 100812 283704
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 94780 3528 94832 3534
rect 94780 3470 94832 3476
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3470
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99840 3460 99892 3466
rect 99840 3402 99892 3408
rect 99852 480 99880 3402
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 283698
rect 102152 3534 102180 293218
rect 106924 290692 106976 290698
rect 106924 290634 106976 290640
rect 104900 287836 104952 287842
rect 104900 287778 104952 287784
rect 102232 286544 102284 286550
rect 102232 286486 102284 286492
rect 102140 3528 102192 3534
rect 102140 3470 102192 3476
rect 102244 480 102272 286486
rect 103520 283824 103572 283830
rect 103520 283766 103572 283772
rect 103532 16574 103560 283766
rect 104912 16574 104940 287778
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 106936 3670 106964 290634
rect 109040 287904 109092 287910
rect 109040 287846 109092 287852
rect 107660 283892 107712 283898
rect 107660 283834 107712 283840
rect 107672 16574 107700 283834
rect 107672 16546 108160 16574
rect 106924 3664 106976 3670
rect 106924 3606 106976 3612
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 106936 480 106964 3470
rect 108132 480 108160 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 287846
rect 110432 6914 110460 293286
rect 115940 289196 115992 289202
rect 115940 289138 115992 289144
rect 111800 287972 111852 287978
rect 111800 287914 111852 287920
rect 110512 285116 110564 285122
rect 110512 285058 110564 285064
rect 110524 16574 110552 285058
rect 111812 16574 111840 287914
rect 114560 285184 114612 285190
rect 114560 285126 114612 285132
rect 114572 16574 114600 285126
rect 115952 16574 115980 289138
rect 116584 254856 116636 254862
rect 116584 254798 116636 254804
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 3664 114060 3670
rect 114008 3606 114060 3612
rect 114020 480 114048 3606
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 116596 3602 116624 254798
rect 116584 3596 116636 3602
rect 116584 3538 116636 3544
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 293354
rect 122840 289332 122892 289338
rect 122840 289274 122892 289280
rect 118700 289264 118752 289270
rect 118700 289206 118752 289212
rect 118712 3602 118740 289206
rect 118792 285252 118844 285258
rect 118792 285194 118844 285200
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 118804 480 118832 285194
rect 121460 252136 121512 252142
rect 121460 252078 121512 252084
rect 121472 16574 121500 252078
rect 122852 16574 122880 289274
rect 124232 16574 124260 294578
rect 160100 282464 160152 282470
rect 160100 282406 160152 282412
rect 155960 282396 156012 282402
rect 155960 282338 156012 282344
rect 151820 280968 151872 280974
rect 151820 280910 151872 280916
rect 149060 280900 149112 280906
rect 149060 280842 149112 280848
rect 144920 279540 144972 279546
rect 144920 279482 144972 279488
rect 142160 278112 142212 278118
rect 142160 278054 142212 278060
rect 138020 274032 138072 274038
rect 138020 273974 138072 273980
rect 131120 272604 131172 272610
rect 131120 272546 131172 272552
rect 126980 265736 127032 265742
rect 126980 265678 127032 265684
rect 125600 260296 125652 260302
rect 125600 260238 125652 260244
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 121092 3596 121144 3602
rect 121092 3538 121144 3544
rect 119908 480 119936 3538
rect 121104 480 121132 3538
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 260238
rect 126992 480 127020 265678
rect 128360 261588 128412 261594
rect 128360 261530 128412 261536
rect 127072 247784 127124 247790
rect 127072 247726 127124 247732
rect 127084 16574 127112 247726
rect 128372 16574 128400 261530
rect 129740 245064 129792 245070
rect 129740 245006 129792 245012
rect 129752 16574 129780 245006
rect 131132 16574 131160 272546
rect 136640 269952 136692 269958
rect 136640 269894 136692 269900
rect 133880 268456 133932 268462
rect 133880 268398 133932 268404
rect 132500 262948 132552 262954
rect 132500 262890 132552 262896
rect 132512 16574 132540 262890
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 268398
rect 135260 249144 135312 249150
rect 135260 249086 135312 249092
rect 135272 480 135300 249086
rect 135352 245132 135404 245138
rect 135352 245074 135404 245080
rect 135364 16574 135392 245074
rect 136652 16574 136680 269894
rect 138032 16574 138060 273974
rect 140780 271312 140832 271318
rect 140780 271254 140832 271260
rect 139400 264376 139452 264382
rect 139400 264318 139452 264324
rect 139412 16574 139440 264318
rect 140792 16574 140820 271254
rect 135364 16546 136496 16574
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136468 480 136496 16546
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 278054
rect 143540 247852 143592 247858
rect 143540 247794 143592 247800
rect 143552 11762 143580 247794
rect 143632 245200 143684 245206
rect 143632 245142 143684 245148
rect 143540 11756 143592 11762
rect 143540 11698 143592 11704
rect 143644 6914 143672 245142
rect 144932 16574 144960 279482
rect 146300 265804 146352 265810
rect 146300 265746 146352 265752
rect 146312 16574 146340 265746
rect 147680 247920 147732 247926
rect 147680 247862 147732 247868
rect 147692 16574 147720 247862
rect 149072 16574 149100 280842
rect 150440 267164 150492 267170
rect 150440 267106 150492 267112
rect 150452 16574 150480 267106
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144736 11756 144788 11762
rect 144736 11698 144788 11704
rect 143552 6886 143672 6914
rect 143552 480 143580 6886
rect 144748 480 144776 11698
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 9674 151860 280910
rect 154580 272672 154632 272678
rect 154580 272614 154632 272620
rect 153200 267232 153252 267238
rect 153200 267174 153252 267180
rect 151912 247988 151964 247994
rect 151912 247930 151964 247936
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 247930
rect 153212 16574 153240 267174
rect 154592 16574 154620 272614
rect 155972 16574 156000 282338
rect 158720 274100 158772 274106
rect 158720 274042 158772 274048
rect 157340 268524 157392 268530
rect 157340 268466 157392 268472
rect 157352 16574 157380 268466
rect 158732 16574 158760 274042
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 480 160140 282406
rect 173900 276956 173952 276962
rect 173900 276898 173952 276904
rect 169760 276888 169812 276894
rect 169760 276830 169812 276836
rect 167000 275460 167052 275466
rect 167000 275402 167052 275408
rect 162860 275392 162912 275398
rect 162860 275334 162912 275340
rect 161480 268592 161532 268598
rect 161480 268534 161532 268540
rect 160192 261656 160244 261662
rect 160192 261598 160244 261604
rect 160204 16574 160232 261598
rect 161492 16574 161520 268534
rect 162872 16574 162900 275334
rect 165620 268660 165672 268666
rect 165620 268602 165672 268608
rect 164240 261724 164292 261730
rect 164240 261666 164292 261672
rect 164252 16574 164280 261666
rect 165632 16574 165660 268602
rect 167012 16574 167040 275402
rect 168380 270020 168432 270026
rect 168380 269962 168432 269968
rect 160204 16546 161336 16574
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161308 480 161336 16546
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 11762 168420 269962
rect 168472 261792 168524 261798
rect 168472 261734 168524 261740
rect 168380 11756 168432 11762
rect 168380 11698 168432 11704
rect 168484 6914 168512 261734
rect 169772 16574 169800 276830
rect 172520 270088 172572 270094
rect 172520 270030 172572 270036
rect 171140 263016 171192 263022
rect 171140 262958 171192 262964
rect 171152 16574 171180 262958
rect 172532 16574 172560 270030
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 169576 11756 169628 11762
rect 169576 11698 169628 11704
rect 168392 6886 168512 6914
rect 168392 480 168420 6886
rect 169588 480 169616 11698
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 276898
rect 174556 267714 174584 443362
rect 178684 308848 178736 308854
rect 178684 308790 178736 308796
rect 178040 307148 178092 307154
rect 178040 307090 178092 307096
rect 176660 278180 176712 278186
rect 176660 278122 176712 278128
rect 174544 267708 174596 267714
rect 174544 267650 174596 267656
rect 175280 263084 175332 263090
rect 175280 263026 175332 263032
rect 174544 250776 174596 250782
rect 174544 250718 174596 250724
rect 174556 3466 174584 250718
rect 175292 16574 175320 263026
rect 175292 16546 175504 16574
rect 174544 3460 174596 3466
rect 174544 3402 174596 3408
rect 175476 480 175504 16546
rect 176672 11762 176700 278122
rect 176752 270156 176804 270162
rect 176752 270098 176804 270104
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 176764 6914 176792 270098
rect 178052 16574 178080 307090
rect 178052 16546 178632 16574
rect 177856 11756 177908 11762
rect 177856 11698 177908 11704
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11698
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3534 178724 308790
rect 178788 150414 178816 445402
rect 217980 445058 218008 565082
rect 218072 465730 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 565146 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700330 267688 703520
rect 283852 700398 283880 703520
rect 300136 700466 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 331232 565146 331260 702986
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 357532 700528 357584 700534
rect 357532 700470 357584 700476
rect 357440 700392 357492 700398
rect 357440 700334 357492 700340
rect 234620 565140 234672 565146
rect 234620 565082 234672 565088
rect 331220 565140 331272 565146
rect 331220 565082 331272 565088
rect 219070 512816 219126 512825
rect 219070 512751 219126 512760
rect 219084 478242 219112 512751
rect 219346 511048 219402 511057
rect 219346 510983 219402 510992
rect 219254 509960 219310 509969
rect 219254 509895 219310 509904
rect 219162 508192 219218 508201
rect 219162 508127 219218 508136
rect 219072 478236 219124 478242
rect 219072 478178 219124 478184
rect 219176 474094 219204 508127
rect 219164 474088 219216 474094
rect 219164 474030 219216 474036
rect 218060 465724 218112 465730
rect 218060 465666 218112 465672
rect 219268 454850 219296 509895
rect 219256 454844 219308 454850
rect 219256 454786 219308 454792
rect 219360 454782 219388 510983
rect 248420 478236 248472 478242
rect 248420 478178 248472 478184
rect 247038 476640 247094 476649
rect 241612 476604 241664 476610
rect 247038 476575 247094 476584
rect 241612 476546 241664 476552
rect 236092 476468 236144 476474
rect 236092 476410 236144 476416
rect 238852 476468 238904 476474
rect 238852 476410 238904 476416
rect 234620 476332 234672 476338
rect 234620 476274 234672 476280
rect 231860 475380 231912 475386
rect 231860 475322 231912 475328
rect 231872 460934 231900 475322
rect 231872 460906 232544 460934
rect 219348 454776 219400 454782
rect 219348 454718 219400 454724
rect 217968 445052 218020 445058
rect 217968 444994 218020 445000
rect 232412 444848 232464 444854
rect 232412 444790 232464 444796
rect 231216 444780 231268 444786
rect 231216 444722 231268 444728
rect 209044 444576 209096 444582
rect 209044 444518 209096 444524
rect 189724 309052 189776 309058
rect 189724 308994 189776 309000
rect 182824 308984 182876 308990
rect 182824 308926 182876 308932
rect 180800 278248 180852 278254
rect 180800 278190 180852 278196
rect 179420 271380 179472 271386
rect 179420 271322 179472 271328
rect 178776 150408 178828 150414
rect 178776 150350 178828 150356
rect 179432 16574 179460 271322
rect 180812 16574 180840 278190
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 178684 3528 178736 3534
rect 178684 3470 178736 3476
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 182836 3670 182864 308926
rect 187700 279608 187752 279614
rect 187700 279550 187752 279556
rect 184940 278316 184992 278322
rect 184940 278258 184992 278264
rect 183560 271448 183612 271454
rect 183560 271390 183612 271396
rect 183572 16574 183600 271390
rect 183572 16546 183784 16574
rect 182824 3664 182876 3670
rect 182824 3606 182876 3612
rect 182548 3460 182600 3466
rect 182548 3402 182600 3408
rect 182560 480 182588 3402
rect 183756 480 183784 16546
rect 184952 480 184980 278258
rect 185032 263152 185084 263158
rect 185032 263094 185084 263100
rect 185044 16574 185072 263094
rect 187712 16574 187740 279550
rect 188344 271516 188396 271522
rect 188344 271458 188396 271464
rect 185044 16546 186176 16574
rect 187712 16546 188292 16574
rect 186148 480 186176 16546
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 187344 480 187372 3538
rect 188264 3482 188292 16546
rect 188356 3602 188384 271458
rect 189080 264444 189132 264450
rect 189080 264386 189132 264392
rect 189092 16574 189120 264386
rect 189092 16546 189304 16574
rect 188344 3596 188396 3602
rect 188344 3538 188396 3544
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189736 3670 189764 308994
rect 207020 307216 207072 307222
rect 207020 307158 207072 307164
rect 205640 281104 205692 281110
rect 205640 281046 205692 281052
rect 198740 281036 198792 281042
rect 198740 280978 198792 280984
rect 196624 279744 196676 279750
rect 196624 279686 196676 279692
rect 191840 279676 191892 279682
rect 191840 279618 191892 279624
rect 191852 16574 191880 279618
rect 193220 272808 193272 272814
rect 193220 272750 193272 272756
rect 192484 272740 192536 272746
rect 192484 272682 192536 272688
rect 191852 16546 192064 16574
rect 189724 3664 189776 3670
rect 189724 3606 189776 3612
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 190840 480 190868 3470
rect 192036 480 192064 16546
rect 192496 3534 192524 272682
rect 193232 3602 193260 272750
rect 195980 264580 196032 264586
rect 195980 264522 196032 264528
rect 193312 264512 193364 264518
rect 193312 264454 193364 264460
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 192484 3528 192536 3534
rect 193324 3482 193352 264454
rect 195992 16574 196020 264522
rect 195992 16546 196572 16574
rect 194416 3596 194468 3602
rect 194416 3538 194468 3544
rect 195612 3596 195664 3602
rect 195612 3538 195664 3544
rect 192484 3470 192536 3476
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3538
rect 195624 480 195652 3538
rect 196544 3482 196572 16546
rect 196636 3602 196664 279686
rect 197360 272876 197412 272882
rect 197360 272818 197412 272824
rect 197372 16574 197400 272818
rect 197372 16546 197952 16574
rect 196624 3596 196676 3602
rect 196624 3538 196676 3544
rect 196544 3454 196848 3482
rect 196820 480 196848 3454
rect 197924 480 197952 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 280978
rect 201500 274168 201552 274174
rect 201500 274110 201552 274116
rect 200120 265872 200172 265878
rect 200120 265814 200172 265820
rect 200132 16574 200160 265814
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 274110
rect 202880 265940 202932 265946
rect 202880 265882 202932 265888
rect 201592 249212 201644 249218
rect 201592 249154 201644 249160
rect 201604 16574 201632 249154
rect 202892 16574 202920 265882
rect 205652 16574 205680 281046
rect 206284 274236 206336 274242
rect 206284 274178 206336 274184
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205088 3188 205140 3194
rect 205088 3130 205140 3136
rect 205100 480 205128 3130
rect 206204 480 206232 16546
rect 206296 3194 206324 274178
rect 206284 3188 206336 3194
rect 206284 3130 206336 3136
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 307158
rect 209056 111790 209084 444518
rect 231124 443556 231176 443562
rect 231124 443498 231176 443504
rect 216128 309120 216180 309126
rect 216128 309062 216180 309068
rect 213552 308916 213604 308922
rect 213552 308858 213604 308864
rect 212448 305856 212500 305862
rect 212448 305798 212500 305804
rect 212356 305720 212408 305726
rect 212356 305662 212408 305668
rect 210882 303376 210938 303385
rect 210882 303311 210938 303320
rect 210792 300416 210844 300422
rect 210792 300358 210844 300364
rect 210700 300348 210752 300354
rect 210700 300290 210752 300296
rect 209688 300144 209740 300150
rect 209688 300086 209740 300092
rect 209700 152590 209728 300086
rect 209780 266008 209832 266014
rect 209780 265950 209832 265956
rect 209688 152584 209740 152590
rect 209688 152526 209740 152532
rect 209044 111784 209096 111790
rect 209044 111726 209096 111732
rect 209792 9674 209820 265950
rect 209872 249280 209924 249286
rect 209872 249222 209924 249228
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 249222
rect 210712 193186 210740 300290
rect 210700 193180 210752 193186
rect 210700 193122 210752 193128
rect 210804 189038 210832 300358
rect 210896 189718 210924 303311
rect 211894 303240 211950 303249
rect 211712 303204 211764 303210
rect 211894 303175 211950 303184
rect 211712 303146 211764 303152
rect 211068 300212 211120 300218
rect 211068 300154 211120 300160
rect 210974 300112 211030 300121
rect 210974 300047 211030 300056
rect 210884 189712 210936 189718
rect 210884 189654 210936 189660
rect 210792 189032 210844 189038
rect 210792 188974 210844 188980
rect 210988 155281 211016 300047
rect 210974 155272 211030 155281
rect 210974 155207 211030 155216
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 208582 3360 208638 3369
rect 208582 3295 208638 3304
rect 208596 480 208624 3295
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 211080 3874 211108 300154
rect 211160 246628 211212 246634
rect 211160 246570 211212 246576
rect 211172 16574 211200 246570
rect 211724 159594 211752 303146
rect 211804 260364 211856 260370
rect 211804 260306 211856 260312
rect 211712 159588 211764 159594
rect 211712 159530 211764 159536
rect 211172 16546 211752 16574
rect 211068 3868 211120 3874
rect 211068 3810 211120 3816
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 211816 3466 211844 260306
rect 211908 158506 211936 303175
rect 211988 303068 212040 303074
rect 211988 303010 212040 303016
rect 212000 158710 212028 303010
rect 212078 302968 212134 302977
rect 212078 302903 212134 302912
rect 211988 158704 212040 158710
rect 211988 158646 212040 158652
rect 211896 158500 211948 158506
rect 211896 158442 211948 158448
rect 212092 158370 212120 302903
rect 212262 302832 212318 302841
rect 212262 302767 212318 302776
rect 212172 300280 212224 300286
rect 212172 300222 212224 300228
rect 212080 158364 212132 158370
rect 212080 158306 212132 158312
rect 212184 155310 212212 300222
rect 212276 158234 212304 302767
rect 212264 158228 212316 158234
rect 212264 158170 212316 158176
rect 212368 155446 212396 305662
rect 212356 155440 212408 155446
rect 212356 155382 212408 155388
rect 212172 155304 212224 155310
rect 212172 155246 212224 155252
rect 211804 3460 211856 3466
rect 211804 3402 211856 3408
rect 212460 3398 212488 305798
rect 213184 303340 213236 303346
rect 213184 303282 213236 303288
rect 213092 302932 213144 302938
rect 213092 302874 213144 302880
rect 213000 245268 213052 245274
rect 213000 245210 213052 245216
rect 213012 168978 213040 245210
rect 213000 168972 213052 168978
rect 213000 168914 213052 168920
rect 213104 158778 213132 302874
rect 213196 159526 213224 303282
rect 213368 303272 213420 303278
rect 213368 303214 213420 303220
rect 213276 300824 213328 300830
rect 213276 300766 213328 300772
rect 213184 159520 213236 159526
rect 213184 159462 213236 159468
rect 213092 158772 213144 158778
rect 213092 158714 213144 158720
rect 213288 155553 213316 300766
rect 213380 155825 213408 303214
rect 213460 300620 213512 300626
rect 213460 300562 213512 300568
rect 213366 155816 213422 155825
rect 213366 155751 213422 155760
rect 213274 155544 213330 155553
rect 213274 155479 213330 155488
rect 213472 152522 213500 300562
rect 213564 159390 213592 308858
rect 214564 306196 214616 306202
rect 214564 306138 214616 306144
rect 213828 303612 213880 303618
rect 213828 303554 213880 303560
rect 213736 303408 213788 303414
rect 213736 303350 213788 303356
rect 213644 245336 213696 245342
rect 213644 245278 213696 245284
rect 213552 159384 213604 159390
rect 213552 159326 213604 159332
rect 213460 152516 213512 152522
rect 213460 152458 213512 152464
rect 213366 3496 213422 3505
rect 213656 3466 213684 245278
rect 213748 4146 213776 303350
rect 213736 4140 213788 4146
rect 213736 4082 213788 4088
rect 213366 3431 213422 3440
rect 213644 3460 213696 3466
rect 212448 3392 212500 3398
rect 212448 3334 212500 3340
rect 213380 480 213408 3431
rect 213644 3402 213696 3408
rect 213840 3330 213868 303554
rect 214472 303544 214524 303550
rect 214472 303486 214524 303492
rect 214380 300552 214432 300558
rect 214380 300494 214432 300500
rect 214392 195294 214420 300494
rect 214380 195288 214432 195294
rect 214380 195230 214432 195236
rect 214484 159662 214512 303486
rect 214472 159656 214524 159662
rect 214472 159598 214524 159604
rect 214472 158840 214524 158846
rect 214472 158782 214524 158788
rect 214484 155038 214512 158782
rect 214576 157962 214604 306138
rect 214840 306060 214892 306066
rect 214840 306002 214892 306008
rect 214656 303136 214708 303142
rect 214656 303078 214708 303084
rect 214668 158846 214696 303078
rect 214746 300248 214802 300257
rect 214746 300183 214802 300192
rect 214656 158840 214708 158846
rect 214656 158782 214708 158788
rect 214654 158672 214710 158681
rect 214654 158607 214710 158616
rect 214564 157956 214616 157962
rect 214564 157898 214616 157904
rect 214668 157894 214696 158607
rect 214656 157888 214708 157894
rect 214656 157830 214708 157836
rect 214472 155032 214524 155038
rect 214472 154974 214524 154980
rect 214760 4010 214788 300183
rect 214748 4004 214800 4010
rect 214748 3946 214800 3952
rect 214470 3496 214526 3505
rect 214470 3431 214526 3440
rect 213828 3324 213880 3330
rect 213828 3266 213880 3272
rect 214484 480 214512 3431
rect 214852 3233 214880 306002
rect 215208 305992 215260 305998
rect 215208 305934 215260 305940
rect 214932 305584 214984 305590
rect 214932 305526 214984 305532
rect 214944 4049 214972 305526
rect 215116 305516 215168 305522
rect 215116 305458 215168 305464
rect 215024 305448 215076 305454
rect 215024 305390 215076 305396
rect 214930 4040 214986 4049
rect 214930 3975 214986 3984
rect 215036 3913 215064 305390
rect 215022 3904 215078 3913
rect 215022 3839 215078 3848
rect 215128 3777 215156 305458
rect 215114 3768 215170 3777
rect 215114 3703 215170 3712
rect 215220 3262 215248 305934
rect 215944 305924 215996 305930
rect 215944 305866 215996 305872
rect 215852 302796 215904 302802
rect 215852 302738 215904 302744
rect 215760 300756 215812 300762
rect 215760 300698 215812 300704
rect 215772 195838 215800 300698
rect 215760 195832 215812 195838
rect 215760 195774 215812 195780
rect 215864 155514 215892 302738
rect 215956 158098 215984 305866
rect 216036 303476 216088 303482
rect 216036 303418 216088 303424
rect 215944 158092 215996 158098
rect 215944 158034 215996 158040
rect 216048 155689 216076 303418
rect 216140 158166 216168 309062
rect 216220 308372 216272 308378
rect 216220 308314 216272 308320
rect 216232 158302 216260 308314
rect 216312 308304 216364 308310
rect 216312 308246 216364 308252
rect 216324 158438 216352 308246
rect 219072 308168 219124 308174
rect 219072 308110 219124 308116
rect 218888 306264 218940 306270
rect 218888 306206 218940 306212
rect 216588 306128 216640 306134
rect 216588 306070 216640 306076
rect 216404 300688 216456 300694
rect 216404 300630 216456 300636
rect 216312 158432 216364 158438
rect 216312 158374 216364 158380
rect 216220 158296 216272 158302
rect 216220 158238 216272 158244
rect 216128 158160 216180 158166
rect 216128 158102 216180 158108
rect 216218 158128 216274 158137
rect 216218 158063 216274 158072
rect 216232 157418 216260 158063
rect 216220 157412 216272 157418
rect 216220 157354 216272 157360
rect 216034 155680 216090 155689
rect 216034 155615 216090 155624
rect 215852 155508 215904 155514
rect 215852 155450 215904 155456
rect 216416 3670 216444 300630
rect 216496 300076 216548 300082
rect 216496 300018 216548 300024
rect 216508 3942 216536 300018
rect 216496 3936 216548 3942
rect 216496 3878 216548 3884
rect 216404 3664 216456 3670
rect 216404 3606 216456 3612
rect 215666 3496 215722 3505
rect 215666 3431 215722 3440
rect 215208 3256 215260 3262
rect 214838 3224 214894 3233
rect 215208 3198 215260 3204
rect 214838 3159 214894 3168
rect 215680 480 215708 3431
rect 216600 3369 216628 306070
rect 217876 305788 217928 305794
rect 217876 305730 217928 305736
rect 217692 305652 217744 305658
rect 217692 305594 217744 305600
rect 217508 304292 217560 304298
rect 217508 304234 217560 304240
rect 217416 302660 217468 302666
rect 217416 302602 217468 302608
rect 217048 300484 217100 300490
rect 217048 300426 217100 300432
rect 217060 193769 217088 300426
rect 217232 259004 217284 259010
rect 217232 258946 217284 258952
rect 217140 243568 217192 243574
rect 217140 243510 217192 243516
rect 217046 193760 217102 193769
rect 217046 193695 217102 193704
rect 216680 193180 216732 193186
rect 216680 193122 216732 193128
rect 216692 192817 216720 193122
rect 216678 192808 216734 192817
rect 216678 192743 216734 192752
rect 216680 189032 216732 189038
rect 216680 188974 216732 188980
rect 216692 188193 216720 188974
rect 216678 188184 216734 188193
rect 216678 188119 216734 188128
rect 217152 155106 217180 243510
rect 217244 169969 217272 258946
rect 217428 195945 217456 302602
rect 217520 196897 217548 304234
rect 217600 296336 217652 296342
rect 217600 296278 217652 296284
rect 217506 196888 217562 196897
rect 217506 196823 217562 196832
rect 217414 195936 217470 195945
rect 217414 195871 217470 195880
rect 217508 195832 217560 195838
rect 217508 195774 217560 195780
rect 217324 195288 217376 195294
rect 217324 195230 217376 195236
rect 217230 169960 217286 169969
rect 217230 169895 217286 169904
rect 217140 155100 217192 155106
rect 217140 155042 217192 155048
rect 217336 4078 217364 195230
rect 217416 168972 217468 168978
rect 217416 168914 217468 168920
rect 217324 4072 217376 4078
rect 217324 4014 217376 4020
rect 216862 3632 216918 3641
rect 216862 3567 216918 3576
rect 216586 3360 216642 3369
rect 216586 3295 216642 3304
rect 216876 480 216904 3567
rect 217428 3534 217456 168914
rect 217520 155242 217548 195774
rect 217612 168065 217640 296278
rect 217704 168337 217732 305594
rect 217784 299940 217836 299946
rect 217784 299882 217836 299888
rect 217690 168328 217746 168337
rect 217690 168263 217746 168272
rect 217598 168056 217654 168065
rect 217598 167991 217654 168000
rect 217796 155417 217824 299882
rect 217888 159458 217916 305730
rect 217968 302864 218020 302870
rect 217968 302806 218020 302812
rect 217876 159452 217928 159458
rect 217876 159394 217928 159400
rect 217980 155961 218008 302806
rect 218794 300384 218850 300393
rect 218794 300319 218850 300328
rect 218704 296268 218756 296274
rect 218704 296210 218756 296216
rect 218428 281172 218480 281178
rect 218428 281114 218480 281120
rect 218440 243545 218468 281114
rect 218520 252204 218572 252210
rect 218520 252146 218572 252152
rect 218426 243536 218482 243545
rect 218426 243471 218482 243480
rect 218532 191049 218560 252146
rect 218612 243636 218664 243642
rect 218612 243578 218664 243584
rect 218518 191040 218574 191049
rect 218518 190975 218574 190984
rect 218060 189712 218112 189718
rect 218060 189654 218112 189660
rect 217966 155952 218022 155961
rect 217966 155887 218022 155896
rect 217782 155408 217838 155417
rect 217782 155343 217838 155352
rect 217508 155236 217560 155242
rect 217508 155178 217560 155184
rect 218072 16574 218100 189654
rect 218624 155174 218652 243578
rect 218716 189961 218744 296210
rect 218702 189952 218758 189961
rect 218702 189887 218758 189896
rect 218808 171134 218836 300319
rect 218716 171106 218836 171134
rect 218716 155378 218744 171106
rect 218796 166320 218848 166326
rect 218796 166262 218848 166268
rect 218808 155650 218836 166262
rect 218900 158030 218928 306206
rect 218980 302728 219032 302734
rect 218980 302670 219032 302676
rect 218992 166326 219020 302670
rect 218980 166320 219032 166326
rect 218980 166262 219032 166268
rect 218978 158672 219034 158681
rect 218978 158607 218980 158616
rect 219032 158607 219034 158616
rect 218980 158578 219032 158584
rect 219084 158574 219112 308110
rect 231136 306338 231164 443498
rect 231228 358766 231256 444722
rect 232228 444644 232280 444650
rect 232228 444586 232280 444592
rect 231308 443488 231360 443494
rect 231308 443430 231360 443436
rect 231320 398818 231348 443430
rect 232240 439550 232268 444586
rect 232424 442626 232452 444790
rect 232516 442762 232544 460906
rect 233240 456136 233292 456142
rect 233240 456078 233292 456084
rect 233148 448588 233200 448594
rect 233148 448530 233200 448536
rect 233160 446758 233188 448530
rect 233148 446752 233200 446758
rect 233148 446694 233200 446700
rect 233252 446690 233280 456078
rect 233332 456068 233384 456074
rect 233332 456010 233384 456016
rect 233240 446684 233292 446690
rect 233240 446626 233292 446632
rect 233344 442762 233372 456010
rect 234632 446690 234660 476274
rect 235906 476232 235962 476241
rect 235906 476167 235962 476176
rect 235920 476134 235948 476167
rect 234712 476128 234764 476134
rect 234712 476070 234764 476076
rect 235908 476128 235960 476134
rect 235908 476070 235960 476076
rect 233884 446684 233936 446690
rect 233884 446626 233936 446632
rect 234620 446684 234672 446690
rect 234620 446626 234672 446632
rect 233896 442762 233924 446626
rect 234724 442762 234752 476070
rect 236104 460934 236132 476410
rect 238760 476400 238812 476406
rect 237470 476368 237526 476377
rect 238760 476342 238812 476348
rect 237470 476303 237526 476312
rect 236104 460906 236224 460934
rect 235540 446684 235592 446690
rect 235540 446626 235592 446632
rect 235552 442762 235580 446626
rect 236196 442762 236224 460906
rect 237484 442762 237512 476303
rect 237562 476232 237618 476241
rect 237562 476167 237618 476176
rect 237576 460934 237604 476167
rect 237576 460906 237696 460934
rect 232516 442734 232806 442762
rect 233344 442734 233542 442762
rect 233896 442734 234278 442762
rect 234724 442734 235106 442762
rect 235552 442734 235842 442762
rect 236196 442734 236578 442762
rect 237406 442734 237512 442762
rect 237668 442762 237696 460906
rect 238772 446622 238800 476342
rect 238760 446616 238812 446622
rect 238760 446558 238812 446564
rect 238864 442762 238892 476410
rect 241520 476264 241572 476270
rect 240138 476232 240194 476241
rect 240138 476167 240194 476176
rect 241426 476232 241482 476241
rect 241520 476206 241572 476212
rect 241426 476167 241482 476176
rect 239404 446616 239456 446622
rect 239404 446558 239456 446564
rect 239416 442762 239444 446558
rect 240152 442762 240180 476167
rect 241440 476134 241468 476167
rect 241428 476128 241480 476134
rect 241428 476070 241480 476076
rect 240232 474088 240284 474094
rect 240232 474030 240284 474036
rect 240244 460934 240272 474030
rect 240244 460906 240824 460934
rect 240796 442762 240824 460906
rect 241532 442762 241560 476206
rect 241624 460934 241652 476546
rect 247052 476542 247080 476575
rect 247040 476536 247092 476542
rect 244278 476504 244334 476513
rect 247040 476478 247092 476484
rect 244278 476439 244280 476448
rect 244332 476439 244334 476448
rect 244280 476410 244332 476416
rect 245752 476400 245804 476406
rect 242898 476368 242954 476377
rect 242898 476303 242900 476312
rect 242952 476303 242954 476312
rect 244278 476368 244334 476377
rect 245752 476342 245804 476348
rect 244278 476303 244334 476312
rect 242900 476274 242952 476280
rect 244292 476270 244320 476303
rect 244280 476264 244332 476270
rect 242806 476232 242862 476241
rect 244280 476206 244332 476212
rect 245658 476232 245714 476241
rect 242806 476167 242808 476176
rect 242860 476167 242862 476176
rect 244924 476196 244976 476202
rect 242808 476138 242860 476144
rect 245658 476167 245714 476176
rect 244924 476138 244976 476144
rect 242900 476128 242952 476134
rect 242900 476070 242952 476076
rect 244372 476128 244424 476134
rect 244372 476070 244424 476076
rect 242912 460934 242940 476070
rect 244384 460934 244412 476070
rect 241624 460906 242296 460934
rect 242912 460906 243216 460934
rect 244384 460906 244688 460934
rect 242268 442762 242296 460906
rect 243188 442762 243216 460906
rect 244280 454844 244332 454850
rect 244280 454786 244332 454792
rect 237668 442734 238142 442762
rect 238864 442734 238970 442762
rect 239416 442734 239706 442762
rect 240152 442734 240442 442762
rect 240796 442734 241270 442762
rect 241532 442734 242006 442762
rect 242268 442734 242742 442762
rect 243188 442734 243570 442762
rect 244292 442748 244320 454786
rect 244660 442762 244688 460906
rect 244936 444990 244964 476138
rect 245672 476134 245700 476167
rect 245660 476128 245712 476134
rect 245660 476070 245712 476076
rect 244924 444984 244976 444990
rect 244924 444926 244976 444932
rect 245764 442762 245792 476342
rect 247222 476232 247278 476241
rect 247222 476167 247278 476176
rect 247236 460934 247264 476167
rect 247236 460906 247816 460934
rect 247132 454776 247184 454782
rect 247132 454718 247184 454724
rect 246580 444984 246632 444990
rect 246580 444926 246632 444932
rect 244660 442734 245134 442762
rect 245764 442734 245870 442762
rect 246592 442748 246620 444926
rect 247040 444712 247092 444718
rect 247040 444654 247092 444660
rect 247052 443698 247080 444654
rect 247040 443692 247092 443698
rect 247040 443634 247092 443640
rect 247144 442762 247172 454718
rect 247788 442762 247816 460906
rect 248432 446758 248460 478178
rect 251180 478168 251232 478174
rect 251180 478110 251232 478116
rect 311900 478168 311952 478174
rect 311900 478110 311952 478116
rect 249798 476640 249854 476649
rect 249798 476575 249854 476584
rect 249812 476542 249840 476575
rect 249800 476536 249852 476542
rect 249800 476478 249852 476484
rect 248512 476332 248564 476338
rect 248512 476274 248564 476280
rect 248420 446752 248472 446758
rect 248420 446694 248472 446700
rect 248524 442762 248552 476274
rect 249798 476232 249854 476241
rect 249798 476167 249854 476176
rect 251086 476232 251142 476241
rect 251086 476167 251088 476176
rect 249812 460934 249840 476167
rect 251140 476167 251142 476176
rect 251088 476138 251140 476144
rect 249812 460906 250024 460934
rect 249340 446752 249392 446758
rect 249340 446694 249392 446700
rect 249352 442762 249380 446694
rect 249996 442762 250024 460906
rect 251192 446758 251220 478110
rect 277766 477048 277822 477057
rect 277766 476983 277822 476992
rect 304998 477048 305054 477057
rect 304998 476983 305054 476992
rect 307758 477048 307814 477057
rect 307758 476983 307814 476992
rect 253846 476912 253902 476921
rect 253846 476847 253902 476856
rect 256606 476912 256662 476921
rect 256606 476847 256662 476856
rect 270498 476912 270554 476921
rect 270498 476847 270554 476856
rect 252558 476640 252614 476649
rect 252558 476575 252560 476584
rect 252612 476575 252614 476584
rect 252652 476604 252704 476610
rect 252560 476546 252612 476552
rect 252652 476546 252704 476552
rect 252374 476368 252430 476377
rect 252664 476320 252692 476546
rect 253860 476474 253888 476847
rect 255410 476776 255466 476785
rect 255410 476711 255466 476720
rect 255320 476536 255372 476542
rect 255320 476478 255372 476484
rect 253848 476468 253900 476474
rect 253848 476410 253900 476416
rect 252374 476303 252430 476312
rect 251272 476264 251324 476270
rect 251272 476206 251324 476212
rect 251180 446752 251232 446758
rect 251180 446694 251232 446700
rect 247144 442734 247434 442762
rect 247788 442734 248170 442762
rect 248524 442734 248906 442762
rect 249352 442734 249734 442762
rect 249996 442734 250470 442762
rect 251284 442748 251312 476206
rect 252388 476134 252416 476303
rect 252572 476292 252692 476320
rect 252466 476232 252522 476241
rect 252466 476167 252522 476176
rect 252376 476128 252428 476134
rect 252376 476070 252428 476076
rect 251732 446752 251784 446758
rect 251732 446694 251784 446700
rect 251744 442762 251772 446694
rect 252480 445262 252508 476167
rect 252572 446758 252600 476292
rect 252652 476196 252704 476202
rect 252652 476138 252704 476144
rect 252560 446752 252612 446758
rect 252560 446694 252612 446700
rect 252468 445256 252520 445262
rect 252468 445198 252520 445204
rect 252664 442762 252692 476138
rect 253940 476128 253992 476134
rect 253940 476070 253992 476076
rect 253952 446758 253980 476070
rect 254032 468512 254084 468518
rect 254032 468454 254084 468460
rect 253204 446752 253256 446758
rect 253204 446694 253256 446700
rect 253940 446752 253992 446758
rect 253940 446694 253992 446700
rect 253216 442762 253244 446694
rect 254044 442762 254072 468454
rect 254676 446752 254728 446758
rect 254676 446694 254728 446700
rect 254688 442762 254716 446694
rect 255332 443204 255360 476478
rect 255424 476406 255452 476711
rect 256620 476678 256648 476847
rect 258356 476740 258408 476746
rect 258356 476682 258408 476688
rect 256608 476672 256660 476678
rect 256608 476614 256660 476620
rect 258080 476468 258132 476474
rect 258080 476410 258132 476416
rect 255412 476400 255464 476406
rect 255412 476342 255464 476348
rect 257986 476368 258042 476377
rect 257986 476303 258042 476312
rect 255962 476232 256018 476241
rect 255962 476167 256018 476176
rect 255872 454708 255924 454714
rect 255872 454650 255924 454656
rect 255884 443204 255912 454650
rect 255976 445738 256004 476167
rect 255964 445732 256016 445738
rect 255964 445674 256016 445680
rect 257436 445256 257488 445262
rect 257436 445198 257488 445204
rect 255332 443176 255544 443204
rect 255884 443176 256280 443204
rect 255516 442762 255544 443176
rect 256252 442762 256280 443176
rect 251744 442734 252034 442762
rect 252664 442734 252770 442762
rect 253216 442734 253598 442762
rect 254044 442734 254334 442762
rect 254688 442734 255070 442762
rect 255516 442734 255898 442762
rect 256252 442734 256634 442762
rect 257448 442748 257476 445198
rect 258000 445126 258028 476303
rect 258092 446758 258120 476410
rect 258262 476368 258318 476377
rect 258262 476303 258264 476312
rect 258316 476303 258318 476312
rect 258264 476274 258316 476280
rect 258170 476232 258226 476241
rect 258170 476167 258172 476176
rect 258224 476167 258226 476176
rect 258172 476138 258224 476144
rect 258368 470594 258396 476682
rect 260104 476672 260156 476678
rect 260104 476614 260156 476620
rect 263598 476640 263654 476649
rect 259552 476468 259604 476474
rect 259552 476410 259604 476416
rect 258184 470566 258396 470594
rect 258080 446752 258132 446758
rect 258080 446694 258132 446700
rect 257988 445120 258040 445126
rect 257988 445062 258040 445068
rect 258184 442748 258212 470566
rect 258540 446752 258592 446758
rect 258540 446694 258592 446700
rect 258552 442762 258580 446694
rect 259564 442762 259592 476410
rect 260116 445738 260144 476614
rect 263598 476575 263600 476584
rect 263652 476575 263654 476584
rect 264978 476640 265034 476649
rect 264978 476575 265034 476584
rect 263600 476546 263652 476552
rect 264992 476542 265020 476575
rect 264980 476536 265032 476542
rect 260746 476504 260802 476513
rect 264980 476478 265032 476484
rect 267830 476504 267886 476513
rect 260746 476439 260802 476448
rect 267830 476439 267832 476448
rect 260760 476338 260788 476439
rect 267884 476439 267886 476448
rect 267832 476410 267884 476416
rect 270512 476406 270540 476847
rect 273166 476640 273222 476649
rect 273166 476575 273222 476584
rect 260932 476400 260984 476406
rect 260838 476368 260894 476377
rect 260748 476332 260800 476338
rect 270500 476400 270552 476406
rect 260932 476342 260984 476348
rect 267646 476368 267702 476377
rect 260838 476303 260894 476312
rect 260748 476274 260800 476280
rect 260852 476270 260880 476303
rect 260840 476264 260892 476270
rect 260746 476232 260802 476241
rect 260840 476206 260892 476212
rect 260746 476167 260802 476176
rect 260760 476134 260788 476167
rect 260748 476128 260800 476134
rect 260748 476070 260800 476076
rect 260104 445732 260156 445738
rect 260104 445674 260156 445680
rect 260472 445664 260524 445670
rect 260472 445606 260524 445612
rect 258552 442734 258934 442762
rect 259564 442734 259762 442762
rect 260484 442748 260512 445606
rect 260944 442762 260972 476342
rect 265624 476332 265676 476338
rect 270500 476342 270552 476348
rect 267646 476303 267702 476312
rect 265624 476274 265676 476280
rect 263692 476264 263744 476270
rect 262126 476232 262182 476241
rect 261484 476196 261536 476202
rect 263506 476232 263562 476241
rect 262126 476167 262182 476176
rect 262220 476196 262272 476202
rect 261484 476138 261536 476144
rect 261496 445330 261524 476138
rect 262140 467838 262168 476167
rect 263692 476206 263744 476212
rect 264886 476232 264942 476241
rect 263506 476167 263562 476176
rect 262220 476138 262272 476144
rect 262128 467832 262180 467838
rect 262128 467774 262180 467780
rect 262232 460934 262260 476138
rect 262864 476128 262916 476134
rect 262864 476070 262916 476076
rect 262232 460906 262352 460934
rect 262036 445732 262088 445738
rect 262036 445674 262088 445680
rect 261484 445324 261536 445330
rect 261484 445266 261536 445272
rect 260944 442734 261326 442762
rect 262048 442748 262076 445674
rect 262324 442762 262352 460906
rect 262876 445738 262904 476070
rect 263520 467226 263548 476167
rect 263508 467220 263560 467226
rect 263508 467162 263560 467168
rect 263704 460934 263732 476206
rect 264886 476167 264942 476176
rect 265164 476196 265216 476202
rect 264900 467294 264928 476167
rect 265164 476138 265216 476144
rect 264888 467288 264940 467294
rect 264888 467230 264940 467236
rect 265176 460934 265204 476138
rect 263704 460906 264008 460934
rect 265176 460906 265480 460934
rect 262864 445732 262916 445738
rect 262864 445674 262916 445680
rect 263600 445120 263652 445126
rect 263600 445062 263652 445068
rect 262324 442734 262798 442762
rect 263612 442748 263640 445062
rect 263980 442762 264008 460906
rect 265072 445324 265124 445330
rect 265072 445266 265124 445272
rect 263980 442734 264362 442762
rect 265084 442748 265112 445266
rect 265452 442762 265480 460906
rect 265636 445670 265664 476274
rect 266266 476232 266322 476241
rect 266266 476167 266322 476176
rect 267554 476232 267610 476241
rect 267554 476167 267610 476176
rect 266280 468586 266308 476167
rect 266268 468580 266320 468586
rect 266268 468522 266320 468528
rect 267568 468518 267596 476167
rect 267660 468654 267688 476303
rect 269026 476232 269082 476241
rect 269026 476167 269082 476176
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 271786 476232 271842 476241
rect 271786 476167 271842 476176
rect 267648 468648 267700 468654
rect 267648 468590 267700 468596
rect 267556 468512 267608 468518
rect 267556 468454 267608 468460
rect 269040 467158 269068 476167
rect 270420 469946 270448 476167
rect 270408 469940 270460 469946
rect 270408 469882 270460 469888
rect 269120 467832 269172 467838
rect 269120 467774 269172 467780
rect 269028 467152 269080 467158
rect 269028 467094 269080 467100
rect 269132 460934 269160 467774
rect 271800 467226 271828 476167
rect 273180 475386 273208 476575
rect 273258 476504 273314 476513
rect 273258 476439 273314 476448
rect 273272 476338 273300 476439
rect 274546 476368 274602 476377
rect 273260 476332 273312 476338
rect 274546 476303 274602 476312
rect 276018 476368 276074 476377
rect 276018 476303 276074 476312
rect 273260 476274 273312 476280
rect 274454 476232 274510 476241
rect 274454 476167 274510 476176
rect 273168 475380 273220 475386
rect 273168 475322 273220 475328
rect 273260 471300 273312 471306
rect 273260 471242 273312 471248
rect 271880 469872 271932 469878
rect 271880 469814 271932 469820
rect 270684 467220 270736 467226
rect 270684 467162 270736 467168
rect 271788 467220 271840 467226
rect 271788 467162 271840 467168
rect 270696 460934 270724 467162
rect 269132 460906 269344 460934
rect 270696 460906 270816 460934
rect 267096 454776 267148 454782
rect 267096 454718 267148 454724
rect 266636 445732 266688 445738
rect 266636 445674 266688 445680
rect 265624 445664 265676 445670
rect 265624 445606 265676 445612
rect 265452 442734 265926 442762
rect 266648 442748 266676 445674
rect 267108 442762 267136 454718
rect 268568 454708 268620 454714
rect 268568 454650 268620 454656
rect 268200 445732 268252 445738
rect 268200 445674 268252 445680
rect 267108 442734 267490 442762
rect 268212 442748 268240 445674
rect 268580 442762 268608 454650
rect 269316 442762 269344 460906
rect 270592 454844 270644 454850
rect 270592 454786 270644 454792
rect 270604 442762 270632 454786
rect 268580 442734 268962 442762
rect 269316 442734 269790 442762
rect 270526 442734 270632 442762
rect 270788 442762 270816 460906
rect 271892 442762 271920 469814
rect 271972 467288 272024 467294
rect 271972 467230 272024 467236
rect 271984 460934 272012 467230
rect 271984 460906 272472 460934
rect 272444 442762 272472 460906
rect 273272 442762 273300 471242
rect 274468 468586 274496 476167
rect 273352 468580 273404 468586
rect 273352 468522 273404 468528
rect 274456 468580 274508 468586
rect 274456 468522 274508 468528
rect 273364 460934 273392 468522
rect 274560 467294 274588 476303
rect 275926 476232 275982 476241
rect 275926 476167 275982 476176
rect 275940 468654 275968 476167
rect 276032 476134 276060 476303
rect 277780 476270 277808 476983
rect 302238 476776 302294 476785
rect 278780 476740 278832 476746
rect 302238 476711 302240 476720
rect 278780 476682 278832 476688
rect 302292 476711 302294 476720
rect 302240 476682 302292 476688
rect 277768 476264 277820 476270
rect 277306 476232 277362 476241
rect 277768 476206 277820 476212
rect 278686 476232 278742 476241
rect 277306 476167 277362 476176
rect 278686 476167 278742 476176
rect 276020 476128 276072 476134
rect 276020 476070 276072 476076
rect 277320 470014 277348 476167
rect 277308 470008 277360 470014
rect 277308 469950 277360 469956
rect 274640 468648 274692 468654
rect 274640 468590 274692 468596
rect 275928 468648 275980 468654
rect 275928 468590 275980 468596
rect 274548 467288 274600 467294
rect 274548 467230 274600 467236
rect 273364 460906 273944 460934
rect 273916 442762 273944 460906
rect 274652 446758 274680 468590
rect 278700 468518 278728 476167
rect 277400 468512 277452 468518
rect 277400 468454 277452 468460
rect 278688 468512 278740 468518
rect 278688 468454 278740 468460
rect 274732 456204 274784 456210
rect 274732 456146 274784 456152
rect 274640 446752 274692 446758
rect 274640 446694 274692 446700
rect 274744 442762 274772 456146
rect 276296 456136 276348 456142
rect 276296 456078 276348 456084
rect 275652 446752 275704 446758
rect 275652 446694 275704 446700
rect 275664 442762 275692 446694
rect 276308 442762 276336 456078
rect 270788 442734 271262 442762
rect 271892 442734 272090 442762
rect 272444 442734 272826 442762
rect 273272 442734 273654 442762
rect 273916 442734 274390 442762
rect 274744 442734 275126 442762
rect 275664 442734 275954 442762
rect 276308 442734 276690 442762
rect 277412 442748 277440 468454
rect 277768 456068 277820 456074
rect 277768 456010 277820 456016
rect 277780 442762 277808 456010
rect 278792 446758 278820 476682
rect 305012 476678 305040 476983
rect 280344 476672 280396 476678
rect 280344 476614 280396 476620
rect 305000 476672 305052 476678
rect 305000 476614 305052 476620
rect 280158 476368 280214 476377
rect 280158 476303 280214 476312
rect 280066 476232 280122 476241
rect 280172 476202 280200 476303
rect 280066 476167 280122 476176
rect 280160 476196 280212 476202
rect 280080 467158 280108 476167
rect 280160 476138 280212 476144
rect 280252 469940 280304 469946
rect 280252 469882 280304 469888
rect 278872 467152 278924 467158
rect 278872 467094 278924 467100
rect 280068 467152 280120 467158
rect 280068 467094 280120 467100
rect 278780 446752 278832 446758
rect 278780 446694 278832 446700
rect 278884 442762 278912 467094
rect 279516 446752 279568 446758
rect 279516 446694 279568 446700
rect 279528 442762 279556 446694
rect 280264 442762 280292 469882
rect 280356 460934 280384 476614
rect 284300 476604 284352 476610
rect 284300 476546 284352 476552
rect 281540 476536 281592 476542
rect 281540 476478 281592 476484
rect 280356 460906 280936 460934
rect 280908 442762 280936 460906
rect 281552 446758 281580 476478
rect 283010 476232 283066 476241
rect 283010 476167 283066 476176
rect 282920 475380 282972 475386
rect 282920 475322 282972 475328
rect 281632 467220 281684 467226
rect 281632 467162 281684 467168
rect 281540 446752 281592 446758
rect 281540 446694 281592 446700
rect 281644 442762 281672 467162
rect 282932 451274 282960 475322
rect 283024 454782 283052 476167
rect 283012 454776 283064 454782
rect 283012 454718 283064 454724
rect 282932 451246 283144 451274
rect 282460 446752 282512 446758
rect 282460 446694 282512 446700
rect 282472 442762 282500 446694
rect 283116 442762 283144 451246
rect 284312 442762 284340 476546
rect 307772 476542 307800 476983
rect 310518 476912 310574 476921
rect 310518 476847 310574 476856
rect 310532 476610 310560 476847
rect 310520 476604 310572 476610
rect 310520 476546 310572 476552
rect 307760 476536 307812 476542
rect 307760 476478 307812 476484
rect 285680 476468 285732 476474
rect 285680 476410 285732 476416
rect 284484 467288 284536 467294
rect 284484 467230 284536 467236
rect 284496 460934 284524 467230
rect 284496 460906 284800 460934
rect 284772 442762 284800 460906
rect 285692 442762 285720 476410
rect 287060 476400 287112 476406
rect 287060 476342 287112 476348
rect 285862 476232 285918 476241
rect 285862 476167 285918 476176
rect 285772 468580 285824 468586
rect 285772 468522 285824 468528
rect 285784 451274 285812 468522
rect 285876 454714 285904 476167
rect 285864 454708 285916 454714
rect 285864 454650 285916 454656
rect 285784 451246 286272 451274
rect 286244 442762 286272 451246
rect 287072 442762 287100 476342
rect 288440 476332 288492 476338
rect 288440 476274 288492 476280
rect 287242 476232 287298 476241
rect 287242 476167 287298 476176
rect 287152 468648 287204 468654
rect 287152 468590 287204 468596
rect 287164 451274 287192 468590
rect 287256 454850 287284 476167
rect 288452 460934 288480 476274
rect 289912 476264 289964 476270
rect 289818 476232 289874 476241
rect 289912 476206 289964 476212
rect 292670 476232 292726 476241
rect 289818 476167 289874 476176
rect 289832 469878 289860 476167
rect 289820 469872 289872 469878
rect 289820 469814 289872 469820
rect 288452 460906 288664 460934
rect 287244 454844 287296 454850
rect 287244 454786 287296 454792
rect 287164 451246 287928 451274
rect 287900 442762 287928 451246
rect 288636 442762 288664 460906
rect 289924 446758 289952 476206
rect 291200 476196 291252 476202
rect 292670 476167 292726 476176
rect 295338 476232 295394 476241
rect 295338 476167 295394 476176
rect 298098 476232 298154 476241
rect 298098 476167 298154 476176
rect 300858 476232 300914 476241
rect 300858 476167 300914 476176
rect 291200 476138 291252 476144
rect 290004 470008 290056 470014
rect 290004 469950 290056 469956
rect 289912 446752 289964 446758
rect 289912 446694 289964 446700
rect 290016 442762 290044 469950
rect 291212 446758 291240 476138
rect 292580 476128 292632 476134
rect 292580 476070 292632 476076
rect 291292 468512 291344 468518
rect 291292 468454 291344 468460
rect 290188 446752 290240 446758
rect 290188 446694 290240 446700
rect 291200 446752 291252 446758
rect 291200 446694 291252 446700
rect 277780 442734 278254 442762
rect 278884 442734 278990 442762
rect 279528 442734 279818 442762
rect 280264 442734 280554 442762
rect 280908 442734 281290 442762
rect 281644 442734 282118 442762
rect 282472 442734 282854 442762
rect 283116 442734 283590 442762
rect 284312 442734 284418 442762
rect 284772 442734 285154 442762
rect 285692 442734 285982 442762
rect 286244 442734 286718 442762
rect 287072 442734 287454 442762
rect 287900 442734 288282 442762
rect 288636 442734 289018 442762
rect 289846 442734 290044 442762
rect 290200 442762 290228 446694
rect 290200 442734 290582 442762
rect 291304 442748 291332 468454
rect 292592 446758 292620 476070
rect 292684 471306 292712 476167
rect 292672 471300 292724 471306
rect 292672 471242 292724 471248
rect 292672 467152 292724 467158
rect 292672 467094 292724 467100
rect 291844 446752 291896 446758
rect 291844 446694 291896 446700
rect 292580 446752 292632 446758
rect 292580 446694 292632 446700
rect 291856 442762 291884 446694
rect 292684 442762 292712 467094
rect 295352 456210 295380 476167
rect 295340 456204 295392 456210
rect 295340 456146 295392 456152
rect 298112 456142 298140 476167
rect 298100 456136 298152 456142
rect 298100 456078 298152 456084
rect 300872 456074 300900 476167
rect 300860 456068 300912 456074
rect 300860 456010 300912 456016
rect 302424 454844 302476 454850
rect 302424 454786 302476 454792
rect 300216 454776 300268 454782
rect 300216 454718 300268 454724
rect 298100 454708 298152 454714
rect 298100 454650 298152 454656
rect 296720 449404 296772 449410
rect 296720 449346 296772 449352
rect 293316 446752 293368 446758
rect 293316 446694 293368 446700
rect 293328 442762 293356 446694
rect 295982 444816 296038 444825
rect 295982 444751 296038 444760
rect 294418 444680 294474 444689
rect 294418 444615 294474 444624
rect 291856 442734 292146 442762
rect 292684 442734 292882 442762
rect 293328 442734 293618 442762
rect 294432 442748 294460 444615
rect 295154 444544 295210 444553
rect 295154 444479 295210 444488
rect 295168 442748 295196 444479
rect 295996 442748 296024 444751
rect 296732 442748 296760 449346
rect 297456 443216 297508 443222
rect 297456 443158 297508 443164
rect 297468 442748 297496 443158
rect 298112 442762 298140 454650
rect 299020 449472 299072 449478
rect 299020 449414 299072 449420
rect 298112 442734 298310 442762
rect 299032 442748 299060 449414
rect 299754 443320 299810 443329
rect 299754 443255 299810 443264
rect 299768 442748 299796 443255
rect 300228 442762 300256 454718
rect 301320 450832 301372 450838
rect 301320 450774 301372 450780
rect 300228 442734 300610 442762
rect 301332 442748 301360 450774
rect 302148 443284 302200 443290
rect 302148 443226 302200 443232
rect 302160 442748 302188 443226
rect 302436 442762 302464 454786
rect 307944 452192 307996 452198
rect 307944 452134 307996 452140
rect 303620 450900 303672 450906
rect 303620 450842 303672 450848
rect 302436 442734 302910 442762
rect 303632 442748 303660 450842
rect 305920 450764 305972 450770
rect 305920 450706 305972 450712
rect 305184 447976 305236 447982
rect 305184 447918 305236 447924
rect 304172 444916 304224 444922
rect 304172 444858 304224 444864
rect 232332 442598 232452 442626
rect 232228 439544 232280 439550
rect 232228 439486 232280 439492
rect 232332 412634 232360 442598
rect 304184 442542 304212 444858
rect 305196 442748 305224 447918
rect 305932 442748 305960 450706
rect 307484 448112 307536 448118
rect 307484 448054 307536 448060
rect 307496 442748 307524 448054
rect 307956 442762 307984 452134
rect 310520 452124 310572 452130
rect 310520 452066 310572 452072
rect 309784 448248 309836 448254
rect 309784 448190 309836 448196
rect 309048 444508 309100 444514
rect 309048 444450 309100 444456
rect 307956 442734 308338 442762
rect 309060 442748 309088 444450
rect 309796 442748 309824 448190
rect 310532 442762 310560 452066
rect 311912 442762 311940 478110
rect 322938 476912 322994 476921
rect 322938 476847 322994 476856
rect 313278 476504 313334 476513
rect 313278 476439 313280 476448
rect 313332 476439 313334 476448
rect 314658 476504 314714 476513
rect 314658 476439 314714 476448
rect 313280 476410 313332 476416
rect 314672 476406 314700 476439
rect 314660 476400 314712 476406
rect 314660 476342 314712 476348
rect 317418 476368 317474 476377
rect 317418 476303 317420 476312
rect 317472 476303 317474 476312
rect 320178 476368 320234 476377
rect 320178 476303 320234 476312
rect 317420 476274 317472 476280
rect 320192 476270 320220 476303
rect 320180 476264 320232 476270
rect 320180 476206 320232 476212
rect 322952 476202 322980 476847
rect 325790 476232 325846 476241
rect 322940 476196 322992 476202
rect 325790 476167 325846 476176
rect 322940 476138 322992 476144
rect 325804 476134 325832 476167
rect 325792 476128 325844 476134
rect 325792 476070 325844 476076
rect 332600 474768 332652 474774
rect 332600 474710 332652 474716
rect 316040 465724 316092 465730
rect 316040 465666 316092 465672
rect 316052 460934 316080 465666
rect 332612 460934 332640 474710
rect 353300 474020 353352 474026
rect 353300 473962 353352 473968
rect 333980 462392 334032 462398
rect 333980 462334 334032 462340
rect 333992 460934 334020 462334
rect 316052 460906 316448 460934
rect 332612 460906 333376 460934
rect 333992 460906 334848 460934
rect 313648 445528 313700 445534
rect 313648 445470 313700 445476
rect 312912 445120 312964 445126
rect 312912 445062 312964 445068
rect 310532 442734 310638 442762
rect 311912 442734 312202 442762
rect 312924 442748 312952 445062
rect 313660 442748 313688 445470
rect 314476 445188 314528 445194
rect 314476 445130 314528 445136
rect 314488 442748 314516 445130
rect 315212 445052 315264 445058
rect 315212 444994 315264 445000
rect 315224 442748 315252 444994
rect 315856 444984 315908 444990
rect 315856 444926 315908 444932
rect 315868 442542 315896 444926
rect 316420 442762 316448 460906
rect 330208 453756 330260 453762
rect 330208 453698 330260 453704
rect 320272 453688 320324 453694
rect 320272 453630 320324 453636
rect 317512 449336 317564 449342
rect 317512 449278 317564 449284
rect 316420 442734 316802 442762
rect 317524 442748 317552 449278
rect 319812 449268 319864 449274
rect 319812 449210 319864 449216
rect 319076 448180 319128 448186
rect 319076 448122 319128 448128
rect 318800 445052 318852 445058
rect 318800 444994 318852 445000
rect 304172 442536 304224 442542
rect 304172 442478 304224 442484
rect 315856 442536 315908 442542
rect 315856 442478 315908 442484
rect 318812 442474 318840 444994
rect 319088 442748 319116 448122
rect 319824 442748 319852 449210
rect 320284 442762 320312 453630
rect 329932 453620 329984 453626
rect 329932 453562 329984 453568
rect 327080 453552 327132 453558
rect 327080 453494 327132 453500
rect 327172 453552 327224 453558
rect 327172 453494 327224 453500
rect 322940 452260 322992 452266
rect 322940 452202 322992 452208
rect 321376 448044 321428 448050
rect 321376 447986 321428 447992
rect 320284 442734 320666 442762
rect 321388 442748 321416 447986
rect 322112 446412 322164 446418
rect 322112 446354 322164 446360
rect 321560 444508 321612 444514
rect 321560 444450 321612 444456
rect 321572 443698 321600 444450
rect 321560 443692 321612 443698
rect 321560 443634 321612 443640
rect 322124 442748 322152 446354
rect 322952 442748 322980 452202
rect 324504 450628 324556 450634
rect 324504 450570 324556 450576
rect 323676 447908 323728 447914
rect 323676 447850 323728 447856
rect 323688 442748 323716 447850
rect 324516 442748 324544 450570
rect 326804 450560 326856 450566
rect 326804 450502 326856 450508
rect 325792 449200 325844 449206
rect 325792 449142 325844 449148
rect 325240 446412 325292 446418
rect 325240 446354 325292 446360
rect 325252 442748 325280 446354
rect 325804 442762 325832 449142
rect 325976 443624 326028 443630
rect 325976 443566 326028 443572
rect 325988 443086 326016 443566
rect 325976 443080 326028 443086
rect 325976 443022 326028 443028
rect 325804 442734 326002 442762
rect 326816 442748 326844 450502
rect 327092 446758 327120 453494
rect 327080 446752 327132 446758
rect 327080 446694 327132 446700
rect 327184 442762 327212 453494
rect 329104 450696 329156 450702
rect 329104 450638 329156 450644
rect 327908 446752 327960 446758
rect 327908 446694 327960 446700
rect 327920 442762 327948 446694
rect 327184 442734 327566 442762
rect 327920 442734 328302 442762
rect 329116 442748 329144 450638
rect 329944 442762 329972 453562
rect 329866 442734 329972 442762
rect 330220 442762 330248 453698
rect 331220 451988 331272 451994
rect 331220 451930 331272 451936
rect 331232 442762 331260 451930
rect 332140 449200 332192 449206
rect 332140 449142 332192 449148
rect 330220 442734 330694 442762
rect 331232 442734 331430 442762
rect 332152 442748 332180 449142
rect 332968 447840 333020 447846
rect 332968 447782 333020 447788
rect 332980 442748 333008 447782
rect 333348 442762 333376 460906
rect 334440 446616 334492 446622
rect 334440 446558 334492 446564
rect 333348 442734 333730 442762
rect 334452 442748 334480 446558
rect 334820 442762 334848 460906
rect 336832 454912 336884 454918
rect 336832 454854 336884 454860
rect 336004 443624 336056 443630
rect 336004 443566 336056 443572
rect 334820 442734 335294 442762
rect 336016 442748 336044 443566
rect 336844 442748 336872 454854
rect 351920 453484 351972 453490
rect 351920 453426 351972 453432
rect 347872 452056 347924 452062
rect 347872 451998 347924 452004
rect 343732 446548 343784 446554
rect 343732 446490 343784 446496
rect 340972 445528 341024 445534
rect 340972 445470 341024 445476
rect 339132 445256 339184 445262
rect 339132 445198 339184 445204
rect 337568 444848 337620 444854
rect 337568 444790 337620 444796
rect 337580 442748 337608 444790
rect 338304 443148 338356 443154
rect 338304 443090 338356 443096
rect 338316 442748 338344 443090
rect 339144 442748 339172 445198
rect 339868 444780 339920 444786
rect 339868 444722 339920 444728
rect 339880 442748 339908 444722
rect 340880 444440 340932 444446
rect 340880 444382 340932 444388
rect 340696 443352 340748 443358
rect 340696 443294 340748 443300
rect 340708 442748 340736 443294
rect 318800 442468 318852 442474
rect 318800 442410 318852 442416
rect 311544 442338 311756 442354
rect 340892 442338 340920 444382
rect 340984 443766 341012 445470
rect 341432 445324 341484 445330
rect 341432 445266 341484 445272
rect 340972 443760 341024 443766
rect 340972 443702 341024 443708
rect 341444 442748 341472 445266
rect 342258 444680 342314 444689
rect 342258 444615 342314 444624
rect 342272 443834 342300 444615
rect 342260 443828 342312 443834
rect 342260 443770 342312 443776
rect 342168 443556 342220 443562
rect 342168 443498 342220 443504
rect 342180 442748 342208 443498
rect 342996 443420 343048 443426
rect 342996 443362 343048 443368
rect 343008 442748 343036 443362
rect 343744 442748 343772 446490
rect 346032 446480 346084 446486
rect 346032 446422 346084 446428
rect 345294 443184 345350 443193
rect 345294 443119 345350 443128
rect 344468 443012 344520 443018
rect 344468 442954 344520 442960
rect 344480 442748 344508 442954
rect 345308 442748 345336 443119
rect 346044 442748 346072 446422
rect 346860 444644 346912 444650
rect 346860 444586 346912 444592
rect 346872 442748 346900 444586
rect 347594 443048 347650 443057
rect 347594 442983 347650 442992
rect 347608 442748 347636 442983
rect 347884 442762 347912 451998
rect 350632 451920 350684 451926
rect 350632 451862 350684 451868
rect 349160 445460 349212 445466
rect 349160 445402 349212 445408
rect 347884 442734 348358 442762
rect 349172 442748 349200 445402
rect 349896 444576 349948 444582
rect 349896 444518 349948 444524
rect 349804 444508 349856 444514
rect 349804 444450 349856 444456
rect 311532 442332 311768 442338
rect 311584 442326 311716 442332
rect 311532 442274 311584 442280
rect 311716 442274 311768 442280
rect 340880 442332 340932 442338
rect 340880 442274 340932 442280
rect 349816 442270 349844 444450
rect 349908 442748 349936 444518
rect 350644 442748 350672 451862
rect 351932 446758 351960 453426
rect 352012 453416 352064 453422
rect 352012 453358 352064 453364
rect 351920 446752 351972 446758
rect 351920 446694 351972 446700
rect 351460 445392 351512 445398
rect 351460 445334 351512 445340
rect 351472 442748 351500 445334
rect 352024 442762 352052 453358
rect 353312 446758 353340 473962
rect 353392 453348 353444 453354
rect 353392 453290 353444 453296
rect 352748 446752 352800 446758
rect 352748 446694 352800 446700
rect 353300 446752 353352 446758
rect 353300 446694 353352 446700
rect 352760 442762 352788 446694
rect 353404 442762 353432 453290
rect 354220 446752 354272 446758
rect 354220 446694 354272 446700
rect 354232 442762 354260 446694
rect 355324 446684 355376 446690
rect 355324 446626 355376 446632
rect 352024 442734 352222 442762
rect 352760 442734 353050 442762
rect 353404 442734 353786 442762
rect 354232 442734 354522 442762
rect 355336 442748 355364 446626
rect 357452 445194 357480 700334
rect 357544 478174 357572 700470
rect 358912 700460 358964 700466
rect 358912 700402 358964 700408
rect 361028 700460 361080 700466
rect 361028 700402 361080 700408
rect 358820 700324 358872 700330
rect 358820 700266 358872 700272
rect 358084 616888 358136 616894
rect 358084 616830 358136 616836
rect 357532 478168 357584 478174
rect 357532 478110 357584 478116
rect 358096 449478 358124 616830
rect 358176 536852 358228 536858
rect 358176 536794 358228 536800
rect 358188 452266 358216 536794
rect 358268 484424 358320 484430
rect 358268 484366 358320 484372
rect 358280 453694 358308 484366
rect 358268 453688 358320 453694
rect 358268 453630 358320 453636
rect 358176 452260 358228 452266
rect 358176 452202 358228 452208
rect 358084 449472 358136 449478
rect 358084 449414 358136 449420
rect 358832 445330 358860 700266
rect 358820 445324 358872 445330
rect 358820 445266 358872 445272
rect 357440 445188 357492 445194
rect 357440 445130 357492 445136
rect 358924 445126 358952 700402
rect 360936 700392 360988 700398
rect 360936 700334 360988 700340
rect 360844 700324 360896 700330
rect 360844 700266 360896 700272
rect 359464 670744 359516 670750
rect 359464 670686 359516 670692
rect 359004 565140 359056 565146
rect 359004 565082 359056 565088
rect 359016 445262 359044 565082
rect 359476 450838 359504 670686
rect 360856 450906 360884 700266
rect 360948 452198 360976 700334
rect 361040 454918 361068 700402
rect 362224 696992 362276 696998
rect 362224 696934 362276 696940
rect 361120 643136 361172 643142
rect 361120 643078 361172 643084
rect 361028 454912 361080 454918
rect 361028 454854 361080 454860
rect 361132 453558 361160 643078
rect 362236 453626 362264 696934
rect 362224 453620 362276 453626
rect 362224 453562 362276 453568
rect 361120 453552 361172 453558
rect 361120 453494 361172 453500
rect 360936 452192 360988 452198
rect 360936 452134 360988 452140
rect 364352 452130 364380 702406
rect 397472 700466 397500 703520
rect 397460 700460 397512 700466
rect 397460 700402 397512 700408
rect 371884 563100 371936 563106
rect 371884 563042 371936 563048
rect 364340 452124 364392 452130
rect 364340 452066 364392 452072
rect 360844 450900 360896 450906
rect 360844 450842 360896 450848
rect 359464 450832 359516 450838
rect 359464 450774 359516 450780
rect 371896 449410 371924 563042
rect 371884 449404 371936 449410
rect 371884 449346 371936 449352
rect 412652 448254 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700398 429884 703520
rect 429844 700392 429896 700398
rect 429844 700334 429896 700340
rect 412640 448248 412692 448254
rect 412640 448190 412692 448196
rect 462332 446622 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 448118 477540 702406
rect 494072 450770 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 450764 494112 450770
rect 494060 450706 494112 450712
rect 527192 449206 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 449200 527232 449206
rect 527180 449142 527232 449148
rect 477500 448112 477552 448118
rect 477500 448054 477552 448060
rect 542372 447982 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 579618 537840 579674 537849
rect 579618 537775 579674 537784
rect 579632 536858 579660 537775
rect 579620 536852 579672 536858
rect 579620 536794 579672 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 454850 580304 683839
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580264 454844 580316 454850
rect 580264 454786 580316 454792
rect 580368 454782 580396 630799
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580356 454776 580408 454782
rect 580356 454718 580408 454724
rect 542360 447976 542412 447982
rect 542360 447918 542412 447924
rect 462320 446616 462372 446622
rect 462320 446558 462372 446564
rect 580460 446418 580488 590951
rect 580538 577688 580594 577697
rect 580538 577623 580594 577632
rect 580552 454714 580580 577623
rect 580540 454708 580592 454714
rect 580540 454650 580592 454656
rect 580448 446412 580500 446418
rect 580448 446354 580500 446360
rect 359004 445256 359056 445262
rect 359004 445198 359056 445204
rect 358912 445120 358964 445126
rect 358912 445062 358964 445068
rect 356796 445052 356848 445058
rect 356796 444994 356848 445000
rect 356060 443488 356112 443494
rect 356060 443430 356112 443436
rect 356072 442748 356100 443430
rect 356808 442748 356836 444994
rect 358360 444984 358412 444990
rect 358360 444926 358412 444932
rect 357624 444440 357676 444446
rect 357624 444382 357676 444388
rect 357636 442748 357664 444382
rect 358372 442748 358400 444926
rect 359924 444916 359976 444922
rect 359924 444858 359976 444864
rect 359188 444508 359240 444514
rect 359188 444450 359240 444456
rect 359200 442748 359228 444450
rect 359936 442748 359964 444858
rect 538862 444816 538918 444825
rect 538862 444751 538918 444760
rect 360660 444712 360712 444718
rect 360660 444654 360712 444660
rect 360672 442748 360700 444654
rect 312084 442264 312136 442270
rect 307022 442232 307078 442241
rect 306774 442190 307022 442218
rect 311374 442212 312084 442218
rect 316040 442264 316092 442270
rect 311374 442206 312136 442212
rect 315974 442212 316040 442218
rect 318524 442264 318576 442270
rect 315974 442206 316092 442212
rect 318366 442212 318524 442218
rect 318366 442206 318576 442212
rect 349804 442264 349856 442270
rect 349804 442206 349856 442212
rect 361210 442232 361266 442241
rect 311374 442190 312124 442206
rect 315974 442190 316080 442206
rect 318366 442190 318564 442206
rect 307022 442167 307078 442176
rect 361946 442232 362002 442241
rect 361266 442190 361514 442218
rect 361210 442167 361266 442176
rect 362002 442190 362250 442218
rect 361946 442167 362002 442176
rect 304448 442128 304500 442134
rect 304448 442070 304500 442076
rect 304460 442068 304488 442070
rect 363696 441856 363748 441862
rect 363696 441798 363748 441804
rect 363604 441788 363656 441794
rect 363604 441730 363656 441736
rect 232240 412606 232360 412634
rect 232240 411262 232268 412606
rect 232228 411256 232280 411262
rect 232228 411198 232280 411204
rect 231308 398812 231360 398818
rect 231308 398754 231360 398760
rect 363616 379506 363644 441730
rect 363708 431934 363736 441798
rect 364984 441720 365036 441726
rect 364984 441662 365036 441668
rect 363696 431928 363748 431934
rect 363696 431870 363748 431876
rect 363604 379500 363656 379506
rect 363604 379442 363656 379448
rect 231216 358760 231268 358766
rect 231216 358702 231268 358708
rect 309258 310554 309456 310570
rect 310638 310554 310836 310570
rect 309258 310548 309468 310554
rect 309258 310542 309416 310548
rect 309416 310490 309468 310496
rect 309784 310548 309836 310554
rect 310638 310548 310848 310554
rect 310638 310542 310796 310548
rect 309784 310490 309836 310496
rect 310796 310490 310848 310496
rect 311164 310548 311216 310554
rect 311164 310490 311216 310496
rect 231872 310406 232530 310434
rect 231768 308440 231820 308446
rect 231768 308382 231820 308388
rect 231780 308106 231808 308382
rect 231768 308100 231820 308106
rect 231768 308042 231820 308048
rect 231124 306332 231176 306338
rect 231124 306274 231176 306280
rect 219348 300008 219400 300014
rect 219348 299950 219400 299956
rect 219256 245404 219308 245410
rect 219256 245346 219308 245352
rect 219164 243704 219216 243710
rect 219164 243646 219216 243652
rect 219072 158568 219124 158574
rect 219072 158510 219124 158516
rect 218888 158024 218940 158030
rect 218888 157966 218940 157972
rect 218796 155644 218848 155650
rect 218796 155586 218848 155592
rect 218704 155372 218756 155378
rect 218704 155314 218756 155320
rect 218612 155168 218664 155174
rect 218612 155110 218664 155116
rect 218072 16546 219112 16574
rect 218794 4040 218850 4049
rect 218794 3975 218850 3984
rect 218808 3641 218836 3975
rect 218794 3632 218850 3641
rect 218794 3567 218850 3576
rect 217416 3528 217468 3534
rect 217416 3470 217468 3476
rect 218058 3496 218114 3505
rect 219084 3482 219112 16546
rect 219176 3806 219204 243646
rect 219164 3800 219216 3806
rect 219164 3742 219216 3748
rect 219268 3618 219296 245346
rect 219360 3738 219388 299950
rect 231872 258738 231900 310406
rect 231952 308440 232004 308446
rect 232700 308394 232728 310420
rect 232884 308446 232912 310420
rect 232976 310406 233174 310434
rect 231952 308382 232004 308388
rect 231860 258732 231912 258738
rect 231860 258674 231912 258680
rect 231964 245002 231992 308382
rect 232056 308366 232728 308394
rect 232872 308440 232924 308446
rect 232872 308382 232924 308388
rect 231952 244996 232004 245002
rect 231952 244938 232004 244944
rect 232056 244934 232084 308366
rect 232976 296714 233004 310406
rect 233344 308632 233372 310420
rect 233252 308604 233372 308632
rect 233436 310406 233634 310434
rect 233148 308508 233200 308514
rect 233148 308450 233200 308456
rect 233160 308038 233188 308450
rect 233252 308417 233280 308604
rect 233332 308508 233384 308514
rect 233332 308450 233384 308456
rect 233238 308408 233294 308417
rect 233238 308343 233294 308352
rect 233148 308032 233200 308038
rect 233148 307974 233200 307980
rect 232148 296686 233004 296714
rect 232148 264246 232176 296686
rect 232136 264240 232188 264246
rect 232136 264182 232188 264188
rect 233344 253230 233372 308450
rect 233436 256018 233464 310406
rect 233516 308440 233568 308446
rect 233516 308382 233568 308388
rect 233528 267034 233556 308382
rect 233804 296714 233832 310420
rect 233896 310406 234094 310434
rect 233896 308446 233924 310406
rect 234264 308514 234292 310420
rect 234540 308582 234568 310420
rect 234528 308576 234580 308582
rect 234528 308518 234580 308524
rect 234252 308508 234304 308514
rect 234252 308450 234304 308456
rect 233884 308440 233936 308446
rect 233884 308382 233936 308388
rect 234724 306320 234752 310420
rect 233712 296686 233832 296714
rect 234632 306292 234752 306320
rect 234816 310406 235014 310434
rect 233516 267028 233568 267034
rect 233516 266970 233568 266976
rect 233424 256012 233476 256018
rect 233424 255954 233476 255960
rect 233332 253224 233384 253230
rect 233332 253166 233384 253172
rect 233712 246362 233740 296686
rect 234632 246430 234660 306292
rect 234712 305380 234764 305386
rect 234712 305322 234764 305328
rect 234724 250510 234752 305322
rect 234816 251870 234844 310406
rect 235184 306882 235212 310420
rect 235276 310406 235474 310434
rect 235172 306876 235224 306882
rect 235172 306818 235224 306824
rect 235080 306672 235132 306678
rect 235080 306614 235132 306620
rect 234896 306332 234948 306338
rect 234896 306274 234948 306280
rect 234908 253298 234936 306274
rect 234988 302252 235040 302258
rect 234988 302194 235040 302200
rect 235000 256086 235028 302194
rect 235092 269822 235120 306614
rect 235276 302258 235304 310406
rect 235644 305386 235672 310420
rect 235736 310406 235934 310434
rect 235736 306338 235764 310406
rect 236104 308106 236132 310420
rect 236380 308718 236408 310420
rect 236368 308712 236420 308718
rect 236368 308654 236420 308660
rect 236092 308100 236144 308106
rect 236092 308042 236144 308048
rect 236092 306468 236144 306474
rect 236092 306410 236144 306416
rect 235724 306332 235776 306338
rect 235724 306274 235776 306280
rect 235632 305380 235684 305386
rect 235632 305322 235684 305328
rect 235264 302252 235316 302258
rect 235264 302194 235316 302200
rect 235080 269816 235132 269822
rect 235080 269758 235132 269764
rect 236104 256154 236132 306410
rect 236276 306400 236328 306406
rect 236276 306342 236328 306348
rect 236184 306332 236236 306338
rect 236184 306274 236236 306280
rect 236196 271182 236224 306274
rect 236288 276690 236316 306342
rect 236564 296714 236592 310420
rect 236656 310406 236854 310434
rect 236656 306338 236684 310406
rect 237024 306406 237052 310420
rect 237116 310406 237314 310434
rect 237116 306474 237144 310406
rect 237104 306468 237156 306474
rect 237104 306410 237156 306416
rect 237012 306400 237064 306406
rect 237012 306342 237064 306348
rect 236644 306332 236696 306338
rect 236644 306274 236696 306280
rect 236380 296686 236592 296714
rect 236276 276684 236328 276690
rect 236276 276626 236328 276632
rect 236184 271176 236236 271182
rect 236184 271118 236236 271124
rect 236092 256148 236144 256154
rect 236092 256090 236144 256096
rect 234988 256080 235040 256086
rect 234988 256022 235040 256028
rect 234896 253292 234948 253298
rect 234896 253234 234948 253240
rect 236380 251938 236408 296686
rect 237484 252006 237512 310420
rect 237576 310406 237774 310434
rect 237576 272542 237604 310406
rect 237944 308038 237972 310420
rect 238036 310406 238234 310434
rect 237932 308032 237984 308038
rect 237932 307974 237984 307980
rect 237748 306400 237800 306406
rect 237748 306342 237800 306348
rect 237656 306332 237708 306338
rect 237656 306274 237708 306280
rect 237668 273970 237696 306274
rect 237760 283626 237788 306342
rect 238036 296714 238064 310406
rect 238404 306338 238432 310420
rect 238496 310406 238694 310434
rect 238496 306406 238524 310406
rect 238484 306400 238536 306406
rect 238484 306342 238536 306348
rect 238392 306332 238444 306338
rect 238392 306274 238444 306280
rect 237852 296686 238064 296714
rect 237748 283620 237800 283626
rect 237748 283562 237800 283568
rect 237656 273964 237708 273970
rect 237656 273906 237708 273912
rect 237564 272536 237616 272542
rect 237564 272478 237616 272484
rect 237852 252074 237880 296686
rect 238864 258806 238892 310420
rect 239048 310406 239154 310434
rect 238944 306332 238996 306338
rect 238944 306274 238996 306280
rect 238956 260166 238984 306274
rect 239048 280838 239076 310406
rect 239324 308650 239352 310420
rect 239416 310406 239614 310434
rect 239312 308644 239364 308650
rect 239312 308586 239364 308592
rect 239128 306400 239180 306406
rect 239128 306342 239180 306348
rect 239140 287706 239168 306342
rect 239416 306338 239444 310406
rect 239404 306332 239456 306338
rect 239404 306274 239456 306280
rect 239784 296714 239812 310420
rect 239968 306406 239996 310420
rect 239956 306400 240008 306406
rect 239956 306342 240008 306348
rect 240244 306320 240272 310420
rect 240442 310406 240548 310434
rect 240416 306332 240468 306338
rect 240244 306292 240364 306320
rect 240232 305380 240284 305386
rect 240232 305322 240284 305328
rect 239232 296686 239812 296714
rect 239128 287700 239180 287706
rect 239128 287642 239180 287648
rect 239036 280832 239088 280838
rect 239036 280774 239088 280780
rect 238944 260160 238996 260166
rect 238944 260102 238996 260108
rect 238852 258800 238904 258806
rect 238852 258742 238904 258748
rect 239232 254590 239260 296686
rect 240244 254862 240272 305322
rect 240336 262886 240364 306292
rect 240416 306274 240468 306280
rect 240428 265674 240456 306274
rect 240520 282198 240548 310406
rect 240704 308786 240732 310420
rect 240692 308780 240744 308786
rect 240692 308722 240744 308728
rect 240888 306338 240916 310420
rect 240980 310406 241178 310434
rect 240876 306332 240928 306338
rect 240876 306274 240928 306280
rect 240980 296714 241008 310406
rect 241348 305386 241376 310420
rect 241336 305380 241388 305386
rect 241336 305322 241388 305328
rect 241520 305108 241572 305114
rect 241520 305050 241572 305056
rect 240612 296686 241008 296714
rect 240508 282192 240560 282198
rect 240508 282134 240560 282140
rect 240416 265668 240468 265674
rect 240416 265610 240468 265616
rect 240324 262880 240376 262886
rect 240324 262822 240376 262828
rect 240232 254856 240284 254862
rect 240232 254798 240284 254804
rect 240612 254658 240640 296686
rect 240600 254652 240652 254658
rect 240600 254594 240652 254600
rect 239220 254584 239272 254590
rect 239220 254526 239272 254532
rect 237840 252068 237892 252074
rect 237840 252010 237892 252016
rect 237472 252000 237524 252006
rect 237472 251942 237524 251948
rect 236368 251932 236420 251938
rect 236368 251874 236420 251880
rect 234804 251864 234856 251870
rect 234804 251806 234856 251812
rect 234712 250504 234764 250510
rect 234712 250446 234764 250452
rect 241532 246566 241560 305050
rect 241520 246560 241572 246566
rect 241520 246502 241572 246508
rect 241624 246498 241652 310420
rect 241808 306320 241836 310420
rect 241716 306292 241836 306320
rect 241900 310406 242098 310434
rect 241716 267102 241744 306292
rect 241796 305380 241848 305386
rect 241796 305322 241848 305328
rect 241808 268394 241836 305322
rect 241900 284986 241928 310406
rect 242268 305114 242296 310420
rect 242360 310406 242558 310434
rect 242360 305386 242388 310406
rect 242348 305380 242400 305386
rect 242348 305322 242400 305328
rect 242256 305108 242308 305114
rect 242256 305050 242308 305056
rect 242728 296714 242756 310420
rect 241992 296686 242756 296714
rect 242912 310406 243018 310434
rect 243202 310406 243308 310434
rect 241992 286346 242020 296686
rect 241980 286340 242032 286346
rect 241980 286282 242032 286288
rect 241888 284980 241940 284986
rect 241888 284922 241940 284928
rect 241796 268388 241848 268394
rect 241796 268330 241848 268336
rect 241704 267096 241756 267102
rect 241704 267038 241756 267044
rect 242912 247722 242940 310406
rect 243280 306474 243308 310406
rect 243372 310406 243478 310434
rect 243268 306468 243320 306474
rect 243268 306410 243320 306416
rect 243084 306400 243136 306406
rect 243084 306342 243136 306348
rect 242992 306332 243044 306338
rect 242992 306274 243044 306280
rect 243004 249082 243032 306274
rect 243096 254794 243124 306342
rect 243372 302682 243400 310406
rect 243452 306468 243504 306474
rect 243452 306410 243504 306416
rect 243188 302654 243400 302682
rect 243084 254788 243136 254794
rect 243084 254730 243136 254736
rect 243188 254726 243216 302654
rect 243464 299474 243492 306410
rect 243648 306338 243676 310420
rect 243740 310406 243938 310434
rect 243636 306332 243688 306338
rect 243636 306274 243688 306280
rect 243280 299446 243492 299474
rect 243280 275330 243308 299446
rect 243740 296714 243768 310406
rect 244108 306406 244136 310420
rect 244096 306400 244148 306406
rect 244096 306342 244148 306348
rect 244384 306338 244412 310420
rect 244568 306354 244596 310420
rect 244372 306332 244424 306338
rect 244372 306274 244424 306280
rect 244476 306326 244596 306354
rect 244660 310406 244858 310434
rect 244372 305312 244424 305318
rect 244372 305254 244424 305260
rect 243372 296686 243768 296714
rect 243372 276826 243400 296686
rect 243360 276820 243412 276826
rect 243360 276762 243412 276768
rect 243268 275324 243320 275330
rect 243268 275266 243320 275272
rect 244384 260234 244412 305254
rect 244476 276758 244504 306326
rect 244556 305380 244608 305386
rect 244556 305322 244608 305328
rect 244568 278050 244596 305322
rect 244660 287774 244688 310406
rect 244740 306332 244792 306338
rect 244740 306274 244792 306280
rect 244648 287768 244700 287774
rect 244648 287710 244700 287716
rect 244556 278044 244608 278050
rect 244556 277986 244608 277992
rect 244464 276752 244516 276758
rect 244464 276694 244516 276700
rect 244372 260228 244424 260234
rect 244372 260170 244424 260176
rect 244752 258874 244780 306274
rect 245028 305318 245056 310420
rect 245120 310406 245318 310434
rect 245120 305386 245148 310406
rect 245488 307086 245516 310420
rect 245476 307080 245528 307086
rect 245476 307022 245528 307028
rect 245660 306332 245712 306338
rect 245660 306274 245712 306280
rect 245108 305380 245160 305386
rect 245108 305322 245160 305328
rect 245016 305312 245068 305318
rect 245016 305254 245068 305260
rect 244740 258868 244792 258874
rect 244740 258810 244792 258816
rect 243176 254720 243228 254726
rect 243176 254662 243228 254668
rect 245672 250578 245700 306274
rect 245764 258942 245792 310420
rect 245948 306354 245976 310420
rect 245856 306326 245976 306354
rect 246040 310406 246238 310434
rect 245856 279478 245884 306326
rect 245936 305380 245988 305386
rect 245936 305322 245988 305328
rect 245948 282266 245976 305322
rect 246040 289134 246068 310406
rect 246408 306338 246436 310420
rect 246500 310406 246698 310434
rect 246396 306332 246448 306338
rect 246396 306274 246448 306280
rect 246500 305386 246528 310406
rect 246488 305380 246540 305386
rect 246488 305322 246540 305328
rect 246868 296714 246896 310420
rect 246132 296686 246896 296714
rect 246132 290494 246160 296686
rect 246120 290488 246172 290494
rect 246120 290430 246172 290436
rect 246028 289128 246080 289134
rect 246028 289070 246080 289076
rect 245936 282260 245988 282266
rect 245936 282202 245988 282208
rect 245844 279472 245896 279478
rect 245844 279414 245896 279420
rect 245752 258936 245804 258942
rect 245752 258878 245804 258884
rect 247052 250646 247080 310420
rect 247224 306468 247276 306474
rect 247224 306410 247276 306416
rect 247132 306400 247184 306406
rect 247132 306342 247184 306348
rect 247144 250714 247172 306342
rect 247236 253366 247264 306410
rect 247328 283694 247356 310420
rect 247408 306332 247460 306338
rect 247408 306274 247460 306280
rect 247420 290630 247448 306274
rect 247408 290624 247460 290630
rect 247408 290566 247460 290572
rect 247512 290562 247540 310420
rect 247604 310406 247802 310434
rect 247604 306406 247632 310406
rect 247972 306474 248000 310420
rect 248064 310406 248262 310434
rect 248446 310406 248644 310434
rect 247960 306468 248012 306474
rect 247960 306410 248012 306416
rect 247592 306400 247644 306406
rect 247592 306342 247644 306348
rect 248064 306338 248092 310406
rect 248616 306746 248644 310406
rect 248604 306740 248656 306746
rect 248604 306682 248656 306688
rect 248604 306536 248656 306542
rect 248604 306478 248656 306484
rect 248512 306400 248564 306406
rect 248512 306342 248564 306348
rect 248052 306332 248104 306338
rect 248052 306274 248104 306280
rect 248420 306332 248472 306338
rect 248420 306274 248472 306280
rect 248432 291854 248460 306274
rect 248420 291848 248472 291854
rect 248420 291790 248472 291796
rect 247500 290556 247552 290562
rect 247500 290498 247552 290504
rect 247316 283688 247368 283694
rect 247316 283630 247368 283636
rect 248524 253434 248552 306342
rect 248616 261526 248644 306478
rect 248708 306406 248736 310420
rect 248696 306400 248748 306406
rect 248696 306342 248748 306348
rect 248696 305380 248748 305386
rect 248696 305322 248748 305328
rect 248708 264314 248736 305322
rect 248892 302234 248920 310420
rect 248984 310406 249182 310434
rect 248984 305386 249012 310406
rect 248972 305380 249024 305386
rect 248972 305322 249024 305328
rect 248800 302206 248920 302234
rect 248800 290698 248828 302206
rect 249352 296714 249380 310420
rect 249444 310406 249642 310434
rect 249444 306338 249472 310406
rect 249708 306672 249760 306678
rect 249708 306614 249760 306620
rect 249432 306332 249484 306338
rect 249432 306274 249484 306280
rect 249720 305266 249748 306614
rect 249812 305386 249840 310420
rect 249996 310406 250102 310434
rect 249892 306604 249944 306610
rect 249892 306546 249944 306552
rect 249800 305380 249852 305386
rect 249800 305322 249852 305328
rect 249720 305238 249840 305266
rect 248892 296686 249380 296714
rect 248788 290692 248840 290698
rect 248788 290634 248840 290640
rect 248696 264308 248748 264314
rect 248696 264250 248748 264256
rect 248604 261520 248656 261526
rect 248604 261462 248656 261468
rect 248892 253502 248920 296686
rect 249812 291922 249840 305238
rect 249800 291916 249852 291922
rect 249800 291858 249852 291864
rect 249904 271250 249932 306546
rect 249996 285054 250024 310406
rect 250272 306678 250300 310420
rect 250364 310406 250562 310434
rect 250260 306672 250312 306678
rect 250260 306614 250312 306620
rect 250364 306610 250392 310406
rect 250352 306604 250404 306610
rect 250352 306546 250404 306552
rect 250732 306490 250760 310420
rect 250088 306462 250760 306490
rect 250824 310406 251022 310434
rect 251206 310406 251312 310434
rect 250088 286414 250116 306462
rect 250824 306354 250852 310406
rect 250180 306326 250852 306354
rect 251180 306400 251232 306406
rect 251180 306342 251232 306348
rect 250180 291990 250208 306326
rect 250260 305380 250312 305386
rect 250260 305322 250312 305328
rect 250168 291984 250220 291990
rect 250168 291926 250220 291932
rect 250076 286408 250128 286414
rect 250076 286350 250128 286356
rect 249984 285048 250036 285054
rect 249984 284990 250036 284996
rect 249892 271244 249944 271250
rect 249892 271186 249944 271192
rect 250272 269890 250300 305322
rect 251192 293282 251220 306342
rect 251180 293276 251232 293282
rect 251180 293218 251232 293224
rect 251284 282334 251312 310406
rect 251468 306354 251496 310420
rect 251364 306332 251416 306338
rect 251468 306326 251588 306354
rect 251364 306274 251416 306280
rect 251376 283762 251404 306274
rect 251456 305380 251508 305386
rect 251456 305322 251508 305328
rect 251468 286550 251496 305322
rect 251456 286544 251508 286550
rect 251456 286486 251508 286492
rect 251560 286482 251588 306326
rect 251548 286476 251600 286482
rect 251548 286418 251600 286424
rect 251364 283756 251416 283762
rect 251364 283698 251416 283704
rect 251272 282328 251324 282334
rect 251272 282270 251324 282276
rect 250260 269884 250312 269890
rect 250260 269826 250312 269832
rect 248880 253496 248932 253502
rect 248880 253438 248932 253444
rect 248512 253428 248564 253434
rect 248512 253370 248564 253376
rect 247224 253360 247276 253366
rect 247224 253302 247276 253308
rect 251652 250782 251680 310420
rect 251744 310406 251942 310434
rect 251744 306338 251772 310406
rect 251732 306332 251784 306338
rect 251732 306274 251784 306280
rect 252112 305386 252140 310420
rect 252204 310406 252402 310434
rect 252586 310406 252692 310434
rect 252204 306406 252232 310406
rect 252192 306400 252244 306406
rect 252192 306342 252244 306348
rect 252100 305380 252152 305386
rect 252100 305322 252152 305328
rect 252664 283830 252692 310406
rect 252744 306400 252796 306406
rect 252744 306342 252796 306348
rect 252756 287910 252784 306342
rect 252744 287904 252796 287910
rect 252744 287846 252796 287852
rect 252848 287842 252876 310420
rect 253032 308854 253060 310420
rect 253124 310406 253322 310434
rect 253020 308848 253072 308854
rect 253020 308790 253072 308796
rect 252928 306332 252980 306338
rect 252928 306274 252980 306280
rect 252940 293350 252968 306274
rect 253124 296714 253152 310406
rect 253204 307896 253256 307902
rect 253204 307838 253256 307844
rect 253032 296686 253152 296714
rect 252928 293344 252980 293350
rect 252928 293286 252980 293292
rect 252836 287836 252888 287842
rect 252836 287778 252888 287784
rect 253032 283898 253060 296686
rect 253020 283892 253072 283898
rect 253020 283834 253072 283840
rect 252652 283824 252704 283830
rect 252652 283766 252704 283772
rect 253216 262954 253244 307838
rect 253492 306406 253520 310420
rect 253584 310406 253782 310434
rect 253966 310406 254072 310434
rect 253480 306400 253532 306406
rect 253480 306342 253532 306348
rect 253584 306338 253612 310406
rect 253572 306332 253624 306338
rect 253572 306274 253624 306280
rect 254044 285122 254072 310406
rect 254136 310406 254242 310434
rect 254136 287978 254164 310406
rect 254412 308990 254440 310420
rect 254400 308984 254452 308990
rect 254400 308926 254452 308932
rect 254216 306400 254268 306406
rect 254596 306354 254624 310420
rect 254688 310406 254886 310434
rect 254688 306406 254716 310406
rect 254768 307828 254820 307834
rect 254768 307770 254820 307776
rect 254216 306342 254268 306348
rect 254228 289202 254256 306342
rect 254308 306332 254360 306338
rect 254308 306274 254360 306280
rect 254412 306326 254624 306354
rect 254676 306400 254728 306406
rect 254676 306342 254728 306348
rect 254320 293418 254348 306274
rect 254308 293412 254360 293418
rect 254308 293354 254360 293360
rect 254216 289196 254268 289202
rect 254216 289138 254268 289144
rect 254124 287972 254176 287978
rect 254124 287914 254176 287920
rect 254412 285190 254440 306326
rect 254780 302234 254808 307770
rect 255056 306338 255084 310420
rect 255044 306332 255096 306338
rect 255044 306274 255096 306280
rect 254596 302206 254808 302234
rect 255332 302234 255360 310420
rect 255332 302206 255452 302234
rect 254400 285184 254452 285190
rect 254400 285126 254452 285132
rect 254032 285116 254084 285122
rect 254032 285058 254084 285064
rect 253204 262948 253256 262954
rect 253204 262890 253256 262896
rect 251640 250776 251692 250782
rect 251640 250718 251692 250724
rect 247132 250708 247184 250714
rect 247132 250650 247184 250656
rect 247040 250640 247092 250646
rect 247040 250582 247092 250588
rect 245660 250572 245712 250578
rect 245660 250514 245712 250520
rect 242992 249076 243044 249082
rect 242992 249018 243044 249024
rect 242900 247716 242952 247722
rect 242900 247658 242952 247664
rect 241612 246492 241664 246498
rect 241612 246434 241664 246440
rect 234620 246424 234672 246430
rect 234620 246366 234672 246372
rect 233700 246356 233752 246362
rect 233700 246298 233752 246304
rect 254596 245138 254624 302206
rect 255424 285258 255452 302206
rect 255516 289270 255544 310420
rect 255792 309058 255820 310420
rect 255780 309052 255832 309058
rect 255780 308994 255832 309000
rect 255688 306400 255740 306406
rect 255688 306342 255740 306348
rect 255596 306332 255648 306338
rect 255596 306274 255648 306280
rect 255608 289338 255636 306274
rect 255700 294642 255728 306342
rect 255976 296714 256004 310420
rect 256068 310406 256266 310434
rect 256068 306338 256096 310406
rect 256436 306406 256464 310420
rect 256424 306400 256476 306406
rect 256424 306342 256476 306348
rect 256056 306332 256108 306338
rect 256712 306320 256740 310420
rect 256910 310406 257016 310434
rect 256712 306292 256924 306320
rect 256056 306274 256108 306280
rect 256700 305380 256752 305386
rect 256700 305322 256752 305328
rect 255792 296686 256004 296714
rect 255688 294636 255740 294642
rect 255688 294578 255740 294584
rect 255596 289332 255648 289338
rect 255596 289274 255648 289280
rect 255504 289264 255556 289270
rect 255504 289206 255556 289212
rect 255412 285252 255464 285258
rect 255412 285194 255464 285200
rect 255792 252142 255820 296686
rect 255780 252136 255832 252142
rect 255780 252078 255832 252084
rect 254584 245132 254636 245138
rect 254584 245074 254636 245080
rect 256712 245070 256740 305322
rect 256792 303748 256844 303754
rect 256792 303690 256844 303696
rect 256804 247790 256832 303690
rect 256896 260302 256924 306292
rect 256988 303226 257016 310406
rect 257172 303754 257200 310420
rect 257160 303748 257212 303754
rect 257160 303690 257212 303696
rect 256988 303198 257108 303226
rect 256976 303000 257028 303006
rect 256976 302942 257028 302948
rect 256988 261594 257016 302942
rect 257080 265742 257108 303198
rect 257356 303006 257384 310420
rect 257448 310406 257646 310434
rect 257448 305386 257476 310406
rect 257436 305380 257488 305386
rect 257436 305322 257488 305328
rect 257344 303000 257396 303006
rect 257344 302942 257396 302948
rect 257816 296714 257844 310420
rect 258092 307902 258120 310420
rect 258080 307896 258132 307902
rect 258080 307838 258132 307844
rect 258276 306320 258304 310420
rect 258460 310406 258566 310434
rect 257172 296686 257844 296714
rect 258184 306292 258304 306320
rect 258356 306332 258408 306338
rect 257172 272610 257200 296686
rect 257160 272604 257212 272610
rect 257160 272546 257212 272552
rect 258184 268462 258212 306292
rect 258356 306274 258408 306280
rect 258264 305380 258316 305386
rect 258264 305322 258316 305328
rect 258276 269958 258304 305322
rect 258368 274038 258396 306274
rect 258356 274032 258408 274038
rect 258356 273974 258408 273980
rect 258264 269952 258316 269958
rect 258264 269894 258316 269900
rect 258172 268456 258224 268462
rect 258172 268398 258224 268404
rect 257068 265736 257120 265742
rect 257068 265678 257120 265684
rect 256976 261588 257028 261594
rect 256976 261530 257028 261536
rect 256884 260296 256936 260302
rect 256884 260238 256936 260244
rect 258460 249150 258488 310406
rect 258736 307834 258764 310420
rect 258828 310406 259026 310434
rect 258724 307828 258776 307834
rect 258724 307770 258776 307776
rect 258828 305386 258856 310406
rect 259196 306338 259224 310420
rect 259472 306626 259500 310420
rect 259670 310406 259776 310434
rect 259472 306598 259684 306626
rect 259552 306468 259604 306474
rect 259552 306410 259604 306416
rect 259184 306332 259236 306338
rect 259184 306274 259236 306280
rect 258816 305380 258868 305386
rect 258816 305322 258868 305328
rect 259460 305380 259512 305386
rect 259460 305322 259512 305328
rect 258448 249144 258500 249150
rect 258448 249086 258500 249092
rect 256792 247784 256844 247790
rect 256792 247726 256844 247732
rect 259472 245206 259500 305322
rect 259564 247858 259592 306410
rect 259656 264382 259684 306598
rect 259748 271318 259776 310406
rect 259840 310406 259946 310434
rect 259840 278118 259868 310406
rect 260116 305386 260144 310420
rect 260208 310406 260406 310434
rect 260208 306474 260236 310406
rect 260196 306468 260248 306474
rect 260196 306410 260248 306416
rect 260104 305380 260156 305386
rect 260104 305322 260156 305328
rect 260576 305266 260604 310420
rect 260656 307828 260708 307834
rect 260656 307770 260708 307776
rect 259932 305238 260604 305266
rect 259932 279546 259960 305238
rect 260668 302234 260696 307770
rect 260852 305386 260880 310420
rect 261036 306320 261064 310420
rect 260944 306292 261064 306320
rect 261220 310406 261326 310434
rect 260840 305380 260892 305386
rect 260840 305322 260892 305328
rect 260840 305244 260892 305250
rect 260840 305186 260892 305192
rect 260116 302206 260696 302234
rect 259920 279540 259972 279546
rect 259920 279482 259972 279488
rect 259828 278112 259880 278118
rect 259828 278054 259880 278060
rect 259736 271312 259788 271318
rect 259736 271254 259788 271260
rect 259644 264376 259696 264382
rect 259644 264318 259696 264324
rect 260116 261662 260144 302206
rect 260104 261656 260156 261662
rect 260104 261598 260156 261604
rect 260852 247994 260880 305186
rect 260840 247988 260892 247994
rect 260840 247930 260892 247936
rect 260944 247926 260972 306292
rect 261220 305538 261248 310406
rect 261220 305510 261340 305538
rect 261024 305380 261076 305386
rect 261024 305322 261076 305328
rect 261208 305380 261260 305386
rect 261208 305322 261260 305328
rect 261036 265810 261064 305322
rect 261116 304020 261168 304026
rect 261116 303962 261168 303968
rect 261128 267170 261156 303962
rect 261220 267238 261248 305322
rect 261312 280906 261340 305510
rect 261496 304026 261524 310420
rect 261680 305250 261708 310420
rect 261772 310406 261970 310434
rect 261668 305244 261720 305250
rect 261668 305186 261720 305192
rect 261484 304020 261536 304026
rect 261484 303962 261536 303968
rect 261772 296714 261800 310406
rect 262140 305386 262168 310420
rect 262324 310406 262430 310434
rect 262128 305380 262180 305386
rect 262128 305322 262180 305328
rect 261404 296686 261800 296714
rect 261404 280974 261432 296686
rect 261392 280968 261444 280974
rect 261392 280910 261444 280916
rect 261300 280900 261352 280906
rect 261300 280842 261352 280848
rect 262324 272678 262352 310406
rect 262404 306400 262456 306406
rect 262404 306342 262456 306348
rect 262416 274106 262444 306342
rect 262496 306332 262548 306338
rect 262496 306274 262548 306280
rect 262508 282470 262536 306274
rect 262496 282464 262548 282470
rect 262496 282406 262548 282412
rect 262600 282402 262628 310420
rect 262692 310406 262890 310434
rect 262588 282396 262640 282402
rect 262588 282338 262640 282344
rect 262404 274100 262456 274106
rect 262404 274042 262456 274048
rect 262312 272672 262364 272678
rect 262312 272614 262364 272620
rect 262692 268530 262720 310406
rect 263060 306406 263088 310420
rect 263152 310406 263350 310434
rect 263048 306400 263100 306406
rect 263048 306342 263100 306348
rect 263152 306338 263180 310406
rect 263520 307834 263548 310420
rect 263692 308576 263744 308582
rect 263692 308518 263744 308524
rect 263600 308508 263652 308514
rect 263600 308450 263652 308456
rect 263508 307828 263560 307834
rect 263508 307770 263560 307776
rect 263140 306332 263192 306338
rect 263140 306274 263192 306280
rect 262680 268524 262732 268530
rect 262680 268466 262732 268472
rect 261208 267232 261260 267238
rect 261208 267174 261260 267180
rect 261116 267164 261168 267170
rect 261116 267106 261168 267112
rect 261024 265804 261076 265810
rect 261024 265746 261076 265752
rect 263612 261730 263640 308450
rect 263704 261798 263732 308518
rect 263796 268598 263824 310420
rect 263876 308440 263928 308446
rect 263876 308382 263928 308388
rect 263888 268666 263916 308382
rect 263980 275398 264008 310420
rect 264072 310406 264270 310434
rect 264072 308514 264100 310406
rect 264060 308508 264112 308514
rect 264060 308450 264112 308456
rect 264440 308446 264468 310420
rect 264532 310406 264730 310434
rect 264428 308440 264480 308446
rect 264428 308382 264480 308388
rect 264532 296714 264560 310406
rect 264900 308582 264928 310420
rect 264888 308576 264940 308582
rect 264888 308518 264940 308524
rect 265072 308576 265124 308582
rect 265072 308518 265124 308524
rect 264980 308236 265032 308242
rect 264980 308178 265032 308184
rect 264072 296686 264560 296714
rect 264072 275466 264100 296686
rect 264060 275460 264112 275466
rect 264060 275402 264112 275408
rect 263968 275392 264020 275398
rect 263968 275334 264020 275340
rect 263876 268660 263928 268666
rect 263876 268602 263928 268608
rect 263784 268592 263836 268598
rect 263784 268534 263836 268540
rect 264992 263090 265020 308178
rect 264980 263084 265032 263090
rect 264980 263026 265032 263032
rect 265084 263022 265112 308518
rect 265176 270026 265204 310420
rect 265374 310406 265480 310434
rect 265348 308508 265400 308514
rect 265348 308450 265400 308456
rect 265256 308440 265308 308446
rect 265256 308382 265308 308388
rect 265268 270094 265296 308382
rect 265360 276962 265388 308450
rect 265348 276956 265400 276962
rect 265348 276898 265400 276904
rect 265452 276894 265480 310406
rect 265544 310406 265650 310434
rect 265544 308582 265572 310406
rect 265532 308576 265584 308582
rect 265532 308518 265584 308524
rect 265820 308446 265848 310420
rect 265912 310406 266110 310434
rect 265912 308514 265940 310406
rect 265900 308508 265952 308514
rect 265900 308450 265952 308456
rect 265808 308440 265860 308446
rect 265808 308382 265860 308388
rect 266280 308242 266308 310420
rect 266464 310406 266570 310434
rect 266268 308236 266320 308242
rect 266268 308178 266320 308184
rect 265440 276888 265492 276894
rect 265440 276830 265492 276836
rect 266464 270162 266492 310406
rect 266544 308440 266596 308446
rect 266740 308394 266768 310420
rect 266544 308382 266596 308388
rect 266556 271386 266584 308382
rect 266648 308366 266768 308394
rect 266648 278186 266676 308366
rect 267016 307154 267044 310420
rect 267200 308446 267228 310420
rect 267292 310406 267490 310434
rect 267188 308440 267240 308446
rect 267188 308382 267240 308388
rect 267004 307148 267056 307154
rect 267004 307090 267056 307096
rect 267292 307034 267320 310406
rect 266740 307006 267320 307034
rect 266740 278254 266768 307006
rect 267660 296714 267688 310420
rect 267832 308576 267884 308582
rect 267832 308518 267884 308524
rect 267740 308508 267792 308514
rect 267740 308450 267792 308456
rect 266832 296686 267688 296714
rect 266728 278248 266780 278254
rect 266728 278190 266780 278196
rect 266636 278180 266688 278186
rect 266636 278122 266688 278128
rect 266544 271380 266596 271386
rect 266544 271322 266596 271328
rect 266452 270156 266504 270162
rect 266452 270098 266504 270104
rect 265256 270088 265308 270094
rect 265256 270030 265308 270036
rect 265164 270020 265216 270026
rect 265164 269962 265216 269968
rect 265072 263016 265124 263022
rect 265072 262958 265124 262964
rect 263692 261792 263744 261798
rect 263692 261734 263744 261740
rect 263600 261724 263652 261730
rect 263600 261666 263652 261672
rect 266832 260370 266860 296686
rect 267752 263158 267780 308450
rect 267844 264450 267872 308518
rect 267936 271454 267964 310420
rect 268016 308440 268068 308446
rect 268016 308382 268068 308388
rect 268028 271522 268056 308382
rect 268120 278322 268148 310420
rect 268212 310406 268410 310434
rect 268212 308514 268240 310406
rect 268200 308508 268252 308514
rect 268200 308450 268252 308456
rect 268580 308446 268608 310420
rect 268568 308440 268620 308446
rect 268568 308382 268620 308388
rect 268764 296714 268792 310420
rect 268856 310406 269054 310434
rect 269238 310406 269436 310434
rect 268856 308582 268884 310406
rect 268844 308576 268896 308582
rect 268844 308518 268896 308524
rect 269120 308576 269172 308582
rect 269120 308518 269172 308524
rect 268212 296686 268792 296714
rect 268212 279614 268240 296686
rect 268200 279608 268252 279614
rect 268200 279550 268252 279556
rect 268108 278316 268160 278322
rect 268108 278258 268160 278264
rect 268016 271516 268068 271522
rect 268016 271458 268068 271464
rect 267924 271448 267976 271454
rect 267924 271390 267976 271396
rect 269132 264586 269160 308518
rect 269212 308508 269264 308514
rect 269212 308450 269264 308456
rect 269120 264580 269172 264586
rect 269120 264522 269172 264528
rect 269224 264518 269252 308450
rect 269304 308440 269356 308446
rect 269304 308382 269356 308388
rect 269316 272814 269344 308382
rect 269304 272808 269356 272814
rect 269304 272750 269356 272756
rect 269408 272746 269436 310406
rect 269500 308394 269528 310420
rect 269684 308514 269712 310420
rect 269776 310406 269974 310434
rect 269672 308508 269724 308514
rect 269672 308450 269724 308456
rect 269776 308446 269804 310406
rect 269764 308440 269816 308446
rect 269500 308366 269620 308394
rect 269764 308382 269816 308388
rect 269488 308236 269540 308242
rect 269488 308178 269540 308184
rect 269500 279750 269528 308178
rect 269488 279744 269540 279750
rect 269488 279686 269540 279692
rect 269592 279682 269620 308366
rect 270144 308242 270172 310420
rect 270236 310406 270434 310434
rect 270618 310406 270816 310434
rect 270236 308582 270264 310406
rect 270224 308576 270276 308582
rect 270224 308518 270276 308524
rect 270500 308576 270552 308582
rect 270500 308518 270552 308524
rect 270132 308236 270184 308242
rect 270132 308178 270184 308184
rect 269580 279676 269632 279682
rect 269580 279618 269632 279624
rect 269396 272740 269448 272746
rect 269396 272682 269448 272688
rect 269212 264512 269264 264518
rect 269212 264454 269264 264460
rect 267832 264444 267884 264450
rect 267832 264386 267884 264392
rect 267740 263152 267792 263158
rect 267740 263094 267792 263100
rect 266820 260364 266872 260370
rect 266820 260306 266872 260312
rect 270512 249218 270540 308518
rect 270684 308508 270736 308514
rect 270684 308450 270736 308456
rect 270592 308440 270644 308446
rect 270592 308382 270644 308388
rect 270604 265878 270632 308382
rect 270696 265946 270724 308450
rect 270788 272882 270816 310406
rect 270880 308394 270908 310420
rect 271064 308446 271092 310420
rect 271156 310406 271354 310434
rect 271052 308440 271104 308446
rect 270880 308366 271000 308394
rect 271052 308382 271104 308388
rect 270868 308236 270920 308242
rect 270868 308178 270920 308184
rect 270880 274174 270908 308178
rect 270972 281042 271000 308366
rect 271156 308242 271184 310406
rect 271524 308582 271552 310420
rect 271616 310406 271814 310434
rect 271998 310406 272104 310434
rect 271512 308576 271564 308582
rect 271512 308518 271564 308524
rect 271616 308514 271644 310406
rect 271604 308508 271656 308514
rect 271604 308450 271656 308456
rect 271972 308508 272024 308514
rect 271972 308450 272024 308456
rect 271144 308236 271196 308242
rect 271144 308178 271196 308184
rect 271696 306400 271748 306406
rect 271696 306342 271748 306348
rect 271708 306202 271736 306342
rect 271696 306196 271748 306202
rect 271696 306138 271748 306144
rect 270960 281036 271012 281042
rect 270960 280978 271012 280984
rect 270868 274168 270920 274174
rect 270868 274110 270920 274116
rect 270776 272876 270828 272882
rect 270776 272818 270828 272824
rect 271984 266014 272012 308450
rect 272076 274242 272104 310406
rect 272156 308440 272208 308446
rect 272156 308382 272208 308388
rect 272064 274236 272116 274242
rect 272064 274178 272116 274184
rect 272168 273873 272196 308382
rect 272260 281110 272288 310420
rect 272444 307222 272472 310420
rect 272536 310406 272734 310434
rect 272536 308446 272564 310406
rect 272524 308440 272576 308446
rect 272524 308382 272576 308388
rect 272432 307216 272484 307222
rect 272432 307158 272484 307164
rect 272904 296714 272932 310420
rect 272996 310406 273194 310434
rect 272996 308514 273024 310406
rect 272984 308508 273036 308514
rect 272984 308450 273036 308456
rect 273364 306354 273392 310420
rect 272352 296686 272932 296714
rect 273272 306326 273392 306354
rect 273456 310406 273654 310434
rect 272248 281104 272300 281110
rect 272248 281046 272300 281052
rect 272154 273864 272210 273873
rect 272154 273799 272210 273808
rect 271972 266008 272024 266014
rect 271972 265950 272024 265956
rect 270684 265940 270736 265946
rect 270684 265882 270736 265888
rect 270592 265872 270644 265878
rect 270592 265814 270644 265820
rect 272352 249286 272380 296686
rect 272340 249280 272392 249286
rect 272340 249222 272392 249228
rect 270500 249212 270552 249218
rect 270500 249154 270552 249160
rect 260932 247920 260984 247926
rect 260932 247862 260984 247868
rect 259552 247852 259604 247858
rect 259552 247794 259604 247800
rect 273272 246634 273300 306326
rect 273456 306218 273484 310406
rect 273824 306354 273852 310420
rect 273364 306190 273484 306218
rect 273548 306326 273852 306354
rect 273916 310406 274114 310434
rect 273364 249121 273392 306190
rect 273444 303748 273496 303754
rect 273444 303690 273496 303696
rect 273456 262857 273484 303690
rect 273548 267073 273576 306326
rect 273916 302234 273944 310406
rect 273640 302206 273944 302234
rect 273640 275233 273668 302206
rect 274284 296714 274312 310420
rect 274376 310406 274574 310434
rect 274376 303754 274404 310406
rect 274364 303748 274416 303754
rect 274364 303690 274416 303696
rect 274744 303385 274772 310420
rect 275020 306105 275048 310420
rect 275204 308961 275232 310420
rect 275190 308952 275246 308961
rect 275190 308887 275246 308896
rect 275006 306096 275062 306105
rect 275006 306031 275062 306040
rect 275480 305454 275508 310420
rect 275664 306241 275692 310420
rect 275940 308689 275968 310420
rect 275926 308680 275982 308689
rect 275926 308615 275982 308624
rect 275650 306232 275706 306241
rect 275650 306167 275706 306176
rect 276124 305590 276152 310420
rect 276112 305584 276164 305590
rect 276112 305526 276164 305532
rect 276308 305522 276336 310420
rect 276584 308825 276612 310420
rect 276570 308816 276626 308825
rect 276570 308751 276626 308760
rect 276768 306406 276796 310420
rect 276756 306400 276808 306406
rect 276756 306342 276808 306348
rect 276296 305516 276348 305522
rect 276296 305458 276348 305464
rect 275468 305448 275520 305454
rect 275468 305390 275520 305396
rect 274730 303376 274786 303385
rect 274730 303311 274786 303320
rect 277044 303249 277072 310420
rect 277228 308553 277256 310420
rect 277214 308544 277270 308553
rect 277214 308479 277270 308488
rect 277504 305969 277532 310420
rect 277490 305960 277546 305969
rect 277490 305895 277546 305904
rect 277030 303240 277086 303249
rect 277030 303175 277086 303184
rect 277688 302977 277716 310420
rect 277964 308174 277992 310420
rect 277952 308168 278004 308174
rect 277952 308110 278004 308116
rect 278148 306066 278176 310420
rect 278136 306060 278188 306066
rect 278136 306002 278188 306008
rect 278424 303113 278452 310420
rect 278608 308310 278636 310420
rect 278596 308304 278648 308310
rect 278596 308246 278648 308252
rect 278884 306134 278912 310420
rect 278872 306128 278924 306134
rect 278872 306070 278924 306076
rect 278410 303104 278466 303113
rect 278410 303039 278466 303048
rect 277674 302968 277730 302977
rect 277674 302903 277730 302912
rect 279068 302841 279096 310420
rect 279344 308378 279372 310420
rect 279332 308372 279384 308378
rect 279332 308314 279384 308320
rect 279528 305998 279556 310420
rect 279516 305992 279568 305998
rect 279516 305934 279568 305940
rect 279804 303618 279832 310420
rect 279988 309126 280016 310420
rect 279976 309120 280028 309126
rect 279976 309062 280028 309068
rect 280264 305930 280292 310420
rect 280252 305924 280304 305930
rect 280252 305866 280304 305872
rect 279792 303612 279844 303618
rect 279792 303554 279844 303560
rect 279054 302832 279110 302841
rect 280448 302802 280476 310420
rect 280724 305697 280752 310420
rect 280908 305833 280936 310420
rect 280894 305824 280950 305833
rect 280894 305759 280950 305768
rect 280710 305688 280766 305697
rect 280710 305623 280766 305632
rect 279054 302767 279110 302776
rect 280436 302796 280488 302802
rect 280436 302738 280488 302744
rect 281184 302734 281212 310420
rect 281368 306338 281396 310420
rect 281356 306332 281408 306338
rect 281356 306274 281408 306280
rect 281644 305726 281672 310420
rect 281632 305720 281684 305726
rect 281632 305662 281684 305668
rect 281828 303210 281856 310420
rect 282104 303550 282132 310420
rect 282288 305862 282316 310420
rect 282276 305856 282328 305862
rect 282276 305798 282328 305804
rect 282092 303544 282144 303550
rect 282092 303486 282144 303492
rect 282564 303346 282592 310420
rect 282748 303414 282776 310420
rect 282736 303408 282788 303414
rect 282736 303350 282788 303356
rect 282552 303340 282604 303346
rect 282552 303282 282604 303288
rect 283024 303278 283052 310420
rect 283012 303272 283064 303278
rect 283012 303214 283064 303220
rect 281816 303204 281868 303210
rect 281816 303146 281868 303152
rect 281172 302728 281224 302734
rect 281172 302670 281224 302676
rect 283208 302234 283236 310420
rect 283392 303482 283420 310420
rect 283380 303476 283432 303482
rect 283380 303418 283432 303424
rect 283668 302870 283696 310420
rect 283656 302864 283708 302870
rect 283656 302806 283708 302812
rect 283852 302234 283880 310420
rect 283116 302206 283236 302234
rect 283300 302206 283880 302234
rect 283944 310406 284142 310434
rect 284326 310406 284524 310434
rect 283116 300257 283144 302206
rect 283300 300393 283328 302206
rect 283944 300830 283972 310406
rect 284300 306400 284352 306406
rect 284300 306342 284352 306348
rect 283932 300824 283984 300830
rect 283932 300766 283984 300772
rect 284312 300626 284340 306342
rect 284392 306332 284444 306338
rect 284392 306274 284444 306280
rect 284300 300620 284352 300626
rect 284300 300562 284352 300568
rect 283286 300384 283342 300393
rect 283286 300319 283342 300328
rect 284404 300286 284432 306274
rect 284496 306218 284524 310406
rect 284588 306354 284616 310420
rect 284588 306326 284708 306354
rect 284772 306338 284800 310420
rect 284864 310406 285062 310434
rect 284496 306190 284616 306218
rect 284484 306128 284536 306134
rect 284484 306070 284536 306076
rect 284392 300280 284444 300286
rect 283102 300248 283158 300257
rect 284392 300222 284444 300228
rect 284496 300218 284524 306070
rect 283102 300183 283158 300192
rect 284484 300212 284536 300218
rect 284484 300154 284536 300160
rect 284588 300121 284616 306190
rect 284680 300150 284708 306326
rect 284760 306332 284812 306338
rect 284760 306274 284812 306280
rect 284864 306134 284892 310406
rect 285232 306406 285260 310420
rect 285324 310406 285522 310434
rect 285706 310406 285812 310434
rect 285220 306400 285272 306406
rect 285220 306342 285272 306348
rect 284852 306128 284904 306134
rect 284852 306070 284904 306076
rect 284668 300144 284720 300150
rect 284574 300112 284630 300121
rect 284668 300086 284720 300092
rect 284574 300047 284630 300056
rect 285324 299946 285352 310406
rect 285680 306468 285732 306474
rect 285680 306410 285732 306416
rect 285692 302234 285720 306410
rect 285784 306270 285812 310406
rect 285968 306746 285996 310420
rect 285956 306740 286008 306746
rect 285956 306682 286008 306688
rect 286152 306626 286180 310420
rect 285876 306598 286180 306626
rect 286244 310406 286442 310434
rect 285772 306264 285824 306270
rect 285772 306206 285824 306212
rect 285692 302206 285812 302234
rect 285312 299940 285364 299946
rect 285312 299882 285364 299888
rect 273732 296686 274312 296714
rect 273732 281178 273760 296686
rect 273720 281172 273772 281178
rect 273720 281114 273772 281120
rect 273626 275224 273682 275233
rect 273626 275159 273682 275168
rect 273534 267064 273590 267073
rect 273534 266999 273590 267008
rect 273442 262848 273498 262857
rect 273442 262783 273498 262792
rect 273350 249112 273406 249121
rect 273350 249047 273406 249056
rect 273260 246628 273312 246634
rect 273260 246570 273312 246576
rect 259460 245200 259512 245206
rect 259460 245142 259512 245148
rect 256700 245064 256752 245070
rect 256700 245006 256752 245012
rect 232044 244928 232096 244934
rect 232044 244870 232096 244876
rect 285784 243642 285812 302206
rect 285876 300762 285904 306598
rect 285956 306536 286008 306542
rect 285956 306478 286008 306484
rect 285864 300756 285916 300762
rect 285864 300698 285916 300704
rect 285968 300082 285996 306478
rect 286244 306474 286272 310406
rect 286232 306468 286284 306474
rect 286232 306410 286284 306416
rect 286612 306354 286640 310420
rect 286888 308922 286916 310420
rect 286876 308916 286928 308922
rect 286876 308858 286928 308864
rect 286060 306326 286640 306354
rect 285956 300076 286008 300082
rect 285956 300018 286008 300024
rect 286060 243710 286088 306326
rect 286140 306264 286192 306270
rect 286140 306206 286192 306212
rect 286152 300558 286180 306206
rect 287072 303142 287100 310420
rect 287152 306536 287204 306542
rect 287152 306478 287204 306484
rect 287164 305794 287192 306478
rect 287348 306354 287376 310420
rect 287532 306542 287560 310420
rect 287624 310406 287822 310434
rect 287520 306536 287572 306542
rect 287520 306478 287572 306484
rect 287244 306332 287296 306338
rect 287348 306326 287560 306354
rect 287244 306274 287296 306280
rect 287152 305788 287204 305794
rect 287152 305730 287204 305736
rect 287060 303136 287112 303142
rect 287060 303078 287112 303084
rect 286140 300552 286192 300558
rect 286140 300494 286192 300500
rect 287256 300014 287284 306274
rect 287336 306264 287388 306270
rect 287336 306206 287388 306212
rect 287244 300008 287296 300014
rect 287244 299950 287296 299956
rect 286048 243704 286100 243710
rect 286048 243646 286100 243652
rect 285772 243636 285824 243642
rect 285772 243578 285824 243584
rect 287348 243574 287376 306206
rect 287428 306196 287480 306202
rect 287428 306138 287480 306144
rect 287440 245410 287468 306138
rect 287532 300694 287560 306326
rect 287624 306270 287652 310406
rect 287992 306338 288020 310420
rect 288084 310406 288282 310434
rect 288466 310406 288572 310434
rect 287980 306332 288032 306338
rect 287980 306274 288032 306280
rect 287612 306264 287664 306270
rect 287612 306206 287664 306212
rect 288084 306202 288112 310406
rect 288440 306332 288492 306338
rect 288440 306274 288492 306280
rect 288072 306196 288124 306202
rect 288072 306138 288124 306144
rect 287520 300688 287572 300694
rect 287520 300630 287572 300636
rect 287428 245404 287480 245410
rect 287428 245346 287480 245352
rect 288452 243574 288480 306274
rect 288544 245342 288572 310406
rect 288636 310406 288742 310434
rect 288532 245336 288584 245342
rect 288532 245278 288584 245284
rect 288636 245274 288664 310406
rect 288912 308922 288940 310420
rect 288900 308916 288952 308922
rect 288900 308858 288952 308864
rect 289188 308378 289216 310420
rect 289176 308372 289228 308378
rect 289176 308314 289228 308320
rect 289372 306338 289400 310420
rect 289464 310406 289662 310434
rect 289846 310406 289952 310434
rect 289360 306332 289412 306338
rect 289360 306274 289412 306280
rect 289464 296714 289492 310406
rect 289820 306332 289872 306338
rect 289820 306274 289872 306280
rect 288728 296686 289492 296714
rect 288728 247722 288756 296686
rect 288716 247716 288768 247722
rect 288716 247658 288768 247664
rect 288624 245268 288676 245274
rect 288624 245210 288676 245216
rect 289832 243642 289860 306274
rect 289924 243710 289952 310406
rect 290016 310406 290122 310434
rect 290016 246566 290044 310406
rect 290292 308650 290320 310420
rect 290280 308644 290332 308650
rect 290280 308586 290332 308592
rect 290476 306338 290504 310420
rect 290752 308786 290780 310420
rect 290740 308780 290792 308786
rect 290740 308722 290792 308728
rect 290936 308718 290964 310420
rect 290924 308712 290976 308718
rect 290924 308654 290976 308660
rect 291212 306354 291240 310420
rect 291396 308582 291424 310420
rect 291488 310406 291686 310434
rect 291384 308576 291436 308582
rect 291384 308518 291436 308524
rect 290464 306332 290516 306338
rect 291212 306326 291424 306354
rect 290464 306274 290516 306280
rect 291200 306264 291252 306270
rect 291200 306206 291252 306212
rect 290004 246560 290056 246566
rect 290004 246502 290056 246508
rect 291212 243778 291240 306206
rect 291292 303612 291344 303618
rect 291292 303554 291344 303560
rect 291304 245206 291332 303554
rect 291396 247790 291424 306326
rect 291488 303618 291516 310406
rect 291476 303612 291528 303618
rect 291476 303554 291528 303560
rect 291476 303476 291528 303482
rect 291476 303418 291528 303424
rect 291488 250646 291516 303418
rect 291856 296714 291884 310420
rect 291948 310406 292146 310434
rect 291948 303482 291976 310406
rect 292316 306270 292344 310420
rect 292592 306354 292620 310420
rect 292790 310406 292988 310434
rect 292592 306326 292896 306354
rect 292304 306264 292356 306270
rect 292304 306206 292356 306212
rect 292764 306264 292816 306270
rect 292764 306206 292816 306212
rect 292580 306196 292632 306202
rect 292580 306138 292632 306144
rect 291936 303476 291988 303482
rect 291936 303418 291988 303424
rect 291580 296686 291884 296714
rect 291476 250640 291528 250646
rect 291476 250582 291528 250588
rect 291580 250510 291608 296686
rect 291568 250504 291620 250510
rect 291568 250446 291620 250452
rect 291384 247784 291436 247790
rect 291384 247726 291436 247732
rect 292592 245274 292620 306138
rect 292672 306128 292724 306134
rect 292672 306070 292724 306076
rect 292684 247926 292712 306070
rect 292672 247920 292724 247926
rect 292672 247862 292724 247868
rect 292776 247858 292804 306206
rect 292868 251190 292896 306326
rect 292856 251184 292908 251190
rect 292856 251126 292908 251132
rect 292960 250986 292988 310406
rect 293052 306202 293080 310420
rect 293236 306270 293264 310420
rect 293328 310406 293526 310434
rect 293224 306264 293276 306270
rect 293224 306206 293276 306212
rect 293040 306196 293092 306202
rect 293040 306138 293092 306144
rect 293328 296714 293356 310406
rect 293696 306134 293724 310420
rect 293972 308854 294000 310420
rect 294170 310406 294276 310434
rect 293960 308848 294012 308854
rect 293960 308790 294012 308796
rect 293960 306400 294012 306406
rect 293960 306342 294012 306348
rect 293684 306128 293736 306134
rect 293684 306070 293736 306076
rect 293052 296686 293356 296714
rect 292948 250980 293000 250986
rect 292948 250922 293000 250928
rect 293052 250714 293080 296686
rect 293040 250708 293092 250714
rect 293040 250650 293092 250656
rect 292764 247852 292816 247858
rect 292764 247794 292816 247800
rect 293972 245342 294000 306342
rect 294144 306332 294196 306338
rect 294144 306274 294196 306280
rect 294052 305788 294104 305794
rect 294052 305730 294104 305736
rect 294064 245410 294092 305730
rect 294156 247654 294184 306274
rect 294248 253502 294276 310406
rect 294432 308689 294460 310420
rect 294418 308680 294474 308689
rect 294418 308615 294474 308624
rect 294616 306338 294644 310420
rect 294708 310406 294906 310434
rect 294708 306406 294736 310406
rect 294696 306400 294748 306406
rect 294696 306342 294748 306348
rect 294604 306332 294656 306338
rect 294604 306274 294656 306280
rect 295076 305794 295104 310420
rect 295352 306354 295380 310420
rect 295352 306326 295472 306354
rect 295340 306264 295392 306270
rect 295340 306206 295392 306212
rect 295064 305788 295116 305794
rect 295064 305730 295116 305736
rect 294236 253496 294288 253502
rect 294236 253438 294288 253444
rect 294144 247648 294196 247654
rect 294144 247590 294196 247596
rect 294052 245404 294104 245410
rect 294052 245346 294104 245352
rect 293960 245336 294012 245342
rect 293960 245278 294012 245284
rect 292580 245268 292632 245274
rect 292580 245210 292632 245216
rect 291292 245200 291344 245206
rect 291292 245142 291344 245148
rect 295352 245041 295380 306206
rect 295444 247586 295472 306326
rect 295536 305130 295564 310420
rect 295812 306270 295840 310420
rect 295800 306264 295852 306270
rect 295800 306206 295852 306212
rect 295536 305102 295748 305130
rect 295524 304972 295576 304978
rect 295524 304914 295576 304920
rect 295432 247580 295484 247586
rect 295432 247522 295484 247528
rect 295338 245032 295394 245041
rect 295338 244967 295394 244976
rect 295536 244905 295564 304914
rect 295616 303204 295668 303210
rect 295616 303146 295668 303152
rect 295628 248266 295656 303146
rect 295720 250306 295748 305102
rect 295996 303210 296024 310420
rect 296088 310406 296286 310434
rect 295984 303204 296036 303210
rect 295984 303146 296036 303152
rect 296088 296714 296116 310406
rect 296456 304978 296484 310420
rect 296732 306354 296760 310420
rect 296930 310406 297128 310434
rect 296732 306326 297036 306354
rect 296720 306264 296772 306270
rect 296720 306206 296772 306212
rect 296444 304972 296496 304978
rect 296444 304914 296496 304920
rect 295812 296686 296116 296714
rect 295812 250918 295840 296686
rect 295800 250912 295852 250918
rect 295800 250854 295852 250860
rect 295708 250300 295760 250306
rect 295708 250242 295760 250248
rect 295616 248260 295668 248266
rect 295616 248202 295668 248208
rect 296732 245449 296760 306206
rect 296904 306196 296956 306202
rect 296904 306138 296956 306144
rect 296812 306128 296864 306134
rect 296812 306070 296864 306076
rect 296824 247994 296852 306070
rect 296812 247988 296864 247994
rect 296812 247930 296864 247936
rect 296718 245440 296774 245449
rect 296718 245375 296774 245384
rect 296916 245177 296944 306138
rect 297008 248130 297036 306326
rect 297100 306320 297128 310406
rect 297192 306610 297220 310420
rect 297272 308916 297324 308922
rect 297272 308858 297324 308864
rect 297284 308582 297312 308858
rect 297272 308576 297324 308582
rect 297272 308518 297324 308524
rect 297180 306604 297232 306610
rect 297180 306546 297232 306552
rect 297100 306292 297312 306320
rect 297088 304360 297140 304366
rect 297088 304302 297140 304308
rect 296996 248124 297048 248130
rect 296996 248066 297048 248072
rect 297100 248062 297128 304302
rect 297284 299474 297312 306292
rect 297376 304366 297404 310420
rect 297468 310406 297666 310434
rect 297364 304360 297416 304366
rect 297364 304302 297416 304308
rect 297192 299446 297312 299474
rect 297192 250850 297220 299446
rect 297468 296714 297496 310406
rect 297836 306202 297864 310420
rect 297824 306196 297876 306202
rect 297824 306138 297876 306144
rect 298020 306134 298048 310420
rect 298192 306400 298244 306406
rect 298192 306342 298244 306348
rect 298296 306354 298324 310420
rect 298480 308825 298508 310420
rect 298572 310406 298770 310434
rect 298466 308816 298522 308825
rect 298466 308751 298522 308760
rect 298100 306332 298152 306338
rect 298100 306274 298152 306280
rect 298008 306128 298060 306134
rect 298008 306070 298060 306076
rect 297284 296686 297496 296714
rect 297180 250844 297232 250850
rect 297180 250786 297232 250792
rect 297284 250442 297312 296686
rect 297272 250436 297324 250442
rect 297272 250378 297324 250384
rect 297088 248056 297140 248062
rect 297088 247998 297140 248004
rect 298112 245313 298140 306274
rect 298204 248198 298232 306342
rect 298296 306326 298416 306354
rect 298284 306264 298336 306270
rect 298284 306206 298336 306212
rect 298296 248334 298324 306206
rect 298388 251122 298416 306326
rect 298572 306270 298600 310406
rect 298560 306264 298612 306270
rect 298560 306206 298612 306212
rect 298940 296714 298968 310420
rect 299032 310406 299230 310434
rect 299032 306338 299060 310406
rect 299400 306406 299428 310420
rect 299480 306468 299532 306474
rect 299480 306410 299532 306416
rect 299388 306400 299440 306406
rect 299388 306342 299440 306348
rect 299020 306332 299072 306338
rect 299020 306274 299072 306280
rect 298480 296686 298968 296714
rect 298376 251116 298428 251122
rect 298376 251058 298428 251064
rect 298480 250782 298508 296686
rect 298468 250776 298520 250782
rect 298468 250718 298520 250724
rect 298284 248328 298336 248334
rect 298284 248270 298336 248276
rect 298192 248192 298244 248198
rect 298192 248134 298244 248140
rect 299492 245585 299520 306410
rect 299572 306332 299624 306338
rect 299572 306274 299624 306280
rect 299584 248169 299612 306274
rect 299676 306134 299704 310420
rect 299860 306474 299888 310420
rect 299952 310406 300150 310434
rect 299848 306468 299900 306474
rect 299848 306410 299900 306416
rect 299952 306354 299980 310406
rect 299768 306326 299980 306354
rect 299664 306128 299716 306134
rect 299664 306070 299716 306076
rect 299664 305992 299716 305998
rect 299664 305934 299716 305940
rect 299570 248160 299626 248169
rect 299570 248095 299626 248104
rect 299478 245576 299534 245585
rect 299478 245511 299534 245520
rect 298098 245304 298154 245313
rect 298098 245239 298154 245248
rect 296902 245168 296958 245177
rect 296902 245103 296958 245112
rect 295522 244896 295578 244905
rect 295522 244831 295578 244840
rect 299676 244769 299704 305934
rect 299768 248402 299796 306326
rect 300320 306252 300348 310420
rect 299860 306224 300348 306252
rect 300412 310406 300610 310434
rect 299860 250889 299888 306224
rect 299940 306128 299992 306134
rect 299940 306070 299992 306076
rect 299952 251054 299980 306070
rect 300412 305998 300440 310406
rect 300780 306338 300808 310420
rect 300768 306332 300820 306338
rect 300768 306274 300820 306280
rect 300952 306332 301004 306338
rect 300952 306274 301004 306280
rect 300400 305992 300452 305998
rect 300400 305934 300452 305940
rect 300860 304972 300912 304978
rect 300860 304914 300912 304920
rect 299940 251048 299992 251054
rect 299940 250990 299992 250996
rect 299846 250880 299902 250889
rect 299846 250815 299902 250824
rect 299756 248396 299808 248402
rect 299756 248338 299808 248344
rect 300872 245614 300900 304914
rect 300860 245608 300912 245614
rect 300860 245550 300912 245556
rect 300964 245546 300992 306274
rect 301056 306270 301084 310420
rect 301240 306354 301268 310420
rect 301148 306326 301268 306354
rect 301332 310406 301530 310434
rect 301332 306338 301360 310406
rect 301320 306332 301372 306338
rect 301044 306264 301096 306270
rect 301044 306206 301096 306212
rect 301044 306128 301096 306134
rect 301044 306070 301096 306076
rect 301056 246265 301084 306070
rect 301148 247518 301176 306326
rect 301320 306274 301372 306280
rect 301228 306264 301280 306270
rect 301228 306206 301280 306212
rect 301240 250374 301268 306206
rect 301700 304978 301728 310420
rect 301792 310406 301990 310434
rect 301688 304972 301740 304978
rect 301688 304914 301740 304920
rect 301792 296714 301820 310406
rect 302160 306134 302188 310420
rect 302252 310406 302450 310434
rect 302148 306128 302200 306134
rect 302148 306070 302200 306076
rect 301332 296686 301820 296714
rect 301332 264217 301360 296686
rect 301318 264208 301374 264217
rect 301318 264143 301374 264152
rect 302252 254697 302280 310406
rect 302620 306354 302648 310420
rect 302344 306326 302648 306354
rect 302712 310406 302910 310434
rect 302344 265577 302372 306326
rect 302516 306264 302568 306270
rect 302516 306206 302568 306212
rect 302424 306196 302476 306202
rect 302424 306138 302476 306144
rect 302330 265568 302386 265577
rect 302330 265503 302386 265512
rect 302238 254688 302294 254697
rect 302238 254623 302294 254632
rect 302436 254561 302464 306138
rect 302528 268666 302556 306206
rect 302712 302234 302740 310406
rect 303080 306202 303108 310420
rect 303172 310406 303370 310434
rect 303172 306270 303200 310406
rect 303160 306264 303212 306270
rect 303160 306206 303212 306212
rect 303068 306196 303120 306202
rect 303068 306138 303120 306144
rect 302620 302206 302740 302234
rect 302620 282169 302648 302206
rect 303540 296714 303568 310420
rect 303816 306610 303844 310420
rect 303804 306604 303856 306610
rect 303804 306546 303856 306552
rect 304000 306490 304028 310420
rect 303724 306462 304028 306490
rect 304092 310406 304290 310434
rect 303620 306332 303672 306338
rect 303620 306274 303672 306280
rect 302712 296686 303568 296714
rect 302712 283529 302740 296686
rect 302698 283520 302754 283529
rect 302698 283455 302754 283464
rect 302606 282160 302662 282169
rect 302606 282095 302662 282104
rect 303632 269958 303660 306274
rect 303620 269952 303672 269958
rect 303620 269894 303672 269900
rect 303724 269793 303752 306462
rect 304092 306218 304120 310406
rect 304172 306604 304224 306610
rect 304172 306546 304224 306552
rect 303816 306190 304120 306218
rect 303816 285258 303844 306190
rect 303896 306128 303948 306134
rect 303896 306070 303948 306076
rect 303908 286550 303936 306070
rect 304184 302234 304212 306546
rect 304000 302206 304212 302234
rect 304000 297401 304028 302206
rect 304460 298994 304488 310420
rect 304552 310406 304750 310434
rect 304552 306338 304580 310406
rect 304540 306332 304592 306338
rect 304540 306274 304592 306280
rect 304920 306134 304948 310420
rect 305104 306490 305132 310420
rect 305012 306462 305132 306490
rect 305196 310406 305394 310434
rect 305012 306270 305040 306462
rect 305196 306354 305224 310406
rect 305564 306354 305592 310420
rect 305104 306326 305224 306354
rect 305288 306326 305592 306354
rect 305656 310406 305854 310434
rect 305000 306264 305052 306270
rect 305000 306206 305052 306212
rect 304908 306128 304960 306134
rect 304908 306070 304960 306076
rect 305000 306128 305052 306134
rect 305000 306070 305052 306076
rect 304448 298988 304500 298994
rect 304448 298930 304500 298936
rect 303986 297392 304042 297401
rect 303986 297327 304042 297336
rect 303896 286544 303948 286550
rect 303896 286486 303948 286492
rect 303804 285252 303856 285258
rect 303804 285194 303856 285200
rect 303710 269784 303766 269793
rect 303710 269719 303766 269728
rect 302516 268660 302568 268666
rect 302516 268602 302568 268608
rect 302422 254552 302478 254561
rect 302422 254487 302478 254496
rect 305012 250578 305040 306070
rect 305104 269890 305132 306326
rect 305184 303204 305236 303210
rect 305184 303146 305236 303152
rect 305196 271386 305224 303146
rect 305288 286482 305316 306326
rect 305368 306264 305420 306270
rect 305368 306206 305420 306212
rect 305380 300558 305408 306206
rect 305656 301481 305684 310406
rect 306024 303210 306052 310420
rect 306116 310406 306314 310434
rect 306116 306134 306144 310406
rect 306380 306604 306432 306610
rect 306380 306546 306432 306552
rect 306104 306128 306156 306134
rect 306104 306070 306156 306076
rect 306012 303204 306064 303210
rect 306012 303146 306064 303152
rect 305642 301472 305698 301481
rect 305642 301407 305698 301416
rect 305368 300552 305420 300558
rect 305368 300494 305420 300500
rect 305276 286476 305328 286482
rect 305276 286418 305328 286424
rect 305184 271380 305236 271386
rect 305184 271322 305236 271328
rect 305092 269884 305144 269890
rect 305092 269826 305144 269832
rect 306392 250753 306420 306546
rect 306484 306338 306512 310420
rect 306576 310406 306774 310434
rect 306472 306332 306524 306338
rect 306472 306274 306524 306280
rect 306472 306196 306524 306202
rect 306472 306138 306524 306144
rect 306484 271250 306512 306138
rect 306576 271318 306604 310406
rect 306944 306610 306972 310420
rect 306932 306604 306984 306610
rect 306932 306546 306984 306552
rect 306656 306400 306708 306406
rect 306656 306342 306708 306348
rect 306668 286414 306696 306342
rect 306748 306332 306800 306338
rect 306748 306274 306800 306280
rect 306760 301714 306788 306274
rect 307220 302977 307248 310420
rect 307404 306202 307432 310420
rect 307496 310406 307694 310434
rect 307496 306406 307524 310406
rect 307760 306876 307812 306882
rect 307760 306818 307812 306824
rect 307484 306400 307536 306406
rect 307484 306342 307536 306348
rect 307392 306196 307444 306202
rect 307392 306138 307444 306144
rect 307206 302968 307262 302977
rect 307206 302903 307262 302912
rect 306748 301708 306800 301714
rect 306748 301650 306800 301656
rect 306656 286408 306708 286414
rect 306656 286350 306708 286356
rect 307772 272678 307800 306818
rect 307864 303249 307892 310420
rect 307956 310406 308154 310434
rect 307956 306882 307984 310406
rect 307944 306876 307996 306882
rect 307944 306818 307996 306824
rect 307944 305380 307996 305386
rect 307944 305322 307996 305328
rect 307850 303240 307906 303249
rect 307850 303175 307906 303184
rect 307852 302796 307904 302802
rect 307852 302738 307904 302744
rect 307760 272672 307812 272678
rect 307760 272614 307812 272620
rect 307864 272610 307892 302738
rect 307956 287842 307984 305322
rect 308324 302234 308352 310420
rect 308600 303113 308628 310420
rect 308586 303104 308642 303113
rect 308586 303039 308642 303048
rect 308784 302802 308812 310420
rect 308876 310406 309074 310434
rect 309336 310406 309534 310434
rect 308876 305386 308904 310406
rect 309336 306490 309364 310406
rect 309152 306462 309364 306490
rect 308864 305380 308916 305386
rect 308864 305322 308916 305328
rect 308772 302796 308824 302802
rect 308772 302738 308824 302744
rect 308048 302206 308352 302234
rect 308048 287910 308076 302206
rect 308036 287904 308088 287910
rect 308036 287846 308088 287852
rect 307944 287836 307996 287842
rect 307944 287778 307996 287784
rect 307852 272604 307904 272610
rect 307852 272546 307904 272552
rect 309152 272542 309180 306462
rect 309704 306354 309732 310420
rect 309232 306332 309284 306338
rect 309232 306274 309284 306280
rect 309336 306326 309732 306354
rect 309244 274174 309272 306274
rect 309336 287774 309364 306326
rect 309796 304201 309824 310490
rect 309980 304502 310008 310420
rect 310164 306338 310192 310420
rect 310256 310406 310454 310434
rect 310716 310406 310914 310434
rect 310152 306332 310204 306338
rect 310152 306274 310204 306280
rect 309968 304496 310020 304502
rect 309968 304438 310020 304444
rect 309782 304192 309838 304201
rect 309782 304127 309838 304136
rect 310256 302234 310284 310406
rect 310716 306490 310744 310406
rect 309428 302206 310284 302234
rect 310532 306462 310744 306490
rect 309428 289338 309456 302206
rect 309416 289332 309468 289338
rect 309416 289274 309468 289280
rect 309324 287768 309376 287774
rect 309324 287710 309376 287716
rect 309232 274168 309284 274174
rect 309232 274110 309284 274116
rect 309140 272536 309192 272542
rect 309140 272478 309192 272484
rect 306564 271312 306616 271318
rect 306564 271254 306616 271260
rect 306472 271244 306524 271250
rect 306472 271186 306524 271192
rect 306378 250744 306434 250753
rect 306378 250679 306434 250688
rect 305000 250572 305052 250578
rect 305000 250514 305052 250520
rect 301228 250368 301280 250374
rect 301228 250310 301280 250316
rect 301136 247512 301188 247518
rect 301136 247454 301188 247460
rect 310532 246498 310560 306462
rect 311084 306354 311112 310420
rect 310612 306332 310664 306338
rect 310612 306274 310664 306280
rect 310716 306326 311112 306354
rect 310624 274106 310652 306274
rect 310716 289270 310744 306326
rect 311176 304434 311204 310490
rect 311360 306105 311388 310420
rect 311544 306338 311572 310420
rect 311636 310406 311834 310434
rect 311532 306332 311584 306338
rect 311532 306274 311584 306280
rect 311346 306096 311402 306105
rect 311346 306031 311402 306040
rect 311164 304428 311216 304434
rect 311164 304370 311216 304376
rect 311636 302234 311664 310406
rect 312004 308922 312032 310420
rect 311992 308916 312044 308922
rect 311992 308858 312044 308864
rect 312188 308530 312216 310420
rect 310808 302206 311664 302234
rect 311912 308502 312216 308530
rect 312280 310406 312478 310434
rect 310704 289264 310756 289270
rect 310704 289206 310756 289212
rect 310808 289202 310836 302206
rect 310796 289196 310848 289202
rect 310796 289138 310848 289144
rect 310612 274100 310664 274106
rect 310612 274042 310664 274048
rect 311912 263090 311940 308502
rect 312280 308394 312308 310406
rect 312360 308916 312412 308922
rect 312360 308858 312412 308864
rect 312084 308372 312136 308378
rect 312084 308314 312136 308320
rect 312188 308366 312308 308394
rect 311992 308304 312044 308310
rect 311992 308246 312044 308252
rect 312004 274038 312032 308246
rect 312096 287706 312124 308314
rect 312188 290698 312216 308366
rect 312372 307290 312400 308858
rect 312360 307284 312412 307290
rect 312360 307226 312412 307232
rect 312648 302841 312676 310420
rect 312740 310406 312938 310434
rect 312740 308310 312768 310406
rect 313108 308378 313136 310420
rect 313292 310406 313398 310434
rect 313096 308372 313148 308378
rect 313096 308314 313148 308320
rect 312728 308304 312780 308310
rect 312728 308246 312780 308252
rect 313292 308174 313320 310406
rect 313568 308394 313596 310420
rect 313384 308366 313596 308394
rect 313660 310406 313858 310434
rect 313280 308168 313332 308174
rect 313280 308110 313332 308116
rect 313280 307420 313332 307426
rect 313280 307362 313332 307368
rect 312634 302832 312690 302841
rect 312634 302767 312690 302776
rect 312176 290692 312228 290698
rect 312176 290634 312228 290640
rect 312084 287700 312136 287706
rect 312084 287642 312136 287648
rect 311992 274032 312044 274038
rect 311992 273974 312044 273980
rect 313292 273970 313320 307362
rect 313384 275534 313412 308366
rect 313660 308258 313688 310406
rect 313476 308230 313688 308258
rect 313476 289134 313504 308230
rect 313648 308168 313700 308174
rect 313648 308110 313700 308116
rect 313556 308100 313608 308106
rect 313556 308042 313608 308048
rect 313568 290630 313596 308042
rect 313660 305969 313688 308110
rect 314028 307222 314056 310420
rect 314120 310406 314318 310434
rect 314120 307426 314148 310406
rect 314488 308106 314516 310420
rect 314660 308372 314712 308378
rect 314660 308314 314712 308320
rect 314476 308100 314528 308106
rect 314476 308042 314528 308048
rect 314672 307850 314700 308314
rect 314764 308038 314792 310420
rect 314948 308394 314976 310420
rect 314856 308366 314976 308394
rect 315040 310406 315238 310434
rect 314752 308032 314804 308038
rect 314752 307974 314804 307980
rect 314672 307822 314792 307850
rect 314660 307760 314712 307766
rect 314660 307702 314712 307708
rect 314108 307420 314160 307426
rect 314108 307362 314160 307368
rect 314016 307216 314068 307222
rect 314016 307158 314068 307164
rect 313646 305960 313702 305969
rect 313646 305895 313702 305904
rect 313556 290624 313608 290630
rect 313556 290566 313608 290572
rect 313464 289128 313516 289134
rect 313464 289070 313516 289076
rect 313372 275528 313424 275534
rect 313372 275470 313424 275476
rect 313280 273964 313332 273970
rect 313280 273906 313332 273912
rect 311900 263084 311952 263090
rect 311900 263026 311952 263032
rect 310520 246492 310572 246498
rect 310520 246434 310572 246440
rect 314672 246430 314700 307702
rect 314764 246634 314792 307822
rect 314856 275466 314884 308366
rect 315040 308258 315068 310406
rect 315408 308378 315436 310420
rect 315500 310406 315698 310434
rect 315396 308372 315448 308378
rect 315396 308314 315448 308320
rect 314948 308230 315068 308258
rect 314948 290562 314976 308230
rect 315028 308168 315080 308174
rect 315028 308110 315080 308116
rect 315040 292058 315068 308110
rect 315120 308032 315172 308038
rect 315120 307974 315172 307980
rect 315132 304366 315160 307974
rect 315500 307766 315528 310406
rect 315868 308174 315896 310420
rect 316144 308922 316172 310420
rect 316132 308916 316184 308922
rect 316132 308858 316184 308864
rect 316328 308802 316356 310420
rect 316236 308774 316356 308802
rect 316420 310406 316618 310434
rect 316132 308372 316184 308378
rect 316132 308314 316184 308320
rect 316040 308304 316092 308310
rect 316040 308246 316092 308252
rect 315856 308168 315908 308174
rect 315856 308110 315908 308116
rect 315488 307760 315540 307766
rect 315488 307702 315540 307708
rect 315120 304360 315172 304366
rect 315120 304302 315172 304308
rect 315028 292052 315080 292058
rect 315028 291994 315080 292000
rect 314936 290556 314988 290562
rect 314936 290498 314988 290504
rect 314844 275460 314896 275466
rect 314844 275402 314896 275408
rect 316052 250617 316080 308246
rect 316144 264450 316172 308314
rect 316236 275398 316264 308774
rect 316420 308310 316448 310406
rect 316788 308378 316816 310420
rect 316880 310406 317078 310434
rect 316776 308372 316828 308378
rect 316776 308314 316828 308320
rect 316408 308304 316460 308310
rect 316408 308246 316460 308252
rect 316880 308156 316908 310406
rect 317052 308916 317104 308922
rect 317052 308858 317104 308864
rect 317064 308174 317092 308858
rect 316328 308128 316908 308156
rect 317052 308168 317104 308174
rect 316328 276894 316356 308128
rect 317052 308110 317104 308116
rect 317248 296714 317276 310420
rect 317420 308916 317472 308922
rect 317420 308858 317472 308864
rect 316420 296686 317276 296714
rect 316420 290494 316448 296686
rect 316408 290488 316460 290494
rect 316408 290430 316460 290436
rect 316316 276888 316368 276894
rect 316316 276830 316368 276836
rect 316224 275392 316276 275398
rect 316224 275334 316276 275340
rect 316132 264444 316184 264450
rect 316132 264386 316184 264392
rect 316038 250608 316094 250617
rect 316038 250543 316094 250552
rect 317432 249286 317460 308858
rect 317524 308310 317552 310420
rect 317708 308394 317736 310420
rect 317800 310406 317998 310434
rect 317800 308922 317828 310406
rect 317788 308916 317840 308922
rect 317788 308858 317840 308864
rect 318168 308394 318196 310420
rect 317616 308366 317736 308394
rect 317800 308366 318196 308394
rect 318260 310406 318458 310434
rect 317512 308304 317564 308310
rect 317512 308246 317564 308252
rect 317512 307556 317564 307562
rect 317512 307498 317564 307504
rect 317524 252074 317552 307498
rect 317616 269822 317644 308366
rect 317696 308236 317748 308242
rect 317696 308178 317748 308184
rect 317708 275330 317736 308178
rect 317800 282402 317828 308366
rect 317880 308304 317932 308310
rect 317880 308246 317932 308252
rect 317892 301646 317920 308246
rect 318260 308242 318288 310406
rect 318248 308236 318300 308242
rect 318248 308178 318300 308184
rect 318064 308168 318116 308174
rect 318064 308110 318116 308116
rect 317880 301640 317932 301646
rect 317880 301582 317932 301588
rect 317788 282396 317840 282402
rect 317788 282338 317840 282344
rect 317696 275324 317748 275330
rect 317696 275266 317748 275272
rect 317604 269816 317656 269822
rect 317604 269758 317656 269764
rect 318076 254726 318104 308110
rect 318628 307562 318656 310420
rect 318800 308984 318852 308990
rect 318800 308926 318852 308932
rect 318616 307556 318668 307562
rect 318616 307498 318668 307504
rect 318064 254720 318116 254726
rect 318064 254662 318116 254668
rect 317512 252068 317564 252074
rect 317512 252010 317564 252016
rect 318812 252006 318840 308926
rect 318904 308310 318932 310420
rect 318984 308916 319036 308922
rect 318984 308858 319036 308864
rect 318892 308304 318944 308310
rect 318892 308246 318944 308252
rect 318892 308168 318944 308174
rect 318892 308110 318944 308116
rect 318800 252000 318852 252006
rect 318800 251942 318852 251948
rect 318904 251938 318932 308110
rect 318996 265878 319024 308858
rect 319088 267238 319116 310420
rect 319180 310406 319378 310434
rect 319180 308990 319208 310406
rect 319168 308984 319220 308990
rect 319168 308926 319220 308932
rect 319548 308922 319576 310420
rect 319536 308916 319588 308922
rect 319536 308858 319588 308864
rect 319732 308394 319760 310420
rect 319180 308366 319760 308394
rect 319824 310406 320022 310434
rect 320206 310406 320312 310434
rect 319180 276826 319208 308366
rect 319260 308304 319312 308310
rect 319260 308246 319312 308252
rect 319272 285190 319300 308246
rect 319824 308174 319852 310406
rect 320180 308916 320232 308922
rect 320180 308858 320232 308864
rect 319812 308168 319864 308174
rect 319812 308110 319864 308116
rect 319260 285184 319312 285190
rect 319260 285126 319312 285132
rect 319168 276820 319220 276826
rect 319168 276762 319220 276768
rect 319076 267232 319128 267238
rect 319076 267174 319128 267180
rect 318984 265872 319036 265878
rect 318984 265814 319036 265820
rect 318892 251932 318944 251938
rect 318892 251874 318944 251880
rect 320192 251870 320220 308858
rect 320284 256222 320312 310406
rect 320468 308360 320496 310420
rect 320652 308922 320680 310420
rect 320744 310406 320942 310434
rect 320640 308916 320692 308922
rect 320640 308858 320692 308864
rect 320468 308332 320680 308360
rect 320456 308168 320508 308174
rect 320652 308156 320680 308332
rect 320456 308110 320508 308116
rect 320560 308128 320680 308156
rect 320364 306604 320416 306610
rect 320364 306546 320416 306552
rect 320376 268598 320404 306546
rect 320468 271182 320496 308110
rect 320560 276758 320588 308128
rect 320744 306610 320772 310406
rect 321112 308174 321140 310420
rect 321204 310406 321402 310434
rect 321586 310406 321692 310434
rect 321100 308168 321152 308174
rect 321100 308110 321152 308116
rect 320732 306604 320784 306610
rect 320732 306546 320784 306552
rect 321204 296714 321232 310406
rect 321560 308372 321612 308378
rect 321560 308314 321612 308320
rect 320652 296686 321232 296714
rect 320652 291990 320680 296686
rect 320640 291984 320692 291990
rect 320640 291926 320692 291932
rect 320548 276752 320600 276758
rect 320548 276694 320600 276700
rect 320456 271176 320508 271182
rect 320456 271118 320508 271124
rect 320364 268592 320416 268598
rect 320364 268534 320416 268540
rect 320272 256216 320324 256222
rect 320272 256158 320324 256164
rect 320180 251864 320232 251870
rect 320180 251806 320232 251812
rect 317420 249280 317472 249286
rect 317420 249222 317472 249228
rect 321572 248033 321600 308314
rect 321664 256154 321692 310406
rect 321756 310406 321862 310434
rect 321756 276690 321784 310406
rect 322032 308394 322060 310420
rect 321848 308366 322060 308394
rect 321848 291922 321876 308366
rect 322308 307970 322336 310420
rect 322492 308378 322520 310420
rect 322584 310406 322782 310434
rect 322966 310406 323072 310434
rect 322480 308372 322532 308378
rect 322480 308314 322532 308320
rect 322296 307964 322348 307970
rect 322296 307906 322348 307912
rect 322584 296714 322612 310406
rect 322940 308372 322992 308378
rect 322940 308314 322992 308320
rect 321940 296686 322612 296714
rect 321940 293486 321968 296686
rect 321928 293480 321980 293486
rect 321928 293422 321980 293428
rect 321836 291916 321888 291922
rect 321836 291858 321888 291864
rect 321744 276684 321796 276690
rect 321744 276626 321796 276632
rect 321652 256148 321704 256154
rect 321652 256090 321704 256096
rect 321558 248024 321614 248033
rect 321558 247959 321614 247968
rect 322952 247761 322980 308314
rect 323044 256086 323072 310406
rect 323136 310406 323242 310434
rect 323032 256080 323084 256086
rect 323032 256022 323084 256028
rect 323136 247897 323164 310406
rect 323412 308394 323440 310420
rect 323688 308417 323716 310420
rect 323228 308366 323440 308394
rect 323674 308408 323730 308417
rect 323228 291854 323256 308366
rect 323872 308378 323900 310420
rect 323964 310406 324162 310434
rect 324346 310406 324544 310434
rect 323674 308343 323730 308352
rect 323860 308372 323912 308378
rect 323860 308314 323912 308320
rect 323964 308156 323992 310406
rect 324320 308372 324372 308378
rect 324320 308314 324372 308320
rect 323320 308128 323992 308156
rect 323320 293418 323348 308128
rect 323584 307964 323636 307970
rect 323584 307906 323636 307912
rect 323596 297634 323624 307906
rect 323584 297628 323636 297634
rect 323584 297570 323636 297576
rect 323308 293412 323360 293418
rect 323308 293354 323360 293360
rect 323216 291848 323268 291854
rect 323216 291790 323268 291796
rect 323122 247888 323178 247897
rect 323122 247823 323178 247832
rect 322938 247752 322994 247761
rect 322938 247687 322994 247696
rect 314752 246628 314804 246634
rect 314752 246570 314804 246576
rect 314660 246424 314712 246430
rect 314660 246366 314712 246372
rect 301042 246256 301098 246265
rect 301042 246191 301098 246200
rect 300952 245540 301004 245546
rect 300952 245482 301004 245488
rect 324332 245138 324360 308314
rect 324412 308304 324464 308310
rect 324412 308246 324464 308252
rect 324424 246362 324452 308246
rect 324516 256018 324544 310406
rect 324608 308378 324636 310420
rect 324596 308372 324648 308378
rect 324596 308314 324648 308320
rect 324596 308236 324648 308242
rect 324596 308178 324648 308184
rect 324608 260302 324636 308178
rect 324792 296714 324820 310420
rect 325068 308553 325096 310420
rect 325054 308544 325110 308553
rect 325054 308479 325110 308488
rect 325252 308242 325280 310420
rect 325344 310406 325542 310434
rect 325726 310406 325924 310434
rect 325344 308310 325372 310406
rect 325792 308372 325844 308378
rect 325792 308314 325844 308320
rect 325332 308304 325384 308310
rect 325332 308246 325384 308252
rect 325700 308304 325752 308310
rect 325700 308246 325752 308252
rect 325240 308236 325292 308242
rect 325240 308178 325292 308184
rect 324700 296686 324820 296714
rect 324700 293350 324728 296686
rect 324688 293344 324740 293350
rect 324688 293286 324740 293292
rect 325712 261730 325740 308246
rect 325804 278254 325832 308314
rect 325896 308122 325924 310406
rect 325988 308258 326016 310420
rect 325988 308230 326108 308258
rect 325896 308094 326016 308122
rect 325884 308032 325936 308038
rect 325884 307974 325936 307980
rect 325896 294778 325924 307974
rect 325988 294846 326016 308094
rect 326080 305697 326108 308230
rect 326172 307154 326200 310420
rect 326264 310406 326462 310434
rect 326264 308038 326292 310406
rect 326632 308310 326660 310420
rect 326816 308378 326844 310420
rect 327092 308378 327120 310420
rect 327276 308394 327304 310420
rect 326804 308372 326856 308378
rect 326804 308314 326856 308320
rect 327080 308372 327132 308378
rect 327080 308314 327132 308320
rect 327184 308366 327304 308394
rect 327368 310406 327566 310434
rect 326620 308304 326672 308310
rect 326620 308246 326672 308252
rect 326252 308032 326304 308038
rect 326252 307974 326304 307980
rect 327080 307964 327132 307970
rect 327080 307906 327132 307912
rect 326160 307148 326212 307154
rect 326160 307090 326212 307096
rect 326066 305688 326122 305697
rect 326066 305623 326122 305632
rect 325976 294840 326028 294846
rect 325976 294782 326028 294788
rect 325884 294772 325936 294778
rect 325884 294714 325936 294720
rect 325792 278248 325844 278254
rect 325792 278190 325844 278196
rect 325700 261724 325752 261730
rect 325700 261666 325752 261672
rect 327092 261594 327120 307906
rect 327184 261662 327212 308366
rect 327264 308304 327316 308310
rect 327264 308246 327316 308252
rect 327276 278118 327304 308246
rect 327368 278186 327396 310406
rect 327448 308372 327500 308378
rect 327448 308314 327500 308320
rect 327460 294710 327488 308314
rect 327736 296714 327764 310420
rect 327828 310406 328026 310434
rect 327828 307970 327856 310406
rect 328196 308310 328224 310420
rect 328472 308922 328500 310420
rect 328460 308916 328512 308922
rect 328460 308858 328512 308864
rect 328656 308394 328684 310420
rect 328472 308366 328684 308394
rect 328748 310406 328946 310434
rect 328184 308304 328236 308310
rect 328184 308246 328236 308252
rect 327816 307964 327868 307970
rect 327816 307906 327868 307912
rect 327552 296686 327764 296714
rect 327552 296206 327580 296686
rect 327540 296200 327592 296206
rect 327540 296142 327592 296148
rect 327448 294704 327500 294710
rect 327448 294646 327500 294652
rect 327356 278180 327408 278186
rect 327356 278122 327408 278128
rect 327264 278112 327316 278118
rect 327264 278054 327316 278060
rect 328472 262954 328500 308366
rect 328552 308304 328604 308310
rect 328748 308258 328776 310406
rect 328828 308916 328880 308922
rect 328828 308858 328880 308864
rect 328552 308246 328604 308252
rect 328564 263022 328592 308246
rect 328656 308230 328776 308258
rect 328656 279682 328684 308230
rect 328736 308168 328788 308174
rect 328736 308110 328788 308116
rect 328644 279676 328696 279682
rect 328644 279618 328696 279624
rect 328748 279614 328776 308110
rect 328840 293282 328868 308858
rect 329116 296714 329144 310420
rect 329208 310406 329406 310434
rect 329208 308310 329236 310406
rect 329196 308304 329248 308310
rect 329196 308246 329248 308252
rect 329576 308174 329604 310420
rect 329852 308394 329880 310420
rect 330050 310406 330248 310434
rect 329852 308366 330064 308394
rect 329840 308304 329892 308310
rect 329840 308246 329892 308252
rect 329564 308168 329616 308174
rect 329564 308110 329616 308116
rect 328932 296686 329144 296714
rect 328932 296138 328960 296686
rect 328920 296132 328972 296138
rect 328920 296074 328972 296080
rect 328828 293276 328880 293282
rect 328828 293218 328880 293224
rect 328736 279608 328788 279614
rect 328736 279550 328788 279556
rect 329852 279546 329880 308246
rect 329932 308236 329984 308242
rect 329932 308178 329984 308184
rect 329944 281042 329972 308178
rect 330036 296070 330064 308366
rect 330116 308372 330168 308378
rect 330116 308314 330168 308320
rect 330128 297566 330156 308314
rect 330220 305833 330248 310406
rect 330312 308310 330340 310420
rect 330496 308378 330524 310420
rect 330484 308372 330536 308378
rect 330484 308314 330536 308320
rect 330300 308304 330352 308310
rect 330300 308246 330352 308252
rect 330772 307086 330800 310420
rect 330956 308242 330984 310420
rect 330944 308236 330996 308242
rect 330944 308178 330996 308184
rect 330760 307080 330812 307086
rect 330760 307022 330812 307028
rect 331232 306134 331260 310420
rect 331416 306320 331444 310420
rect 331324 306292 331444 306320
rect 331508 310406 331706 310434
rect 331220 306128 331272 306134
rect 331220 306070 331272 306076
rect 331220 305992 331272 305998
rect 331220 305934 331272 305940
rect 330206 305824 330262 305833
rect 330206 305759 330262 305768
rect 330116 297560 330168 297566
rect 330116 297502 330168 297508
rect 330024 296064 330076 296070
rect 330024 296006 330076 296012
rect 329932 281036 329984 281042
rect 329932 280978 329984 280984
rect 329840 279540 329892 279546
rect 329840 279482 329892 279488
rect 328552 263016 328604 263022
rect 328552 262958 328604 262964
rect 328460 262948 328512 262954
rect 328460 262890 328512 262896
rect 327172 261656 327224 261662
rect 327172 261598 327224 261604
rect 327080 261588 327132 261594
rect 327080 261530 327132 261536
rect 324596 260296 324648 260302
rect 324596 260238 324648 260244
rect 324504 256012 324556 256018
rect 324504 255954 324556 255960
rect 331232 253434 331260 305934
rect 331324 262886 331352 306292
rect 331404 306196 331456 306202
rect 331404 306138 331456 306144
rect 331416 264382 331444 306138
rect 331508 280974 331536 310406
rect 331588 306332 331640 306338
rect 331588 306274 331640 306280
rect 331496 280968 331548 280974
rect 331496 280910 331548 280916
rect 331600 280906 331628 306274
rect 331680 306128 331732 306134
rect 331680 306070 331732 306076
rect 331692 297498 331720 306070
rect 331876 305998 331904 310420
rect 331968 310406 332166 310434
rect 331968 306202 331996 310406
rect 332336 306338 332364 310420
rect 332324 306332 332376 306338
rect 332612 306320 332640 310420
rect 332810 310406 332916 310434
rect 332784 306332 332836 306338
rect 332612 306292 332732 306320
rect 332324 306274 332376 306280
rect 331956 306196 332008 306202
rect 331956 306138 332008 306144
rect 332600 306196 332652 306202
rect 332600 306138 332652 306144
rect 331864 305992 331916 305998
rect 331864 305934 331916 305940
rect 331680 297492 331732 297498
rect 331680 297434 331732 297440
rect 331588 280900 331640 280906
rect 331588 280842 331640 280848
rect 331404 264376 331456 264382
rect 331404 264318 331456 264324
rect 331312 262880 331364 262886
rect 331312 262822 331364 262828
rect 331220 253428 331272 253434
rect 331220 253370 331272 253376
rect 332612 247625 332640 306138
rect 332704 253366 332732 306292
rect 332784 306274 332836 306280
rect 332692 253360 332744 253366
rect 332692 253302 332744 253308
rect 332796 253298 332824 306274
rect 332888 264314 332916 310406
rect 333072 309134 333100 310420
rect 333072 309106 333192 309134
rect 332968 304224 333020 304230
rect 332968 304166 333020 304172
rect 332876 264308 332928 264314
rect 332876 264250 332928 264256
rect 332980 264246 333008 304166
rect 333164 299474 333192 309106
rect 333256 306338 333284 310420
rect 333348 310406 333546 310434
rect 333244 306332 333296 306338
rect 333244 306274 333296 306280
rect 333348 304230 333376 310406
rect 333716 306202 333744 310420
rect 333704 306196 333756 306202
rect 333704 306138 333756 306144
rect 333336 304224 333388 304230
rect 333336 304166 333388 304172
rect 333072 299446 333192 299474
rect 333072 282334 333100 299446
rect 333900 297430 333928 310420
rect 333992 310406 334190 310434
rect 333888 297424 333940 297430
rect 333888 297366 333940 297372
rect 333060 282328 333112 282334
rect 333060 282270 333112 282276
rect 332968 264240 333020 264246
rect 332968 264182 333020 264188
rect 333992 260234 334020 310406
rect 334164 306400 334216 306406
rect 334164 306342 334216 306348
rect 334072 306332 334124 306338
rect 334072 306274 334124 306280
rect 334084 265674 334112 306274
rect 334176 282198 334204 306342
rect 334360 306320 334388 310420
rect 334268 306292 334388 306320
rect 334452 310406 334650 310434
rect 334268 282266 334296 306292
rect 334452 302234 334480 310406
rect 334820 306338 334848 310420
rect 334912 310406 335110 310434
rect 334912 306406 334940 310406
rect 334900 306400 334952 306406
rect 334900 306342 334952 306348
rect 334808 306332 334860 306338
rect 334808 306274 334860 306280
rect 334360 302206 334480 302234
rect 334360 283830 334388 302206
rect 335280 298926 335308 310420
rect 335452 306400 335504 306406
rect 335452 306342 335504 306348
rect 335360 306332 335412 306338
rect 335360 306274 335412 306280
rect 335268 298920 335320 298926
rect 335268 298862 335320 298868
rect 334348 283824 334400 283830
rect 334348 283766 334400 283772
rect 334256 282260 334308 282266
rect 334256 282202 334308 282208
rect 334164 282192 334216 282198
rect 334164 282134 334216 282140
rect 334072 265668 334124 265674
rect 334072 265610 334124 265616
rect 333980 260228 334032 260234
rect 333980 260170 334032 260176
rect 332784 253292 332836 253298
rect 332784 253234 332836 253240
rect 335372 249082 335400 306274
rect 335464 249150 335492 306342
rect 335556 305946 335584 310420
rect 335740 306406 335768 310420
rect 335832 310406 336030 310434
rect 335728 306400 335780 306406
rect 335728 306342 335780 306348
rect 335728 305992 335780 305998
rect 335556 305918 335676 305946
rect 335728 305934 335780 305940
rect 335544 305856 335596 305862
rect 335544 305798 335596 305804
rect 335556 265742 335584 305798
rect 335648 265810 335676 305918
rect 335740 298790 335768 305934
rect 335832 298858 335860 310406
rect 336200 305862 336228 310420
rect 336292 310406 336490 310434
rect 336292 306338 336320 310406
rect 336280 306332 336332 306338
rect 336280 306274 336332 306280
rect 336660 305998 336688 310420
rect 336936 306746 336964 310420
rect 336924 306740 336976 306746
rect 336924 306682 336976 306688
rect 337120 306626 337148 310420
rect 336752 306598 337148 306626
rect 337212 310406 337410 310434
rect 336648 305992 336700 305998
rect 336648 305934 336700 305940
rect 336188 305856 336240 305862
rect 336188 305798 336240 305804
rect 335820 298852 335872 298858
rect 335820 298794 335872 298800
rect 335728 298784 335780 298790
rect 335728 298726 335780 298732
rect 335636 265804 335688 265810
rect 335636 265746 335688 265752
rect 335544 265736 335596 265742
rect 335544 265678 335596 265684
rect 336752 249218 336780 306598
rect 336924 306468 336976 306474
rect 336924 306410 336976 306416
rect 336832 306400 336884 306406
rect 336832 306342 336884 306348
rect 336844 250481 336872 306342
rect 336936 261526 336964 306410
rect 337016 306332 337068 306338
rect 337016 306274 337068 306280
rect 337028 267102 337056 306274
rect 337108 303340 337160 303346
rect 337108 303282 337160 303288
rect 337120 278050 337148 303282
rect 337212 300286 337240 310406
rect 337580 306338 337608 310420
rect 337672 310406 337870 310434
rect 337568 306332 337620 306338
rect 337568 306274 337620 306280
rect 337672 303346 337700 310406
rect 338040 306406 338068 310420
rect 338132 310406 338330 310434
rect 338028 306400 338080 306406
rect 338028 306342 338080 306348
rect 337660 303340 337712 303346
rect 337660 303282 337712 303288
rect 337200 300280 337252 300286
rect 337200 300222 337252 300228
rect 337108 278044 337160 278050
rect 337108 277986 337160 277992
rect 337016 267096 337068 267102
rect 337016 267038 337068 267044
rect 338132 267034 338160 310406
rect 338212 306332 338264 306338
rect 338500 306320 338528 310420
rect 338212 306274 338264 306280
rect 338316 306292 338528 306320
rect 338592 310406 338790 310434
rect 338224 267170 338252 306274
rect 338316 283694 338344 306292
rect 338396 306196 338448 306202
rect 338396 306138 338448 306144
rect 338304 283688 338356 283694
rect 338304 283630 338356 283636
rect 338408 283626 338436 306138
rect 338592 302234 338620 310406
rect 338960 306338 338988 310420
rect 339052 310406 339250 310434
rect 338948 306332 339000 306338
rect 338948 306274 339000 306280
rect 339052 306202 339080 310406
rect 339040 306196 339092 306202
rect 339040 306138 339092 306144
rect 338500 302206 338620 302234
rect 338500 294642 338528 302206
rect 339420 300218 339448 310420
rect 339604 310406 339710 310434
rect 339500 306332 339552 306338
rect 339500 306274 339552 306280
rect 339408 300212 339460 300218
rect 339408 300154 339460 300160
rect 338488 294636 338540 294642
rect 338488 294578 338540 294584
rect 338396 283620 338448 283626
rect 338396 283562 338448 283568
rect 338212 267164 338264 267170
rect 338212 267106 338264 267112
rect 338120 267028 338172 267034
rect 338120 266970 338172 266976
rect 336924 261520 336976 261526
rect 336924 261462 336976 261468
rect 336830 250472 336886 250481
rect 336830 250407 336886 250416
rect 336740 249212 336792 249218
rect 336740 249154 336792 249160
rect 335452 249144 335504 249150
rect 335452 249086 335504 249092
rect 335360 249076 335412 249082
rect 335360 249018 335412 249024
rect 332598 247616 332654 247625
rect 332598 247551 332654 247560
rect 324412 246356 324464 246362
rect 324412 246298 324464 246304
rect 324320 245132 324372 245138
rect 324320 245074 324372 245080
rect 339512 245070 339540 306274
rect 339604 268530 339632 310406
rect 339880 306320 339908 310420
rect 339696 306292 339908 306320
rect 339972 310406 340170 310434
rect 339696 279478 339724 306292
rect 339776 306196 339828 306202
rect 339776 306138 339828 306144
rect 339788 283762 339816 306138
rect 339972 302234 340000 310406
rect 340340 306338 340368 310420
rect 340432 310406 340630 310434
rect 340328 306332 340380 306338
rect 340328 306274 340380 306280
rect 340432 306202 340460 310406
rect 340420 306196 340472 306202
rect 340420 306138 340472 306144
rect 339880 302206 340000 302234
rect 339880 300150 339908 302206
rect 340800 301578 340828 310420
rect 340892 310406 341090 310434
rect 340788 301572 340840 301578
rect 340788 301514 340840 301520
rect 339868 300144 339920 300150
rect 339868 300086 339920 300092
rect 339776 283756 339828 283762
rect 339776 283698 339828 283704
rect 339684 279472 339736 279478
rect 339684 279414 339736 279420
rect 339592 268524 339644 268530
rect 339592 268466 339644 268472
rect 339500 245064 339552 245070
rect 339500 245006 339552 245012
rect 340892 245002 340920 310406
rect 341260 306354 341288 310420
rect 340972 306332 341024 306338
rect 340972 306274 341024 306280
rect 341076 306326 341288 306354
rect 340880 244996 340932 245002
rect 340880 244938 340932 244944
rect 340984 244934 341012 306274
rect 341076 280838 341104 306326
rect 341156 306264 341208 306270
rect 341156 306206 341208 306212
rect 341168 285054 341196 306206
rect 341248 306196 341300 306202
rect 341248 306138 341300 306144
rect 341260 296002 341288 306138
rect 341444 301510 341472 310420
rect 341536 310406 341734 310434
rect 341536 306338 341564 310406
rect 341524 306332 341576 306338
rect 341524 306274 341576 306280
rect 341904 306270 341932 310420
rect 341996 310406 342194 310434
rect 342378 310406 342576 310434
rect 341892 306264 341944 306270
rect 341892 306206 341944 306212
rect 341996 306202 342024 310406
rect 342260 306400 342312 306406
rect 342260 306342 342312 306348
rect 341984 306196 342036 306202
rect 341984 306138 342036 306144
rect 341432 301504 341484 301510
rect 341432 301446 341484 301452
rect 341248 295996 341300 296002
rect 341248 295938 341300 295944
rect 341156 285048 341208 285054
rect 341156 284990 341208 284996
rect 341064 280832 341116 280838
rect 341064 280774 341116 280780
rect 342272 253230 342300 306342
rect 342444 306332 342496 306338
rect 342444 306274 342496 306280
rect 342352 305380 342404 305386
rect 342352 305322 342404 305328
rect 342364 254658 342392 305322
rect 342456 268394 342484 306274
rect 342548 268462 342576 310406
rect 342640 284986 342668 310420
rect 342824 306406 342852 310420
rect 342916 310406 343114 310434
rect 342812 306400 342864 306406
rect 342812 306342 342864 306348
rect 342916 306338 342944 310406
rect 342904 306332 342956 306338
rect 342904 306274 342956 306280
rect 343284 296714 343312 310420
rect 343376 310406 343574 310434
rect 343758 310406 343864 310434
rect 343376 305386 343404 310406
rect 343364 305380 343416 305386
rect 343364 305322 343416 305328
rect 343640 303748 343692 303754
rect 343640 303690 343692 303696
rect 342732 296686 343312 296714
rect 342732 285122 342760 296686
rect 343652 296342 343680 303690
rect 343640 296336 343692 296342
rect 343640 296278 343692 296284
rect 342720 285116 342772 285122
rect 342720 285058 342772 285064
rect 342628 284980 342680 284986
rect 342628 284922 342680 284928
rect 342536 268456 342588 268462
rect 342536 268398 342588 268404
rect 342444 268388 342496 268394
rect 342444 268330 342496 268336
rect 343836 260166 343864 310406
rect 343928 310406 344034 310434
rect 343928 286346 343956 310406
rect 344204 302234 344232 310420
rect 344480 305658 344508 310420
rect 344468 305652 344520 305658
rect 344468 305594 344520 305600
rect 344664 303754 344692 310420
rect 344756 310406 344954 310434
rect 344652 303748 344704 303754
rect 344652 303690 344704 303696
rect 344020 302206 344232 302234
rect 343916 286340 343968 286346
rect 343916 286282 343968 286288
rect 343824 260160 343876 260166
rect 343824 260102 343876 260108
rect 342352 254652 342404 254658
rect 342352 254594 342404 254600
rect 344020 254590 344048 302206
rect 344756 296714 344784 310406
rect 345124 309097 345152 310420
rect 345110 309088 345166 309097
rect 345110 309023 345166 309032
rect 345400 308990 345428 310420
rect 345388 308984 345440 308990
rect 345388 308926 345440 308932
rect 345584 305658 345612 310420
rect 345572 305652 345624 305658
rect 345572 305594 345624 305600
rect 345860 303074 345888 310420
rect 346044 308961 346072 310420
rect 346030 308952 346086 308961
rect 346320 308922 346348 310420
rect 346030 308887 346086 308896
rect 346308 308916 346360 308922
rect 346308 308858 346360 308864
rect 346504 303142 346532 310420
rect 346492 303136 346544 303142
rect 346492 303078 346544 303084
rect 345848 303068 345900 303074
rect 345848 303010 345900 303016
rect 346780 302938 346808 310420
rect 346768 302932 346820 302938
rect 346768 302874 346820 302880
rect 346964 300422 346992 310420
rect 347240 305522 347268 310420
rect 347228 305516 347280 305522
rect 347228 305458 347280 305464
rect 347424 303074 347452 310420
rect 347700 303346 347728 310420
rect 347780 306332 347832 306338
rect 347780 306274 347832 306280
rect 347688 303340 347740 303346
rect 347688 303282 347740 303288
rect 347412 303068 347464 303074
rect 347412 303010 347464 303016
rect 346952 300416 347004 300422
rect 346952 300358 347004 300364
rect 344112 296686 344784 296714
rect 344112 259010 344140 296686
rect 344100 259004 344152 259010
rect 344100 258946 344152 258952
rect 344008 254584 344060 254590
rect 344008 254526 344060 254532
rect 342260 253224 342312 253230
rect 342260 253166 342312 253172
rect 347792 252210 347820 306274
rect 347884 296274 347912 310420
rect 348160 306241 348188 310420
rect 348146 306232 348202 306241
rect 348146 306167 348202 306176
rect 348344 302938 348372 310420
rect 348528 303550 348556 310420
rect 348620 310406 348818 310434
rect 348620 306338 348648 310406
rect 348608 306332 348660 306338
rect 348608 306274 348660 306280
rect 348988 305930 349016 310420
rect 348976 305924 349028 305930
rect 348976 305866 349028 305872
rect 348516 303544 348568 303550
rect 348516 303486 348568 303492
rect 349264 303210 349292 310420
rect 349252 303204 349304 303210
rect 349252 303146 349304 303152
rect 349448 302988 349476 310420
rect 349724 305862 349752 310420
rect 349712 305856 349764 305862
rect 349712 305798 349764 305804
rect 349908 303278 349936 310420
rect 350000 310406 350198 310434
rect 349896 303272 349948 303278
rect 349896 303214 349948 303220
rect 349172 302960 349476 302988
rect 348332 302932 348384 302938
rect 348332 302874 348384 302880
rect 349172 300354 349200 302960
rect 350000 302234 350028 310406
rect 350368 306134 350396 310420
rect 350356 306128 350408 306134
rect 350356 306070 350408 306076
rect 350644 303006 350672 310420
rect 350632 303000 350684 303006
rect 350632 302942 350684 302948
rect 350828 302666 350856 310420
rect 351104 305318 351132 310420
rect 351092 305312 351144 305318
rect 351092 305254 351144 305260
rect 351288 303414 351316 310420
rect 351564 304298 351592 310420
rect 351748 305386 351776 310420
rect 351736 305380 351788 305386
rect 351736 305322 351788 305328
rect 351552 304292 351604 304298
rect 351552 304234 351604 304240
rect 352024 303482 352052 310420
rect 352208 306066 352236 310420
rect 352196 306060 352248 306066
rect 352196 306002 352248 306008
rect 352484 303618 352512 310420
rect 352668 307970 352696 310420
rect 352656 307964 352708 307970
rect 352656 307906 352708 307912
rect 352944 305726 352972 310420
rect 353128 309058 353156 310420
rect 353116 309052 353168 309058
rect 353116 308994 353168 309000
rect 353404 306270 353432 310420
rect 353588 308310 353616 310420
rect 353576 308304 353628 308310
rect 353576 308246 353628 308252
rect 353392 306264 353444 306270
rect 353392 306206 353444 306212
rect 353864 306202 353892 310420
rect 354048 308174 354076 310420
rect 354036 308168 354088 308174
rect 354036 308110 354088 308116
rect 353852 306196 353904 306202
rect 353852 306138 353904 306144
rect 352932 305720 352984 305726
rect 352932 305662 352984 305668
rect 354324 305590 354352 310420
rect 354508 308038 354536 310420
rect 354784 308938 354812 310420
rect 354968 309126 354996 310420
rect 354956 309120 355008 309126
rect 354956 309062 355008 309068
rect 354784 308910 354904 308938
rect 354772 308848 354824 308854
rect 354772 308790 354824 308796
rect 354680 308712 354732 308718
rect 354680 308654 354732 308660
rect 354692 308514 354720 308654
rect 354680 308508 354732 308514
rect 354680 308450 354732 308456
rect 354784 308106 354812 308790
rect 354772 308100 354824 308106
rect 354772 308042 354824 308048
rect 354496 308032 354548 308038
rect 354496 307974 354548 307980
rect 354876 306338 354904 308910
rect 354864 306332 354916 306338
rect 354864 306274 354916 306280
rect 354312 305584 354364 305590
rect 354312 305526 354364 305532
rect 355244 305454 355272 310420
rect 355428 308854 355456 310420
rect 355626 310406 355824 310434
rect 355416 308848 355468 308854
rect 355416 308790 355468 308796
rect 355416 308712 355468 308718
rect 355416 308654 355468 308660
rect 355324 308576 355376 308582
rect 355324 308518 355376 308524
rect 355232 305448 355284 305454
rect 355232 305390 355284 305396
rect 352472 303612 352524 303618
rect 352472 303554 352524 303560
rect 352012 303476 352064 303482
rect 352012 303418 352064 303424
rect 351276 303408 351328 303414
rect 351276 303350 351328 303356
rect 350816 302660 350868 302666
rect 350816 302602 350868 302608
rect 349264 302206 350028 302234
rect 349264 300490 349292 302206
rect 349252 300484 349304 300490
rect 349252 300426 349304 300432
rect 349160 300348 349212 300354
rect 349160 300290 349212 300296
rect 347872 296268 347924 296274
rect 347872 296210 347924 296216
rect 347780 252204 347832 252210
rect 347780 252146 347832 252152
rect 340972 244928 341024 244934
rect 340972 244870 341024 244876
rect 299662 244760 299718 244769
rect 299662 244695 299718 244704
rect 355336 244186 355364 308518
rect 355324 244180 355376 244186
rect 355324 244122 355376 244128
rect 355428 243846 355456 308654
rect 355692 308644 355744 308650
rect 355692 308586 355744 308592
rect 355600 308508 355652 308514
rect 355600 308450 355652 308456
rect 355508 308100 355560 308106
rect 355508 308042 355560 308048
rect 355520 243953 355548 308042
rect 355612 244594 355640 308450
rect 355600 244588 355652 244594
rect 355600 244530 355652 244536
rect 355704 244322 355732 308586
rect 355796 308582 355824 310406
rect 355784 308576 355836 308582
rect 355784 308518 355836 308524
rect 355888 308514 355916 310420
rect 355968 308576 356020 308582
rect 355968 308518 356020 308524
rect 355876 308508 355928 308514
rect 355876 308450 355928 308456
rect 355784 308236 355836 308242
rect 355784 308178 355836 308184
rect 355796 245478 355824 308178
rect 355980 302802 356008 308518
rect 356072 302870 356100 310420
rect 356348 308378 356376 310420
rect 356546 310406 356744 310434
rect 356336 308372 356388 308378
rect 356336 308314 356388 308320
rect 356060 302864 356112 302870
rect 356060 302806 356112 302812
rect 355968 302796 356020 302802
rect 355968 302738 356020 302744
rect 356716 302234 356744 310406
rect 356808 308582 356836 310420
rect 356796 308576 356848 308582
rect 356796 308518 356848 308524
rect 356992 302734 357020 310420
rect 357268 308718 357296 310420
rect 357256 308712 357308 308718
rect 357256 308654 357308 308660
rect 357452 305182 357480 310420
rect 357532 308304 357584 308310
rect 357532 308246 357584 308252
rect 357544 307970 357572 308246
rect 357532 307964 357584 307970
rect 357532 307906 357584 307912
rect 357728 306610 357756 310420
rect 357716 306604 357768 306610
rect 357716 306546 357768 306552
rect 357912 306490 357940 310420
rect 357544 306462 357940 306490
rect 358004 310406 358202 310434
rect 357440 305176 357492 305182
rect 357440 305118 357492 305124
rect 356980 302728 357032 302734
rect 356980 302670 357032 302676
rect 356716 302206 356836 302234
rect 356704 247648 356756 247654
rect 356704 247590 356756 247596
rect 355784 245472 355836 245478
rect 355784 245414 355836 245420
rect 356334 245304 356390 245313
rect 356334 245239 356390 245248
rect 356348 244633 356376 245239
rect 356610 245168 356666 245177
rect 356610 245103 356666 245112
rect 356334 244624 356390 244633
rect 356334 244559 356390 244568
rect 356624 244497 356652 245103
rect 356610 244488 356666 244497
rect 356610 244423 356666 244432
rect 355692 244316 355744 244322
rect 355692 244258 355744 244264
rect 355506 243944 355562 243953
rect 355506 243879 355562 243888
rect 355416 243840 355468 243846
rect 355416 243782 355468 243788
rect 291200 243772 291252 243778
rect 291200 243714 291252 243720
rect 289912 243704 289964 243710
rect 289912 243646 289964 243652
rect 289820 243636 289872 243642
rect 289820 243578 289872 243584
rect 287336 243568 287388 243574
rect 287336 243510 287388 243516
rect 288440 243568 288492 243574
rect 288440 243510 288492 243516
rect 277030 159896 277086 159905
rect 277030 159831 277086 159840
rect 278134 159896 278190 159905
rect 278134 159831 278190 159840
rect 279238 159896 279294 159905
rect 279238 159831 279294 159840
rect 285954 159896 286010 159905
rect 285954 159831 286010 159840
rect 356244 159860 356296 159866
rect 256700 159656 256752 159662
rect 256054 159624 256110 159633
rect 255320 159588 255372 159594
rect 256700 159598 256752 159604
rect 271050 159624 271106 159633
rect 256054 159559 256110 159568
rect 255320 159530 255372 159536
rect 239588 158772 239640 158778
rect 239588 158714 239640 158720
rect 238116 158704 238168 158710
rect 227718 158672 227774 158681
rect 220820 158636 220872 158642
rect 220820 158578 220872 158584
rect 224224 158636 224276 158642
rect 238114 158672 238116 158681
rect 239600 158681 239628 158714
rect 238168 158672 238170 158681
rect 227718 158607 227774 158616
rect 229100 158636 229152 158642
rect 224224 158578 224276 158584
rect 219440 157888 219492 157894
rect 219440 157830 219492 157836
rect 219452 16574 219480 157830
rect 220832 16574 220860 158578
rect 224236 157962 224264 158578
rect 224314 158264 224370 158273
rect 224314 158199 224370 158208
rect 224224 157956 224276 157962
rect 224224 157898 224276 157904
rect 224328 157729 224356 158199
rect 224958 157856 225014 157865
rect 224958 157791 225014 157800
rect 224314 157720 224370 157729
rect 224314 157655 224370 157664
rect 223580 157412 223632 157418
rect 223580 157354 223632 157360
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219348 3732 219400 3738
rect 219348 3674 219400 3680
rect 219268 3602 219388 3618
rect 219268 3596 219400 3602
rect 219268 3590 219348 3596
rect 219348 3538 219400 3544
rect 219346 3496 219402 3505
rect 219084 3454 219296 3482
rect 218058 3431 218114 3440
rect 218072 480 218100 3431
rect 219268 480 219296 3454
rect 219346 3431 219402 3440
rect 219360 3233 219388 3431
rect 219346 3224 219402 3233
rect 219346 3159 219402 3168
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222750 3904 222806 3913
rect 222750 3839 222806 3848
rect 222764 480 222792 3839
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 157354
rect 224972 16574 225000 157791
rect 227732 16574 227760 158607
rect 238114 158607 238170 158616
rect 239586 158672 239642 158681
rect 239586 158607 239642 158616
rect 242438 158672 242494 158681
rect 242438 158607 242494 158616
rect 244278 158672 244334 158681
rect 244278 158607 244334 158616
rect 248326 158672 248382 158681
rect 248326 158607 248382 158616
rect 250902 158672 250958 158681
rect 250902 158607 250958 158616
rect 252098 158672 252154 158681
rect 252098 158607 252154 158616
rect 229100 158578 229152 158584
rect 229112 16574 229140 158578
rect 234620 158568 234672 158574
rect 231858 158536 231914 158545
rect 230480 158500 230532 158506
rect 234620 158510 234672 158516
rect 231858 158471 231914 158480
rect 230480 158442 230532 158448
rect 230492 16574 230520 158442
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 225156 480 225184 16546
rect 227534 3768 227590 3777
rect 227534 3703 227590 3712
rect 226338 3632 226394 3641
rect 226338 3567 226394 3576
rect 226352 480 226380 3567
rect 227548 480 227576 3703
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 158471
rect 233238 158400 233294 158409
rect 233238 158335 233294 158344
rect 233252 16574 233280 158335
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11762 234660 158510
rect 238760 158432 238812 158438
rect 238760 158374 238812 158380
rect 240598 158400 240654 158409
rect 234712 158364 234764 158370
rect 234712 158306 234764 158312
rect 234620 11756 234672 11762
rect 234620 11698 234672 11704
rect 234724 6914 234752 158306
rect 237378 158264 237434 158273
rect 237378 158199 237434 158208
rect 237392 16574 237420 158199
rect 238772 16574 238800 158374
rect 240598 158335 240654 158344
rect 240612 155922 240640 158335
rect 241520 158228 241572 158234
rect 241520 158170 241572 158176
rect 240600 155916 240652 155922
rect 240600 155858 240652 155864
rect 241532 16574 241560 158170
rect 242452 157350 242480 158607
rect 242992 158296 243044 158302
rect 242992 158238 243044 158244
rect 242440 157344 242492 157350
rect 242440 157286 242492 157292
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 235816 11756 235868 11762
rect 235816 11698 235868 11704
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11698
rect 237010 3496 237066 3505
rect 237010 3431 237066 3440
rect 237024 480 237052 3431
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240506 3360 240562 3369
rect 240506 3295 240562 3304
rect 240520 480 240548 3295
rect 241716 480 241744 16546
rect 243004 6914 243032 158238
rect 244292 157282 244320 158607
rect 245660 158160 245712 158166
rect 245660 158102 245712 158108
rect 246762 158128 246818 158137
rect 245566 157856 245622 157865
rect 245566 157791 245622 157800
rect 244280 157276 244332 157282
rect 244280 157218 244332 157224
rect 245580 155582 245608 157791
rect 245568 155576 245620 155582
rect 245568 155518 245620 155524
rect 245672 16574 245700 158102
rect 246762 158063 246818 158072
rect 247040 158092 247092 158098
rect 246776 155854 246804 158063
rect 247040 158034 247092 158040
rect 246764 155848 246816 155854
rect 246764 155790 246816 155796
rect 247052 16574 247080 158034
rect 247774 157856 247830 157865
rect 247774 157791 247830 157800
rect 247788 155718 247816 157791
rect 248340 157214 248368 158607
rect 249798 158264 249854 158273
rect 249798 158199 249854 158208
rect 248694 157856 248750 157865
rect 248694 157791 248750 157800
rect 248328 157208 248380 157214
rect 248328 157150 248380 157156
rect 248708 155786 248736 157791
rect 248696 155780 248748 155786
rect 248696 155722 248748 155728
rect 247776 155712 247828 155718
rect 247776 155654 247828 155660
rect 248420 155508 248472 155514
rect 248420 155450 248472 155456
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 245200 3324 245252 3330
rect 245200 3266 245252 3272
rect 244096 3256 244148 3262
rect 244096 3198 244148 3204
rect 244108 480 244136 3198
rect 245212 480 245240 3266
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 155450
rect 249812 16574 249840 158199
rect 250718 157856 250774 157865
rect 250718 157791 250774 157800
rect 250732 155514 250760 157791
rect 250916 157146 250944 158607
rect 251178 157992 251234 158001
rect 251178 157927 251234 157936
rect 250904 157140 250956 157146
rect 250904 157082 250956 157088
rect 250720 155508 250772 155514
rect 250720 155450 250772 155456
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 157927
rect 252112 157078 252140 158607
rect 252560 158024 252612 158030
rect 252560 157966 252612 157972
rect 252100 157072 252152 157078
rect 252100 157014 252152 157020
rect 251272 155644 251324 155650
rect 251272 155586 251324 155592
rect 251284 16574 251312 155586
rect 252572 16574 252600 157966
rect 253478 157856 253534 157865
rect 253478 157791 253534 157800
rect 253492 155650 253520 157791
rect 253480 155644 253532 155650
rect 253480 155586 253532 155592
rect 253940 155440 253992 155446
rect 253940 155382 253992 155388
rect 253952 16574 253980 155382
rect 255332 16574 255360 159530
rect 256068 155446 256096 159559
rect 256056 155440 256108 155446
rect 256056 155382 256108 155388
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 159598
rect 271050 159559 271106 159568
rect 275834 159624 275890 159633
rect 275834 159559 275890 159568
rect 259552 159520 259604 159526
rect 259552 159462 259604 159468
rect 257342 158672 257398 158681
rect 257342 158607 257398 158616
rect 257356 157010 257384 158607
rect 257344 157004 257396 157010
rect 257344 156946 257396 156952
rect 259564 6914 259592 159462
rect 268384 158704 268436 158710
rect 259918 158672 259974 158681
rect 259918 158607 259974 158616
rect 261758 158672 261814 158681
rect 261758 158607 261814 158616
rect 264334 158672 264390 158681
rect 264334 158607 264390 158616
rect 265898 158672 265954 158681
rect 265898 158607 265954 158616
rect 268382 158672 268384 158681
rect 268436 158672 268438 158681
rect 268382 158607 268438 158616
rect 268750 158672 268806 158681
rect 268750 158607 268752 158616
rect 259932 156874 259960 158607
rect 261206 157584 261262 157593
rect 261206 157519 261262 157528
rect 259920 156868 259972 156874
rect 259920 156810 259972 156816
rect 260838 155816 260894 155825
rect 260838 155751 260894 155760
rect 260852 16574 260880 155751
rect 261220 154562 261248 157519
rect 261772 156942 261800 158607
rect 263690 157584 263746 157593
rect 263690 157519 263746 157528
rect 261760 156936 261812 156942
rect 261760 156878 261812 156884
rect 263598 155680 263654 155689
rect 263598 155615 263654 155624
rect 261208 154556 261260 154562
rect 261208 154498 261260 154504
rect 263612 16574 263640 155615
rect 263704 154494 263732 157519
rect 264348 156806 264376 158607
rect 264336 156800 264388 156806
rect 264336 156742 264388 156748
rect 265912 156738 265940 158607
rect 268804 158607 268806 158616
rect 269854 158672 269910 158681
rect 269854 158607 269910 158616
rect 268752 158578 268804 158584
rect 269868 158098 269896 158607
rect 269856 158092 269908 158098
rect 269856 158034 269908 158040
rect 266634 157720 266690 157729
rect 266634 157655 266690 157664
rect 265990 157584 266046 157593
rect 265990 157519 266046 157528
rect 265900 156732 265952 156738
rect 265900 156674 265952 156680
rect 264978 155952 265034 155961
rect 264978 155887 265034 155896
rect 263692 154488 263744 154494
rect 263692 154430 263744 154436
rect 260852 16546 261800 16574
rect 263612 16546 264192 16574
rect 259472 6886 259592 6914
rect 258264 3392 258316 3398
rect 258264 3334 258316 3340
rect 258276 480 258304 3334
rect 259472 480 259500 6886
rect 260656 4140 260708 4146
rect 260656 4082 260708 4088
rect 260668 480 260696 4082
rect 261772 480 261800 16546
rect 262956 4004 263008 4010
rect 262956 3946 263008 3952
rect 262968 480 262996 3946
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 155887
rect 266004 154426 266032 157519
rect 266648 155378 266676 157655
rect 271064 156670 271092 159559
rect 273352 158908 273404 158914
rect 273352 158850 273404 158856
rect 273364 158681 273392 158850
rect 275848 158846 275876 159559
rect 277044 159050 277072 159831
rect 277032 159044 277084 159050
rect 277032 158986 277084 158992
rect 278148 158982 278176 159831
rect 279252 159118 279280 159831
rect 284392 159452 284444 159458
rect 284392 159394 284444 159400
rect 281540 159384 281592 159390
rect 281540 159326 281592 159332
rect 279240 159112 279292 159118
rect 279240 159054 279292 159060
rect 278136 158976 278188 158982
rect 278136 158918 278188 158924
rect 275836 158840 275888 158846
rect 275836 158782 275888 158788
rect 274456 158772 274508 158778
rect 274456 158714 274508 158720
rect 274468 158681 274496 158714
rect 271142 158672 271198 158681
rect 271142 158607 271198 158616
rect 272246 158672 272302 158681
rect 272246 158607 272302 158616
rect 273350 158672 273406 158681
rect 273350 158607 273406 158616
rect 274454 158672 274510 158681
rect 274454 158607 274510 158616
rect 276110 158672 276166 158681
rect 276110 158607 276166 158616
rect 281078 158672 281134 158681
rect 281078 158607 281134 158616
rect 271156 158302 271184 158607
rect 272260 158574 272288 158607
rect 272248 158568 272300 158574
rect 272248 158510 272300 158516
rect 271144 158296 271196 158302
rect 271144 158238 271196 158244
rect 273718 157720 273774 157729
rect 273718 157655 273774 157664
rect 271052 156664 271104 156670
rect 271052 156606 271104 156612
rect 267738 155544 267794 155553
rect 267738 155479 267794 155488
rect 266360 155372 266412 155378
rect 266360 155314 266412 155320
rect 266636 155372 266688 155378
rect 266636 155314 266688 155320
rect 265992 154420 266044 154426
rect 265992 154362 266044 154368
rect 266372 16574 266400 155314
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 155479
rect 273732 155310 273760 157655
rect 276124 156602 276152 158607
rect 278502 157720 278558 157729
rect 278502 157655 278558 157664
rect 276112 156596 276164 156602
rect 276112 156538 276164 156544
rect 274638 155408 274694 155417
rect 274638 155343 274694 155352
rect 270500 155304 270552 155310
rect 267830 155272 267886 155281
rect 270500 155246 270552 155252
rect 273720 155304 273772 155310
rect 273720 155246 273772 155252
rect 267830 155207 267886 155216
rect 267844 16574 267872 155207
rect 269120 152584 269172 152590
rect 269120 152526 269172 152532
rect 269132 16574 269160 152526
rect 270512 16574 270540 155246
rect 273260 152516 273312 152522
rect 273260 152458 273312 152464
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 272444 480 272472 3810
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 152458
rect 274652 16574 274680 155343
rect 278516 155242 278544 157655
rect 277400 155236 277452 155242
rect 277400 155178 277452 155184
rect 278504 155236 278556 155242
rect 278504 155178 278556 155184
rect 277412 16574 277440 155178
rect 281092 155174 281120 158607
rect 278780 155168 278832 155174
rect 278780 155110 278832 155116
rect 281080 155168 281132 155174
rect 281080 155110 281132 155116
rect 278792 16574 278820 155110
rect 274652 16546 274864 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 274836 480 274864 16546
rect 276020 4072 276072 4078
rect 276020 4014 276072 4020
rect 276032 480 276060 4014
rect 277124 3936 277176 3942
rect 277124 3878 277176 3884
rect 277136 480 277164 3878
rect 278332 480 278360 16546
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 280724 480 280752 3742
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 159326
rect 283654 158672 283710 158681
rect 283654 158607 283710 158616
rect 283668 156534 283696 158607
rect 283656 156528 283708 156534
rect 283656 156470 283708 156476
rect 282920 155032 282972 155038
rect 282920 154974 282972 154980
rect 282932 16574 282960 154974
rect 284404 16574 284432 159394
rect 285968 159254 285996 159831
rect 356244 159802 356296 159808
rect 291014 159624 291070 159633
rect 291014 159559 291070 159568
rect 317696 159588 317748 159594
rect 285956 159248 286008 159254
rect 285956 159190 286008 159196
rect 291028 159186 291056 159559
rect 317696 159530 317748 159536
rect 314660 159520 314712 159526
rect 314660 159462 314712 159468
rect 307852 159452 307904 159458
rect 307852 159394 307904 159400
rect 292580 159384 292632 159390
rect 292580 159326 292632 159332
rect 291016 159180 291068 159186
rect 291016 159122 291068 159128
rect 292592 158574 292620 159326
rect 293590 158672 293646 158681
rect 293590 158607 293646 158616
rect 295982 158672 296038 158681
rect 295982 158607 296038 158616
rect 298558 158672 298614 158681
rect 298558 158607 298614 158616
rect 301042 158672 301098 158681
rect 301042 158607 301098 158616
rect 303526 158672 303582 158681
rect 303526 158607 303582 158616
rect 306102 158672 306158 158681
rect 306102 158607 306158 158616
rect 292580 158568 292632 158574
rect 292580 158510 292632 158516
rect 293604 158030 293632 158607
rect 293592 158024 293644 158030
rect 293592 157966 293644 157972
rect 288254 157584 288310 157593
rect 288254 157519 288310 157528
rect 288268 155106 288296 157519
rect 295996 156466 296024 158607
rect 298572 158574 298600 158607
rect 298560 158568 298612 158574
rect 298560 158510 298612 158516
rect 301056 158506 301084 158607
rect 301044 158500 301096 158506
rect 301044 158442 301096 158448
rect 303540 158438 303568 158607
rect 303528 158432 303580 158438
rect 303528 158374 303580 158380
rect 306116 158370 306144 158607
rect 306104 158364 306156 158370
rect 306104 158306 306156 158312
rect 307864 158302 307892 159394
rect 308678 158672 308734 158681
rect 308678 158607 308734 158616
rect 311070 158672 311126 158681
rect 311070 158607 311126 158616
rect 313462 158672 313518 158681
rect 313462 158607 313518 158616
rect 308692 158302 308720 158607
rect 307852 158296 307904 158302
rect 307852 158238 307904 158244
rect 308680 158296 308732 158302
rect 308680 158238 308732 158244
rect 311084 158234 311112 158607
rect 311072 158228 311124 158234
rect 311072 158170 311124 158176
rect 313476 158166 313504 158607
rect 313464 158160 313516 158166
rect 313464 158102 313516 158108
rect 314672 158098 314700 159462
rect 315854 158672 315910 158681
rect 315854 158607 315910 158616
rect 315868 158098 315896 158607
rect 314660 158092 314712 158098
rect 314660 158034 314712 158040
rect 315856 158092 315908 158098
rect 315856 158034 315908 158040
rect 317708 158030 317736 159530
rect 355324 159316 355376 159322
rect 355324 159258 355376 159264
rect 355336 158982 355364 159258
rect 355324 158976 355376 158982
rect 355324 158918 355376 158924
rect 355416 158976 355468 158982
rect 355416 158918 355468 158924
rect 355428 158778 355456 158918
rect 355416 158772 355468 158778
rect 355416 158714 355468 158720
rect 355508 158772 355560 158778
rect 355508 158714 355560 158720
rect 318614 158672 318670 158681
rect 318614 158607 318670 158616
rect 321006 158672 321062 158681
rect 321006 158607 321062 158616
rect 323398 158672 323454 158681
rect 323398 158607 323454 158616
rect 325974 158672 326030 158681
rect 325974 158607 326030 158616
rect 318628 158030 318656 158607
rect 317696 158024 317748 158030
rect 317696 157966 317748 157972
rect 318616 158024 318668 158030
rect 318616 157966 318668 157972
rect 321020 157962 321048 158607
rect 321008 157956 321060 157962
rect 321008 157898 321060 157904
rect 323412 157894 323440 158607
rect 323400 157888 323452 157894
rect 323400 157830 323452 157836
rect 325988 157826 326016 158607
rect 355520 157865 355548 158714
rect 356256 158574 356284 159802
rect 356244 158568 356296 158574
rect 356244 158510 356296 158516
rect 355506 157856 355562 157865
rect 325976 157820 326028 157826
rect 355506 157791 355562 157800
rect 325976 157762 326028 157768
rect 295984 156460 296036 156466
rect 295984 156402 296036 156408
rect 285680 155100 285732 155106
rect 285680 155042 285732 155048
rect 288256 155100 288308 155106
rect 288256 155042 288308 155048
rect 285692 16574 285720 155042
rect 282932 16546 283144 16574
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 283116 480 283144 16546
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 284312 480 284340 3606
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 307944 9648 307996 9654
rect 307944 9590 307996 9596
rect 306748 9580 306800 9586
rect 306748 9522 306800 9528
rect 305552 9512 305604 9518
rect 305552 9454 305604 9460
rect 304356 9444 304408 9450
rect 304356 9386 304408 9392
rect 299664 9376 299716 9382
rect 299664 9318 299716 9324
rect 297272 9308 297324 9314
rect 297272 9250 297324 9256
rect 296076 9104 296128 9110
rect 296076 9046 296128 9052
rect 294880 9036 294932 9042
rect 294880 8978 294932 8984
rect 293684 8968 293736 8974
rect 293684 8910 293736 8916
rect 292580 6180 292632 6186
rect 292580 6122 292632 6128
rect 287796 3732 287848 3738
rect 287796 3674 287848 3680
rect 287808 480 287836 3674
rect 288992 3596 289044 3602
rect 288992 3538 289044 3544
rect 289004 480 289032 3538
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 290188 3460 290240 3466
rect 290188 3402 290240 3408
rect 290200 480 290228 3402
rect 291396 480 291424 3470
rect 292592 480 292620 6122
rect 293696 480 293724 8910
rect 294892 480 294920 8978
rect 296088 480 296116 9046
rect 297284 480 297312 9250
rect 298468 9172 298520 9178
rect 298468 9114 298520 9120
rect 298480 480 298508 9114
rect 299676 480 299704 9318
rect 301964 9240 302016 9246
rect 301964 9182 302016 9188
rect 300768 8900 300820 8906
rect 300768 8842 300820 8848
rect 300780 480 300808 8842
rect 301976 480 302004 9182
rect 303160 8832 303212 8838
rect 303160 8774 303212 8780
rect 303172 480 303200 8774
rect 304368 480 304396 9386
rect 305564 480 305592 9454
rect 306760 480 306788 9522
rect 307956 480 307984 9590
rect 319718 8936 319774 8945
rect 319718 8871 319774 8880
rect 316224 8764 316276 8770
rect 316224 8706 316276 8712
rect 313832 6588 313884 6594
rect 313832 6530 313884 6536
rect 312636 6452 312688 6458
rect 312636 6394 312688 6400
rect 311440 6384 311492 6390
rect 311440 6326 311492 6332
rect 310244 6316 310296 6322
rect 310244 6258 310296 6264
rect 309048 6248 309100 6254
rect 309048 6190 309100 6196
rect 309060 480 309088 6190
rect 310256 480 310284 6258
rect 311452 480 311480 6326
rect 312648 480 312676 6394
rect 313844 480 313872 6530
rect 315028 6520 315080 6526
rect 315028 6462 315080 6468
rect 315040 480 315068 6462
rect 316236 480 316264 8706
rect 317328 6792 317380 6798
rect 317328 6734 317380 6740
rect 317340 480 317368 6734
rect 318524 6656 318576 6662
rect 318524 6598 318576 6604
rect 318536 480 318564 6598
rect 319732 480 319760 8871
rect 323308 6860 323360 6866
rect 323308 6802 323360 6808
rect 320916 6724 320968 6730
rect 320916 6666 320968 6672
rect 320928 480 320956 6666
rect 322112 3460 322164 3466
rect 322112 3402 322164 3408
rect 322124 480 322152 3402
rect 323320 480 323348 6802
rect 350446 6760 350502 6769
rect 350446 6695 350502 6704
rect 348054 6624 348110 6633
rect 348054 6559 348110 6568
rect 344558 6488 344614 6497
rect 344558 6423 344614 6432
rect 340970 6352 341026 6361
rect 340970 6287 341026 6296
rect 337474 6216 337530 6225
rect 337474 6151 337530 6160
rect 326804 6112 326856 6118
rect 326804 6054 326856 6060
rect 325608 3664 325660 3670
rect 325608 3606 325660 3612
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 324424 480 324452 3470
rect 325620 480 325648 3606
rect 326816 480 326844 6054
rect 330392 6044 330444 6050
rect 330392 5986 330444 5992
rect 329196 3596 329248 3602
rect 329196 3538 329248 3544
rect 327998 3360 328054 3369
rect 327998 3295 328054 3304
rect 328012 480 328040 3295
rect 329208 480 329236 3538
rect 330404 480 330432 5986
rect 333888 5976 333940 5982
rect 333888 5918 333940 5924
rect 332692 3732 332744 3738
rect 332692 3674 332744 3680
rect 331586 3496 331642 3505
rect 331586 3431 331642 3440
rect 331600 480 331628 3431
rect 332704 480 332732 3674
rect 333900 480 333928 5918
rect 336280 3800 336332 3806
rect 336280 3742 336332 3748
rect 335082 3632 335138 3641
rect 335082 3567 335138 3576
rect 335096 480 335124 3567
rect 336292 480 336320 3742
rect 337488 480 337516 6151
rect 339868 3868 339920 3874
rect 339868 3810 339920 3816
rect 338670 3768 338726 3777
rect 338670 3703 338726 3712
rect 338684 480 338712 3703
rect 339880 480 339908 3810
rect 340984 480 341012 6287
rect 342168 4004 342220 4010
rect 342168 3946 342220 3952
rect 342180 480 342208 3946
rect 343364 3936 343416 3942
rect 343364 3878 343416 3884
rect 343376 480 343404 3878
rect 344572 480 344600 6423
rect 346952 4072 347004 4078
rect 345754 4040 345810 4049
rect 346952 4014 347004 4020
rect 345754 3975 345810 3984
rect 345768 480 345796 3975
rect 346964 480 346992 4014
rect 348068 480 348096 6559
rect 349250 3224 349306 3233
rect 349250 3159 349306 3168
rect 349264 480 349292 3159
rect 350460 480 350488 6695
rect 354036 4140 354088 4146
rect 354036 4082 354088 4088
rect 351642 3904 351698 3913
rect 351642 3839 351698 3848
rect 351656 480 351684 3839
rect 352840 3256 352892 3262
rect 352840 3198 352892 3204
rect 352852 480 352880 3198
rect 354048 480 354076 4082
rect 356242 3768 356298 3777
rect 356242 3703 356298 3712
rect 355508 3596 355560 3602
rect 355508 3538 355560 3544
rect 355232 3392 355284 3398
rect 355232 3334 355284 3340
rect 355244 480 355272 3334
rect 355520 3330 355548 3538
rect 355508 3324 355560 3330
rect 355508 3266 355560 3272
rect 356256 3233 356284 3703
rect 356716 3534 356744 247590
rect 356808 159594 356836 302206
rect 357440 245608 357492 245614
rect 356886 245576 356942 245585
rect 356886 245511 356942 245520
rect 357438 245576 357440 245585
rect 357492 245576 357494 245585
rect 357438 245511 357494 245520
rect 356900 245177 356928 245511
rect 356886 245168 356942 245177
rect 356886 245103 356942 245112
rect 356796 159588 356848 159594
rect 356796 159530 356848 159536
rect 357438 158808 357494 158817
rect 357438 158743 357494 158752
rect 356704 3528 356756 3534
rect 356704 3470 356756 3476
rect 356336 3460 356388 3466
rect 356336 3402 356388 3408
rect 356242 3224 356298 3233
rect 356242 3159 356298 3168
rect 356348 480 356376 3402
rect 357452 3262 357480 158743
rect 357544 158506 357572 306462
rect 358004 306218 358032 310406
rect 358084 308508 358136 308514
rect 358084 308450 358136 308456
rect 358096 308242 358124 308450
rect 358268 308440 358320 308446
rect 358268 308382 358320 308388
rect 358084 308236 358136 308242
rect 358084 308178 358136 308184
rect 358084 306604 358136 306610
rect 358084 306546 358136 306552
rect 357636 306190 358032 306218
rect 357636 158642 357664 306190
rect 358096 306116 358124 306546
rect 357912 306088 358124 306116
rect 357716 305788 357768 305794
rect 357716 305730 357768 305736
rect 357624 158636 357676 158642
rect 357624 158578 357676 158584
rect 357532 158500 357584 158506
rect 357532 158442 357584 158448
rect 357728 158438 357756 305730
rect 357808 305244 357860 305250
rect 357808 305186 357860 305192
rect 357820 159526 357848 305186
rect 357808 159520 357860 159526
rect 357808 159462 357860 159468
rect 357912 158778 357940 306088
rect 357992 305176 358044 305182
rect 357992 305118 358044 305124
rect 358004 159866 358032 305118
rect 358176 245540 358228 245546
rect 358176 245482 358228 245488
rect 358188 245449 358216 245482
rect 358174 245440 358230 245449
rect 358084 245404 358136 245410
rect 358174 245375 358230 245384
rect 358084 245346 358136 245352
rect 357992 159860 358044 159866
rect 357992 159802 358044 159808
rect 357900 158772 357952 158778
rect 357900 158714 357952 158720
rect 357716 158432 357768 158438
rect 357716 158374 357768 158380
rect 358096 3602 358124 245346
rect 358280 245342 358308 308382
rect 358372 305794 358400 310420
rect 358556 310406 358662 310434
rect 358846 310406 359044 310434
rect 358360 305788 358412 305794
rect 358360 305730 358412 305736
rect 358452 305788 358504 305794
rect 358452 305730 358504 305736
rect 358464 305386 358492 305730
rect 358452 305380 358504 305386
rect 358452 305322 358504 305328
rect 358556 305250 358584 310406
rect 358912 306536 358964 306542
rect 358912 306478 358964 306484
rect 358728 306400 358780 306406
rect 358634 306368 358690 306377
rect 358728 306342 358780 306348
rect 358634 306303 358690 306312
rect 358648 306134 358676 306303
rect 358740 306270 358768 306342
rect 358728 306264 358780 306270
rect 358728 306206 358780 306212
rect 358636 306128 358688 306134
rect 358636 306070 358688 306076
rect 358544 305244 358596 305250
rect 358544 305186 358596 305192
rect 358820 251184 358872 251190
rect 358820 251126 358872 251132
rect 358360 247580 358412 247586
rect 358360 247522 358412 247528
rect 358176 245336 358228 245342
rect 358176 245278 358228 245284
rect 358268 245336 358320 245342
rect 358268 245278 358320 245284
rect 358188 6866 358216 245278
rect 358268 243772 358320 243778
rect 358268 243714 358320 243720
rect 358176 6860 358228 6866
rect 358176 6802 358228 6808
rect 358280 6322 358308 243714
rect 358268 6316 358320 6322
rect 358268 6258 358320 6264
rect 358372 3670 358400 247522
rect 358832 6390 358860 251126
rect 358924 158302 358952 306478
rect 359016 306354 359044 310406
rect 359108 306474 359136 310420
rect 359292 306542 359320 310420
rect 359384 310406 359582 310434
rect 359280 306536 359332 306542
rect 359280 306478 359332 306484
rect 359096 306468 359148 306474
rect 359096 306410 359148 306416
rect 359384 306354 359412 310406
rect 359648 308440 359700 308446
rect 359648 308382 359700 308388
rect 359464 306468 359516 306474
rect 359464 306410 359516 306416
rect 359016 306326 359136 306354
rect 359004 302660 359056 302666
rect 359004 302602 359056 302608
rect 358912 158296 358964 158302
rect 358912 158238 358964 158244
rect 359016 158234 359044 302602
rect 359108 158370 359136 306326
rect 359200 306326 359412 306354
rect 359200 159390 359228 306326
rect 359280 305380 359332 305386
rect 359280 305322 359332 305328
rect 359188 159384 359240 159390
rect 359188 159326 359240 159332
rect 359292 158914 359320 305322
rect 359476 296714 359504 306410
rect 359384 296686 359504 296714
rect 359384 159458 359412 296686
rect 359464 245268 359516 245274
rect 359464 245210 359516 245216
rect 359372 159452 359424 159458
rect 359372 159394 359424 159400
rect 359280 158908 359332 158914
rect 359280 158850 359332 158856
rect 359096 158364 359148 158370
rect 359096 158306 359148 158312
rect 359004 158228 359056 158234
rect 359004 158170 359056 158176
rect 359476 6594 359504 245210
rect 359556 243704 359608 243710
rect 359556 243646 359608 243652
rect 359568 9314 359596 243646
rect 359660 158166 359688 308382
rect 359752 302666 359780 310420
rect 359844 310406 360042 310434
rect 359844 305386 359872 310406
rect 360212 308446 360240 310420
rect 360304 310406 360502 310434
rect 360200 308440 360252 308446
rect 360200 308382 360252 308388
rect 360304 307902 360332 310406
rect 360672 308530 360700 310420
rect 360488 308502 360700 308530
rect 360764 310406 360962 310434
rect 360384 308372 360436 308378
rect 360384 308314 360436 308320
rect 360292 307896 360344 307902
rect 360292 307838 360344 307844
rect 360106 306368 360162 306377
rect 360106 306303 360162 306312
rect 360120 306134 360148 306303
rect 360108 306128 360160 306134
rect 360108 306070 360160 306076
rect 359924 306060 359976 306066
rect 359924 306002 359976 306008
rect 359936 305726 359964 306002
rect 359924 305720 359976 305726
rect 359924 305662 359976 305668
rect 360016 305720 360068 305726
rect 360016 305662 360068 305668
rect 359832 305380 359884 305386
rect 359832 305322 359884 305328
rect 360028 305318 360056 305662
rect 360016 305312 360068 305318
rect 360016 305254 360068 305260
rect 359740 302660 359792 302666
rect 359740 302602 359792 302608
rect 360200 250980 360252 250986
rect 360200 250922 360252 250928
rect 359648 158160 359700 158166
rect 359648 158102 359700 158108
rect 359556 9308 359608 9314
rect 359556 9250 359608 9256
rect 359464 6588 359516 6594
rect 359464 6530 359516 6536
rect 360212 6458 360240 250922
rect 360292 250300 360344 250306
rect 360292 250242 360344 250248
rect 360200 6452 360252 6458
rect 360200 6394 360252 6400
rect 358820 6384 358872 6390
rect 358820 6326 358872 6332
rect 360304 6118 360332 250242
rect 360396 158030 360424 308314
rect 360488 158098 360516 308502
rect 360568 307964 360620 307970
rect 360568 307906 360620 307912
rect 360580 159050 360608 307906
rect 360660 307896 360712 307902
rect 360660 307838 360712 307844
rect 360568 159044 360620 159050
rect 360568 158986 360620 158992
rect 360672 158982 360700 307838
rect 360660 158976 360712 158982
rect 360660 158918 360712 158924
rect 360764 158846 360792 310406
rect 361028 308440 361080 308446
rect 361028 308382 361080 308388
rect 360844 247920 360896 247926
rect 360844 247862 360896 247868
rect 360752 158840 360804 158846
rect 360752 158782 360804 158788
rect 360476 158092 360528 158098
rect 360476 158034 360528 158040
rect 360384 158024 360436 158030
rect 360384 157966 360436 157972
rect 360856 6798 360884 247862
rect 360936 243636 360988 243642
rect 360936 243578 360988 243584
rect 360948 8906 360976 243578
rect 361040 157962 361068 308382
rect 361132 308378 361160 310420
rect 361224 310406 361422 310434
rect 361120 308372 361172 308378
rect 361120 308314 361172 308320
rect 361224 307970 361252 310406
rect 361304 308848 361356 308854
rect 361304 308790 361356 308796
rect 361316 308378 361344 308790
rect 361592 308446 361620 310420
rect 361684 310406 361882 310434
rect 361580 308440 361632 308446
rect 361580 308382 361632 308388
rect 361304 308372 361356 308378
rect 361304 308314 361356 308320
rect 361212 307964 361264 307970
rect 361212 307906 361264 307912
rect 361684 307834 361712 310406
rect 362052 308394 362080 310420
rect 361776 308366 362080 308394
rect 362144 310406 362342 310434
rect 361672 307828 361724 307834
rect 361672 307770 361724 307776
rect 361672 248260 361724 248266
rect 361672 248202 361724 248208
rect 361028 157956 361080 157962
rect 361028 157898 361080 157904
rect 360936 8900 360988 8906
rect 360936 8842 360988 8848
rect 360844 6792 360896 6798
rect 360844 6734 360896 6740
rect 360292 6112 360344 6118
rect 360292 6054 360344 6060
rect 358360 3664 358412 3670
rect 358360 3606 358412 3612
rect 358726 3632 358782 3641
rect 358084 3596 358136 3602
rect 358726 3567 358782 3576
rect 358084 3538 358136 3544
rect 357530 3496 357586 3505
rect 357530 3431 357586 3440
rect 357440 3256 357492 3262
rect 357440 3198 357492 3204
rect 357544 480 357572 3431
rect 358740 480 358768 3567
rect 359922 3496 359978 3505
rect 359922 3431 359978 3440
rect 361118 3496 361174 3505
rect 361118 3431 361174 3440
rect 359936 480 359964 3431
rect 361132 480 361160 3431
rect 361684 3330 361712 248202
rect 361776 157894 361804 308366
rect 361948 307828 362000 307834
rect 361948 307770 362000 307776
rect 361856 307760 361908 307766
rect 361856 307702 361908 307708
rect 361764 157888 361816 157894
rect 361764 157830 361816 157836
rect 361868 157826 361896 307702
rect 361960 159322 361988 307770
rect 362144 296714 362172 310406
rect 362406 308816 362462 308825
rect 362406 308751 362462 308760
rect 362420 306374 362448 308751
rect 362512 307766 362540 310420
rect 363694 309088 363750 309097
rect 363694 309023 363750 309032
rect 362500 307760 362552 307766
rect 362500 307702 362552 307708
rect 362420 306346 362540 306374
rect 362408 305516 362460 305522
rect 362408 305458 362460 305464
rect 362052 296686 362172 296714
rect 361948 159316 362000 159322
rect 361948 159258 362000 159264
rect 362052 159118 362080 296686
rect 362132 247852 362184 247858
rect 362132 247794 362184 247800
rect 362040 159112 362092 159118
rect 362040 159054 362092 159060
rect 361856 157820 361908 157826
rect 361856 157762 361908 157768
rect 362144 6526 362172 247794
rect 362316 244316 362368 244322
rect 362316 244258 362368 244264
rect 362224 244180 362276 244186
rect 362224 244122 362276 244128
rect 362132 6520 362184 6526
rect 362132 6462 362184 6468
rect 362236 6186 362264 244122
rect 362328 9382 362356 244258
rect 362420 155582 362448 305458
rect 362408 155576 362460 155582
rect 362408 155518 362460 155524
rect 362316 9376 362368 9382
rect 362316 9318 362368 9324
rect 362224 6180 362276 6186
rect 362224 6122 362276 6128
rect 362512 4010 362540 306346
rect 363144 250912 363196 250918
rect 363144 250854 363196 250860
rect 362960 248328 363012 248334
rect 362960 248270 363012 248276
rect 362500 4004 362552 4010
rect 362500 3946 362552 3952
rect 362972 3942 363000 248270
rect 363052 247512 363104 247518
rect 363052 247454 363104 247460
rect 362960 3936 363012 3942
rect 362960 3878 363012 3884
rect 362314 3496 362370 3505
rect 363064 3466 363092 247454
rect 363156 6050 363184 250854
rect 363236 250436 363288 250442
rect 363236 250378 363288 250384
rect 363248 6225 363276 250378
rect 363328 248396 363380 248402
rect 363328 248338 363380 248344
rect 363340 6769 363368 248338
rect 363512 244588 363564 244594
rect 363512 244530 363564 244536
rect 363418 243944 363474 243953
rect 363418 243879 363474 243888
rect 363326 6760 363382 6769
rect 363326 6695 363382 6704
rect 363432 6662 363460 243879
rect 363524 8838 363552 244530
rect 363604 243568 363656 243574
rect 363604 243510 363656 243516
rect 363616 9042 363644 243510
rect 363708 157457 363736 309023
rect 363786 308952 363842 308961
rect 363786 308887 363842 308896
rect 363800 158545 363828 308887
rect 364996 273222 365024 441662
rect 369216 309120 369268 309126
rect 369216 309062 369268 309068
rect 366456 309052 366508 309058
rect 366456 308994 366508 309000
rect 365810 308680 365866 308689
rect 365810 308615 365866 308624
rect 365076 308032 365128 308038
rect 365076 307974 365128 307980
rect 364984 273216 365036 273222
rect 364984 273158 365036 273164
rect 364708 251116 364760 251122
rect 364708 251058 364760 251064
rect 364616 248192 364668 248198
rect 364616 248134 364668 248140
rect 364340 248124 364392 248130
rect 364340 248066 364392 248072
rect 363786 158536 363842 158545
rect 363786 158471 363842 158480
rect 363694 157448 363750 157457
rect 363694 157383 363750 157392
rect 363604 9036 363656 9042
rect 363604 8978 363656 8984
rect 363512 8832 363564 8838
rect 363512 8774 363564 8780
rect 363420 6656 363472 6662
rect 363420 6598 363472 6604
rect 363234 6216 363290 6225
rect 363234 6151 363290 6160
rect 363144 6044 363196 6050
rect 363144 5986 363196 5992
rect 364352 3738 364380 248066
rect 364524 248056 364576 248062
rect 364524 247998 364576 248004
rect 364432 247988 364484 247994
rect 364432 247930 364484 247936
rect 364444 3874 364472 247930
rect 364432 3868 364484 3874
rect 364432 3810 364484 3816
rect 364536 3806 364564 247998
rect 364628 4078 364656 248134
rect 364720 6361 364748 251058
rect 364800 250844 364852 250850
rect 364800 250786 364852 250792
rect 364706 6352 364762 6361
rect 364706 6287 364762 6296
rect 364812 5982 364840 250786
rect 364892 250708 364944 250714
rect 364892 250650 364944 250656
rect 364904 8770 364932 250650
rect 364984 247716 365036 247722
rect 364984 247658 365036 247664
rect 364996 9110 365024 247658
rect 365088 156874 365116 307974
rect 365168 305448 365220 305454
rect 365168 305390 365220 305396
rect 365180 159254 365208 305390
rect 365720 268660 365772 268666
rect 365720 268602 365772 268608
rect 365258 159624 365314 159633
rect 365258 159559 365314 159568
rect 365168 159248 365220 159254
rect 365168 159190 365220 159196
rect 365076 156868 365128 156874
rect 365076 156810 365128 156816
rect 364984 9104 365036 9110
rect 364984 9046 365036 9052
rect 364892 8764 364944 8770
rect 364892 8706 364944 8712
rect 364800 5976 364852 5982
rect 364800 5918 364852 5924
rect 365272 4146 365300 159559
rect 365260 4140 365312 4146
rect 365260 4082 365312 4088
rect 364616 4072 364668 4078
rect 364616 4014 364668 4020
rect 364524 3800 364576 3806
rect 364524 3742 364576 3748
rect 364340 3732 364392 3738
rect 364340 3674 364392 3680
rect 364614 3632 364670 3641
rect 364614 3567 364670 3576
rect 363510 3496 363566 3505
rect 362314 3431 362370 3440
rect 363052 3460 363104 3466
rect 361672 3324 361724 3330
rect 361672 3266 361724 3272
rect 362328 480 362356 3431
rect 363510 3431 363566 3440
rect 363052 3402 363104 3408
rect 363524 480 363552 3431
rect 364628 480 364656 3567
rect 365732 1290 365760 268602
rect 365824 6730 365852 308615
rect 366272 308304 366324 308310
rect 366272 308246 366324 308252
rect 366180 308168 366232 308174
rect 366180 308110 366232 308116
rect 365996 253496 366048 253502
rect 365996 253438 366048 253444
rect 365904 250368 365956 250374
rect 365904 250310 365956 250316
rect 365812 6724 365864 6730
rect 365812 6666 365864 6672
rect 365810 3632 365866 3641
rect 365810 3567 365866 3576
rect 365720 1284 365772 1290
rect 365720 1226 365772 1232
rect 365824 480 365852 3567
rect 365916 3398 365944 250310
rect 366008 8945 366036 253438
rect 366088 247784 366140 247790
rect 366088 247726 366140 247732
rect 366100 9450 366128 247726
rect 366192 157010 366220 308110
rect 366284 158137 366312 308246
rect 366364 308100 366416 308106
rect 366364 308042 366416 308048
rect 366376 159225 366404 308042
rect 366362 159216 366418 159225
rect 366362 159151 366418 159160
rect 366468 159089 366496 308994
rect 366548 308984 366600 308990
rect 366548 308926 366600 308932
rect 366454 159080 366510 159089
rect 366454 159015 366510 159024
rect 366560 158817 366588 308926
rect 368756 308916 368808 308922
rect 368756 308858 368808 308864
rect 367468 308644 367520 308650
rect 367468 308586 367520 308592
rect 367192 251048 367244 251054
rect 367192 250990 367244 250996
rect 367100 250776 367152 250782
rect 367100 250718 367152 250724
rect 366546 158808 366602 158817
rect 366546 158743 366602 158752
rect 366270 158128 366326 158137
rect 366270 158063 366326 158072
rect 366180 157004 366232 157010
rect 366180 156946 366232 156952
rect 366088 9444 366140 9450
rect 366088 9386 366140 9392
rect 365994 8936 366050 8945
rect 365994 8871 366050 8880
rect 367112 6497 367140 250718
rect 367204 6633 367232 250990
rect 367284 246560 367336 246566
rect 367284 246502 367336 246508
rect 367296 9178 367324 246502
rect 367376 245336 367428 245342
rect 367376 245278 367428 245284
rect 367388 9518 367416 245278
rect 367480 155378 367508 308586
rect 367560 308576 367612 308582
rect 367560 308518 367612 308524
rect 367572 156738 367600 308518
rect 367836 308236 367888 308242
rect 367836 308178 367888 308184
rect 367744 306128 367796 306134
rect 367744 306070 367796 306076
rect 367652 305924 367704 305930
rect 367652 305866 367704 305872
rect 367560 156732 367612 156738
rect 367560 156674 367612 156680
rect 367664 155718 367692 305866
rect 367652 155712 367704 155718
rect 367652 155654 367704 155660
rect 367756 155514 367784 306070
rect 367848 159361 367876 308178
rect 367928 303544 367980 303550
rect 367928 303486 367980 303492
rect 367834 159352 367890 159361
rect 367834 159287 367890 159296
rect 367940 157350 367968 303486
rect 368480 250640 368532 250646
rect 368480 250582 368532 250588
rect 367928 157344 367980 157350
rect 367928 157286 367980 157292
rect 367744 155508 367796 155514
rect 367744 155450 367796 155456
rect 367468 155372 367520 155378
rect 367468 155314 367520 155320
rect 367376 9512 367428 9518
rect 367376 9454 367428 9460
rect 367284 9172 367336 9178
rect 367284 9114 367336 9120
rect 367190 6624 367246 6633
rect 367190 6559 367246 6568
rect 367098 6488 367154 6497
rect 367098 6423 367154 6432
rect 368492 6254 368520 250582
rect 368572 245472 368624 245478
rect 368572 245414 368624 245420
rect 368584 8974 368612 245414
rect 368664 245200 368716 245206
rect 368664 245142 368716 245148
rect 368676 9586 368704 245142
rect 368768 157282 368796 308858
rect 368848 308440 368900 308446
rect 368848 308382 368900 308388
rect 368756 157276 368808 157282
rect 368756 157218 368808 157224
rect 368860 156806 368888 308382
rect 368940 308372 368992 308378
rect 368940 308314 368992 308320
rect 368952 156942 368980 308314
rect 369030 306232 369086 306241
rect 369030 306167 369086 306176
rect 368940 156936 368992 156942
rect 368940 156878 368992 156884
rect 368848 156800 368900 156806
rect 368848 156742 368900 156748
rect 369044 155854 369072 306167
rect 369124 305856 369176 305862
rect 369124 305798 369176 305804
rect 369032 155848 369084 155854
rect 369032 155790 369084 155796
rect 369136 155786 369164 305798
rect 369228 158001 369256 309062
rect 431222 308544 431278 308553
rect 431222 308479 431278 308488
rect 377404 307284 377456 307290
rect 377404 307226 377456 307232
rect 370136 306332 370188 306338
rect 370136 306274 370188 306280
rect 370044 305584 370096 305590
rect 370044 305526 370096 305532
rect 369308 303340 369360 303346
rect 369308 303282 369360 303288
rect 369214 157992 369270 158001
rect 369214 157927 369270 157936
rect 369320 155922 369348 303282
rect 369860 250504 369912 250510
rect 369860 250446 369912 250452
rect 369308 155916 369360 155922
rect 369308 155858 369360 155864
rect 369124 155780 369176 155786
rect 369124 155722 369176 155728
rect 369872 9654 369900 250446
rect 369952 243840 370004 243846
rect 369952 243782 370004 243788
rect 369860 9648 369912 9654
rect 369860 9590 369912 9596
rect 368664 9580 368716 9586
rect 368664 9522 368716 9528
rect 369964 9246 369992 243782
rect 370056 155174 370084 305526
rect 370148 156602 370176 306274
rect 371700 306264 371752 306270
rect 371700 306206 371752 306212
rect 371516 306196 371568 306202
rect 371516 306138 371568 306144
rect 371332 306060 371384 306066
rect 371332 306002 371384 306008
rect 370412 305788 370464 305794
rect 370412 305730 370464 305736
rect 370228 305652 370280 305658
rect 370228 305594 370280 305600
rect 370240 157214 370268 305594
rect 370320 302796 370372 302802
rect 370320 302738 370372 302744
rect 370228 157208 370280 157214
rect 370228 157150 370280 157156
rect 370136 156596 370188 156602
rect 370136 156538 370188 156544
rect 370044 155168 370096 155174
rect 370044 155110 370096 155116
rect 370332 155106 370360 302738
rect 370424 158409 370452 305730
rect 370504 303136 370556 303142
rect 370504 303078 370556 303084
rect 370410 158400 370466 158409
rect 370410 158335 370466 158344
rect 370516 157146 370544 303078
rect 370688 303068 370740 303074
rect 370688 303010 370740 303016
rect 370596 302728 370648 302734
rect 370596 302670 370648 302676
rect 370504 157140 370556 157146
rect 370504 157082 370556 157088
rect 370608 156466 370636 302670
rect 370700 158953 370728 303010
rect 371240 285252 371292 285258
rect 371240 285194 371292 285200
rect 370686 158944 370742 158953
rect 370686 158879 370742 158888
rect 370596 156460 370648 156466
rect 370596 156402 370648 156408
rect 370320 155100 370372 155106
rect 370320 155042 370372 155048
rect 369952 9240 370004 9246
rect 369952 9182 370004 9188
rect 368572 8968 368624 8974
rect 368572 8910 368624 8916
rect 368480 6248 368532 6254
rect 368480 6190 368532 6196
rect 368202 3632 368258 3641
rect 368202 3567 368258 3576
rect 369398 3632 369454 3641
rect 369398 3567 369454 3576
rect 370594 3632 370650 3641
rect 370594 3567 370650 3576
rect 365904 3392 365956 3398
rect 365904 3334 365956 3340
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 367020 480 367048 1226
rect 368216 480 368244 3567
rect 369412 480 369440 3567
rect 370608 480 370636 3567
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 285194
rect 371344 155310 371372 306002
rect 371424 305992 371476 305998
rect 371424 305934 371476 305940
rect 371436 155650 371464 305934
rect 371424 155644 371476 155650
rect 371424 155586 371476 155592
rect 371332 155304 371384 155310
rect 371332 155246 371384 155252
rect 371528 155242 371556 306138
rect 371608 305720 371660 305726
rect 371608 305662 371660 305668
rect 371620 157078 371648 305662
rect 371608 157072 371660 157078
rect 371608 157014 371660 157020
rect 371712 156534 371740 306206
rect 371792 303612 371844 303618
rect 371792 303554 371844 303560
rect 371804 156670 371832 303554
rect 373080 303476 373132 303482
rect 373080 303418 373132 303424
rect 372712 303408 372764 303414
rect 372712 303350 372764 303356
rect 371884 302864 371936 302870
rect 371884 302806 371936 302812
rect 371896 159186 371924 302806
rect 372620 298988 372672 298994
rect 372620 298930 372672 298936
rect 371884 159180 371936 159186
rect 371884 159122 371936 159128
rect 371792 156664 371844 156670
rect 371792 156606 371844 156612
rect 371700 156528 371752 156534
rect 371700 156470 371752 156476
rect 371516 155236 371568 155242
rect 371516 155178 371568 155184
rect 372632 16574 372660 298930
rect 372724 154426 372752 303350
rect 372804 303272 372856 303278
rect 372804 303214 372856 303220
rect 372816 154562 372844 303214
rect 372896 303000 372948 303006
rect 372896 302942 372948 302948
rect 372804 154556 372856 154562
rect 372804 154498 372856 154504
rect 372908 154494 372936 302942
rect 372988 302932 373040 302938
rect 372988 302874 373040 302880
rect 373000 155446 373028 302874
rect 373092 158710 373120 303418
rect 373172 303204 373224 303210
rect 373172 303146 373224 303152
rect 373080 158704 373132 158710
rect 373080 158646 373132 158652
rect 373184 158273 373212 303146
rect 375380 300552 375432 300558
rect 375380 300494 375432 300500
rect 374000 286544 374052 286550
rect 374000 286486 374052 286492
rect 373170 158264 373226 158273
rect 373170 158199 373226 158208
rect 372988 155440 373040 155446
rect 372988 155382 373040 155388
rect 372896 154488 372948 154494
rect 372896 154430 372948 154436
rect 372712 154420 372764 154426
rect 372712 154362 372764 154368
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3534 374040 286486
rect 374092 269952 374144 269958
rect 374092 269894 374144 269900
rect 374000 3528 374052 3534
rect 374000 3470 374052 3476
rect 374104 480 374132 269894
rect 375392 16574 375420 300494
rect 376760 269884 376812 269890
rect 376760 269826 376812 269832
rect 376772 16574 376800 269826
rect 375392 16546 376064 16574
rect 376772 16546 377352 16574
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 375300 480 375328 3470
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377324 3482 377352 16546
rect 377416 3602 377444 307226
rect 422300 307216 422352 307222
rect 422300 307158 422352 307164
rect 407118 306096 407174 306105
rect 407118 306031 407174 306040
rect 400220 304496 400272 304502
rect 400220 304438 400272 304444
rect 386418 302968 386474 302977
rect 386418 302903 386474 302912
rect 382280 301708 382332 301714
rect 382280 301650 382332 301656
rect 378140 286476 378192 286482
rect 378140 286418 378192 286424
rect 378152 16574 378180 286418
rect 380900 271380 380952 271386
rect 380900 271322 380952 271328
rect 380912 16574 380940 271322
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 377404 3596 377456 3602
rect 377404 3538 377456 3544
rect 377324 3454 377720 3482
rect 377692 480 377720 3454
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379978 3904 380034 3913
rect 379978 3839 380034 3848
rect 379992 480 380020 3839
rect 381188 480 381216 16546
rect 382292 3466 382320 301650
rect 383660 271312 383712 271318
rect 383660 271254 383712 271260
rect 382372 250572 382424 250578
rect 382372 250514 382424 250520
rect 382280 3460 382332 3466
rect 382280 3402 382332 3408
rect 382384 480 382412 250514
rect 383672 16574 383700 271254
rect 385038 250744 385094 250753
rect 385038 250679 385094 250688
rect 385052 16574 385080 250679
rect 386432 16574 386460 302903
rect 391940 287904 391992 287910
rect 391940 287846 391992 287852
rect 389180 286408 389232 286414
rect 389180 286350 389232 286356
rect 387800 271244 387852 271250
rect 387800 271186 387852 271192
rect 387064 246628 387116 246634
rect 387064 246570 387116 246576
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 383568 3460 383620 3466
rect 383568 3402 383620 3408
rect 383580 480 383608 3402
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387076 3398 387104 246570
rect 387064 3392 387116 3398
rect 387064 3334 387116 3340
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 271186
rect 389192 16574 389220 286350
rect 390560 272672 390612 272678
rect 390560 272614 390612 272620
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3466 390600 272614
rect 391952 16574 391980 287846
rect 396080 287836 396132 287842
rect 396080 287778 396132 287784
rect 394700 272604 394752 272610
rect 394700 272546 394752 272552
rect 394712 16574 394740 272546
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 390650 3496 390706 3505
rect 390560 3460 390612 3466
rect 390650 3431 390706 3440
rect 391848 3460 391900 3466
rect 390560 3402 390612 3408
rect 390664 480 390692 3431
rect 391848 3402 391900 3408
rect 391860 480 391888 3402
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394238 3632 394294 3641
rect 394238 3567 394294 3576
rect 394252 480 394280 3567
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 287778
rect 398840 287768 398892 287774
rect 398840 287710 398892 287716
rect 398852 3534 398880 287710
rect 398932 272536 398984 272542
rect 398932 272478 398984 272484
rect 398840 3528 398892 3534
rect 398840 3470 398892 3476
rect 397734 3360 397790 3369
rect 397734 3295 397790 3304
rect 397748 480 397776 3295
rect 398944 480 398972 272478
rect 400232 16574 400260 304438
rect 404360 304428 404412 304434
rect 404360 304370 404412 304376
rect 402980 289332 403032 289338
rect 402980 289274 403032 289280
rect 401600 274168 401652 274174
rect 401600 274110 401652 274116
rect 401612 16574 401640 274110
rect 402992 16574 403020 289274
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400140 480 400168 3470
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 304370
rect 405740 246492 405792 246498
rect 405740 246434 405792 246440
rect 405752 16574 405780 246434
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3534 407160 306031
rect 418158 305960 418214 305969
rect 418158 305895 418214 305904
rect 415398 302832 415454 302841
rect 415398 302767 415454 302776
rect 414020 290692 414072 290698
rect 414020 290634 414072 290640
rect 407212 289264 407264 289270
rect 407212 289206 407264 289212
rect 407120 3528 407172 3534
rect 407120 3470 407172 3476
rect 407224 480 407252 289206
rect 409880 289196 409932 289202
rect 409880 289138 409932 289144
rect 408500 274100 408552 274106
rect 408500 274042 408552 274048
rect 408512 16574 408540 274042
rect 409892 16574 409920 289138
rect 412640 263084 412692 263090
rect 412640 263026 412692 263032
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 411916 480 411944 3538
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 263026
rect 414032 16574 414060 290634
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3346 415440 302767
rect 416780 287700 416832 287706
rect 416780 287642 416832 287648
rect 415492 274032 415544 274038
rect 415492 273974 415544 273980
rect 415504 3534 415532 273974
rect 416792 16574 416820 287642
rect 418172 16574 418200 305895
rect 420920 289128 420972 289134
rect 420920 289070 420972 289076
rect 419540 275528 419592 275534
rect 419540 275470 419592 275476
rect 419552 16574 419580 275470
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 415412 3318 415532 3346
rect 415504 480 415532 3318
rect 416700 480 416728 3470
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 289070
rect 422312 16574 422340 307158
rect 425060 304360 425112 304366
rect 425060 304302 425112 304308
rect 423680 290624 423732 290630
rect 423680 290566 423732 290572
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3534 423720 290566
rect 423772 273964 423824 273970
rect 423772 273906 423824 273912
rect 423680 3528 423732 3534
rect 423680 3470 423732 3476
rect 423784 480 423812 273906
rect 425072 16574 425100 304302
rect 427820 290556 427872 290562
rect 427820 290498 427872 290504
rect 426440 275460 426492 275466
rect 426440 275402 426492 275408
rect 426452 16574 426480 275402
rect 427832 16574 427860 290498
rect 430580 246424 430632 246430
rect 430580 246366 430632 246372
rect 430592 16574 430620 246366
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 424980 480 425008 3470
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 3460 429712 3466
rect 429660 3402 429712 3408
rect 429672 480 429700 3402
rect 430868 480 430896 16546
rect 431236 3738 431264 308479
rect 471978 308408 472034 308417
rect 471978 308343 472034 308352
rect 442262 305824 442318 305833
rect 442262 305759 442318 305768
rect 440240 301640 440292 301646
rect 440240 301582 440292 301588
rect 431960 292052 432012 292058
rect 431960 291994 432012 292000
rect 431224 3732 431276 3738
rect 431224 3674 431276 3680
rect 431972 3346 432000 291994
rect 438860 290488 438912 290494
rect 438860 290430 438912 290436
rect 437480 276888 437532 276894
rect 437480 276830 437532 276836
rect 433340 275392 433392 275398
rect 433340 275334 433392 275340
rect 432604 263016 432656 263022
rect 432604 262958 432656 262964
rect 432052 254720 432104 254726
rect 432052 254662 432104 254668
rect 432064 3534 432092 254662
rect 432052 3528 432104 3534
rect 432052 3470 432104 3476
rect 432616 3466 432644 262958
rect 433352 16574 433380 275334
rect 436100 264444 436152 264450
rect 436100 264386 436152 264392
rect 434718 250608 434774 250617
rect 434718 250543 434774 250552
rect 434732 16574 434760 250543
rect 436112 16574 436140 264386
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 432604 3460 432656 3466
rect 432604 3402 432656 3408
rect 431972 3318 432092 3346
rect 432064 480 432092 3318
rect 433260 480 433288 3470
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 276830
rect 438872 16574 438900 290430
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3346 440280 301582
rect 440332 269816 440384 269822
rect 440332 269758 440384 269764
rect 440344 3534 440372 269758
rect 441620 249280 441672 249286
rect 441620 249222 441672 249228
rect 441632 16574 441660 249222
rect 441632 16546 442212 16574
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442184 3482 442212 16546
rect 442276 3602 442304 305759
rect 465080 297628 465132 297634
rect 465080 297570 465132 297576
rect 459560 291984 459612 291990
rect 459560 291926 459612 291932
rect 447140 285184 447192 285190
rect 447140 285126 447192 285132
rect 443000 282396 443052 282402
rect 443000 282338 443052 282344
rect 443012 16574 443040 282338
rect 444380 275324 444432 275330
rect 444380 275266 444432 275272
rect 444392 16574 444420 275266
rect 445760 252068 445812 252074
rect 445760 252010 445812 252016
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 442264 3596 442316 3602
rect 442264 3538 442316 3544
rect 440252 3318 440372 3346
rect 440344 480 440372 3318
rect 441540 480 441568 3470
rect 442184 3454 442672 3482
rect 442644 480 442672 3454
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 252010
rect 447152 16574 447180 285126
rect 451280 276820 451332 276826
rect 451280 276762 451332 276768
rect 448520 267232 448572 267238
rect 448520 267174 448572 267180
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3346 448560 267174
rect 449900 265872 449952 265878
rect 449900 265814 449952 265820
rect 448612 252000 448664 252006
rect 448612 251942 448664 251948
rect 448624 3534 448652 251942
rect 449912 16574 449940 265814
rect 451292 16574 451320 276762
rect 455420 276752 455472 276758
rect 455420 276694 455472 276700
rect 454040 256216 454092 256222
rect 454040 256158 454092 256164
rect 452660 251932 452712 251938
rect 452660 251874 452712 251880
rect 452672 16574 452700 251874
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 448532 3318 448652 3346
rect 448624 480 448652 3318
rect 449820 480 449848 3470
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 256158
rect 455432 16574 455460 276694
rect 458180 271176 458232 271182
rect 458180 271118 458232 271124
rect 456800 268592 456852 268598
rect 456800 268534 456852 268540
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3602 456840 268534
rect 457444 264376 457496 264382
rect 457444 264318 457496 264324
rect 456892 251864 456944 251870
rect 456892 251806 456944 251812
rect 456800 3596 456852 3602
rect 456800 3538 456852 3544
rect 456904 480 456932 251806
rect 457456 3670 457484 264318
rect 458192 16574 458220 271118
rect 459572 16574 459600 291926
rect 463700 291916 463752 291922
rect 463700 291858 463752 291864
rect 462320 276684 462372 276690
rect 462320 276626 462372 276632
rect 460940 256148 460992 256154
rect 460940 256090 460992 256096
rect 460952 16574 460980 256090
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 457444 3664 457496 3670
rect 457444 3606 457496 3612
rect 458088 3596 458140 3602
rect 458088 3538 458140 3544
rect 458100 480 458128 3538
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 276626
rect 463712 16574 463740 291858
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 6914 465120 297570
rect 466460 293480 466512 293486
rect 466460 293422 466512 293428
rect 465170 248024 465226 248033
rect 465170 247959 465226 247968
rect 465184 16574 465212 247959
rect 466472 16574 466500 293422
rect 470600 291848 470652 291854
rect 470600 291790 470652 291796
rect 467104 264308 467156 264314
rect 467104 264250 467156 264256
rect 465184 16546 465856 16574
rect 466472 16546 467052 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467024 3482 467052 16546
rect 467116 3670 467144 264250
rect 467840 256080 467892 256086
rect 467840 256022 467892 256028
rect 467852 16574 467880 256022
rect 469218 247888 469274 247897
rect 469218 247823 469274 247832
rect 469232 16574 469260 247823
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 467104 3664 467156 3670
rect 467104 3606 467156 3612
rect 467024 3454 467512 3482
rect 467484 480 467512 3454
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 291790
rect 471992 16574 472020 308343
rect 484400 307148 484452 307154
rect 484400 307090 484452 307096
rect 483018 305688 483074 305697
rect 483018 305623 483074 305632
rect 481640 294840 481692 294846
rect 481640 294782 481692 294788
rect 473360 293412 473412 293418
rect 473360 293354 473412 293360
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3398 473400 293354
rect 477500 293344 477552 293350
rect 477500 293286 477552 293292
rect 476764 264240 476816 264246
rect 476764 264182 476816 264188
rect 474740 256012 474792 256018
rect 474740 255954 474792 255960
rect 473450 247752 473506 247761
rect 473450 247687 473506 247696
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 247687
rect 474752 16574 474780 255954
rect 476120 245132 476172 245138
rect 476120 245074 476172 245080
rect 476132 16574 476160 245074
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 474188 3392 474240 3398
rect 474188 3334 474240 3340
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3334
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 476776 3806 476804 264182
rect 477512 16574 477540 293286
rect 480260 260296 480312 260302
rect 480260 260238 480312 260244
rect 480272 16574 480300 260238
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 476764 3800 476816 3806
rect 476764 3742 476816 3748
rect 478156 480 478184 16546
rect 479340 3732 479392 3738
rect 479340 3674 479392 3680
rect 479352 480 479380 3674
rect 480548 480 480576 16546
rect 481652 3398 481680 294782
rect 481732 246356 481784 246362
rect 481732 246298 481784 246304
rect 481640 3392 481692 3398
rect 481640 3334 481692 3340
rect 481744 480 481772 246298
rect 483032 16574 483060 305623
rect 484412 16574 484440 307090
rect 507860 307080 507912 307086
rect 507860 307022 507912 307028
rect 506480 297560 506532 297566
rect 506480 297502 506532 297508
rect 492680 296200 492732 296206
rect 492680 296142 492732 296148
rect 485780 294772 485832 294778
rect 485780 294714 485832 294720
rect 485792 16574 485820 294714
rect 489920 294704 489972 294710
rect 489920 294646 489972 294652
rect 488540 278248 488592 278254
rect 488540 278190 488592 278196
rect 487160 261724 487212 261730
rect 487160 261666 487212 261672
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 482468 3392 482520 3398
rect 482468 3334 482520 3340
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3334
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 261666
rect 488552 16574 488580 278190
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 480 489960 294646
rect 491300 278180 491352 278186
rect 491300 278122 491352 278128
rect 490012 261656 490064 261662
rect 490012 261598 490064 261604
rect 490024 16574 490052 261598
rect 491312 16574 491340 278122
rect 492692 16574 492720 296142
rect 499580 296132 499632 296138
rect 499580 296074 499632 296080
rect 496820 293276 496872 293282
rect 496820 293218 496872 293224
rect 495440 278112 495492 278118
rect 495440 278054 495492 278060
rect 494060 261588 494112 261594
rect 494060 261530 494112 261536
rect 494072 16574 494100 261530
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 278054
rect 496084 265804 496136 265810
rect 496084 265746 496136 265752
rect 496096 3942 496124 265746
rect 496832 16574 496860 293218
rect 498200 279676 498252 279682
rect 498200 279618 498252 279624
rect 496832 16546 497136 16574
rect 496084 3936 496136 3942
rect 496084 3878 496136 3884
rect 497108 480 497136 16546
rect 498212 3398 498240 279618
rect 498292 262948 498344 262954
rect 498292 262890 498344 262896
rect 498200 3392 498252 3398
rect 498200 3334 498252 3340
rect 498304 3210 498332 262890
rect 499592 16574 499620 296074
rect 503720 296064 503772 296070
rect 503720 296006 503772 296012
rect 502340 279608 502392 279614
rect 502340 279550 502392 279556
rect 499592 16546 500632 16574
rect 499028 3392 499080 3398
rect 499028 3334 499080 3340
rect 498212 3182 498332 3210
rect 498212 480 498240 3182
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3334
rect 500604 480 500632 16546
rect 502352 6914 502380 279550
rect 502984 265736 503036 265742
rect 502984 265678 503036 265684
rect 502996 16574 503024 265678
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 501788 3460 501840 3466
rect 501788 3402 501840 3408
rect 501800 480 501828 3402
rect 502996 480 503024 6886
rect 503088 4010 503116 16546
rect 503076 4004 503128 4010
rect 503076 3946 503128 3952
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 296006
rect 506492 3534 506520 297502
rect 506572 279540 506624 279546
rect 506572 279482 506624 279488
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 505388 480 505416 3470
rect 506584 3346 506612 279482
rect 507872 16574 507900 307022
rect 531320 298920 531372 298926
rect 531320 298862 531372 298868
rect 510620 297492 510672 297498
rect 510620 297434 510672 297440
rect 509240 281036 509292 281042
rect 509240 280978 509292 280984
rect 508504 267164 508556 267170
rect 508504 267106 508556 267112
rect 507872 16546 508452 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 508424 3482 508452 16546
rect 508516 3738 508544 267106
rect 509252 16574 509280 280978
rect 510632 16574 510660 297434
rect 524420 297424 524472 297430
rect 524420 297366 524472 297372
rect 520280 282328 520332 282334
rect 520280 282270 520332 282276
rect 513380 280968 513432 280974
rect 513380 280910 513432 280916
rect 512000 262880 512052 262886
rect 512000 262822 512052 262828
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 508504 3732 508556 3738
rect 508504 3674 508556 3680
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508424 3454 508912 3482
rect 508884 480 508912 3454
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 262822
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 280910
rect 516140 280900 516192 280906
rect 516140 280842 516192 280848
rect 514852 253428 514904 253434
rect 514852 253370 514904 253376
rect 514864 6914 514892 253370
rect 516152 16574 516180 280842
rect 516784 268524 516836 268530
rect 516784 268466 516836 268472
rect 516152 16546 516732 16574
rect 514772 6886 514892 6914
rect 514772 480 514800 6886
rect 515956 3596 516008 3602
rect 515956 3538 516008 3544
rect 515968 480 515996 3538
rect 516704 3482 516732 16546
rect 516796 3874 516824 268466
rect 517520 253360 517572 253366
rect 517520 253302 517572 253308
rect 517532 16574 517560 253302
rect 517532 16546 517928 16574
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 516704 3454 517192 3482
rect 517164 480 517192 3454
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3664 519596 3670
rect 519544 3606 519596 3612
rect 519556 480 519584 3606
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 282270
rect 520924 268456 520976 268462
rect 520924 268398 520976 268404
rect 520936 3466 520964 268398
rect 521660 253292 521712 253298
rect 521660 253234 521712 253240
rect 520924 3460 520976 3466
rect 520924 3402 520976 3408
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 253234
rect 523130 247616 523186 247625
rect 523130 247551 523186 247560
rect 523144 16574 523172 247551
rect 524432 16574 524460 297366
rect 528560 283824 528612 283830
rect 528560 283766 528612 283772
rect 527180 282260 527232 282266
rect 527180 282202 527232 282208
rect 525064 268388 525116 268394
rect 525064 268330 525116 268336
rect 523144 16546 523816 16574
rect 524432 16546 525012 16574
rect 523040 3800 523092 3806
rect 523040 3742 523092 3748
rect 523052 480 523080 3742
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 524984 3482 525012 16546
rect 525076 3602 525104 268330
rect 525800 260228 525852 260234
rect 525800 260170 525852 260176
rect 525812 16574 525840 260170
rect 527192 16574 527220 282202
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524984 3454 525472 3482
rect 525444 480 525472 3454
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 283766
rect 529940 265668 529992 265674
rect 529940 265610 529992 265616
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 265610
rect 531332 3602 531360 298862
rect 535460 298852 535512 298858
rect 535460 298794 535512 298800
rect 531412 282192 531464 282198
rect 531412 282134 531464 282140
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531424 3482 531452 282134
rect 534724 249212 534776 249218
rect 534724 249154 534776 249160
rect 534080 249144 534132 249150
rect 534080 249086 534132 249092
rect 534092 16574 534120 249086
rect 534092 16546 534488 16574
rect 533712 3936 533764 3942
rect 533712 3878 533764 3884
rect 532148 3596 532200 3602
rect 532148 3538 532200 3544
rect 531332 3454 531452 3482
rect 531332 480 531360 3454
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3538
rect 533724 480 533752 3878
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3670 534764 249154
rect 535472 16574 535500 298794
rect 538220 249076 538272 249082
rect 538220 249018 538272 249024
rect 535472 16546 536144 16574
rect 534724 3664 534776 3670
rect 534724 3606 534776 3612
rect 536116 480 536144 16546
rect 537208 4004 537260 4010
rect 537208 3946 537260 3952
rect 537220 480 537248 3946
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 249018
rect 538876 3602 538904 444751
rect 581000 443828 581052 443834
rect 581000 443770 581052 443776
rect 580632 443760 580684 443766
rect 580632 443702 580684 443708
rect 580540 443692 580592 443698
rect 580540 443634 580592 443640
rect 580356 443284 580408 443290
rect 580356 443226 580408 443232
rect 580264 443216 580316 443222
rect 580264 443158 580316 443164
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 579620 379500 579672 379506
rect 579620 379442 579672 379448
rect 579632 378457 579660 379442
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 560300 301572 560352 301578
rect 560300 301514 560352 301520
rect 542360 300280 542412 300286
rect 542360 300222 542412 300228
rect 539600 298784 539652 298790
rect 539600 298726 539652 298732
rect 538956 283756 539008 283762
rect 538956 283698 539008 283704
rect 538968 3806 538996 283698
rect 538956 3800 539008 3806
rect 538956 3742 539008 3748
rect 538864 3596 538916 3602
rect 538864 3538 538916 3544
rect 539612 480 539640 298726
rect 539692 261520 539744 261526
rect 539692 261462 539744 261468
rect 539704 16574 539732 261462
rect 542372 16574 542400 300222
rect 553400 300212 553452 300218
rect 553400 300154 553452 300160
rect 549260 294636 549312 294642
rect 549260 294578 549312 294584
rect 547880 283688 547932 283694
rect 547880 283630 547932 283636
rect 545120 278044 545172 278050
rect 545120 277986 545172 277992
rect 543740 267096 543792 267102
rect 543740 267038 543792 267044
rect 543752 16574 543780 267038
rect 545132 16574 545160 277986
rect 546498 250472 546554 250481
rect 546498 250407 546554 250416
rect 539704 16546 540376 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 3664 542044 3670
rect 541992 3606 542044 3612
rect 542004 480 542032 3606
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 250407
rect 547892 3398 547920 283630
rect 547972 267028 548024 267034
rect 547972 266970 548024 266976
rect 547880 3392 547932 3398
rect 547880 3334 547932 3340
rect 547984 3210 548012 266970
rect 549272 16574 549300 294578
rect 552664 285116 552716 285122
rect 552664 285058 552716 285064
rect 552020 283620 552072 283626
rect 552020 283562 552072 283568
rect 549272 16546 550312 16574
rect 548708 3392 548760 3398
rect 548708 3334 548760 3340
rect 547892 3182 548012 3210
rect 547892 480 547920 3182
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3334
rect 550284 480 550312 16546
rect 552032 6914 552060 283562
rect 552676 16574 552704 285058
rect 553412 16574 553440 300154
rect 556160 300144 556212 300150
rect 556160 300086 556212 300092
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 551468 3732 551520 3738
rect 551468 3674 551520 3680
rect 551480 480 551508 3674
rect 552676 480 552704 6886
rect 552768 3670 552796 16546
rect 552756 3664 552808 3670
rect 552756 3606 552808 3612
rect 553780 480 553808 16546
rect 554964 3868 555016 3874
rect 554964 3810 555016 3816
rect 554976 480 555004 3810
rect 556172 3398 556200 300086
rect 556252 279472 556304 279478
rect 556252 279414 556304 279420
rect 556160 3392 556212 3398
rect 556160 3334 556212 3340
rect 556264 3210 556292 279414
rect 557540 245064 557592 245070
rect 557540 245006 557592 245012
rect 557552 16574 557580 245006
rect 560312 16574 560340 301514
rect 564440 301504 564492 301510
rect 564440 301446 564492 301452
rect 563060 280832 563112 280838
rect 563060 280774 563112 280780
rect 561680 244996 561732 245002
rect 561680 244938 561732 244944
rect 561692 16574 561720 244938
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556988 3392 557040 3398
rect 556988 3334 557040 3340
rect 556172 3182 556292 3210
rect 556172 480 556200 3182
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557000 354 557028 3334
rect 558564 480 558592 16546
rect 559748 3800 559800 3806
rect 559748 3742 559800 3748
rect 559760 480 559788 3742
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 280774
rect 564452 480 564480 301446
rect 567200 295996 567252 296002
rect 567200 295938 567252 295944
rect 565820 285048 565872 285054
rect 565820 284990 565872 284996
rect 564532 244928 564584 244934
rect 564532 244870 564584 244876
rect 564544 16574 564572 244870
rect 565832 16574 565860 284990
rect 567212 16574 567240 295938
rect 576860 286340 576912 286346
rect 576860 286282 576912 286288
rect 569960 284980 570012 284986
rect 569960 284922 570012 284928
rect 569972 16574 570000 284922
rect 575480 260160 575532 260166
rect 575480 260102 575532 260108
rect 574100 254652 574152 254658
rect 574100 254594 574152 254600
rect 571340 253224 571392 253230
rect 571340 253166 571392 253172
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 3460 569184 3466
rect 569132 3402 569184 3408
rect 569144 480 569172 3402
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 253166
rect 574112 16574 574140 254594
rect 575492 16574 575520 260102
rect 576872 16574 576900 286282
rect 579620 273216 579672 273222
rect 579620 273158 579672 273164
rect 579632 272241 579660 273158
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 578240 254584 578292 254590
rect 578240 254526 578292 254532
rect 578252 16574 578280 254526
rect 580276 33153 580304 443158
rect 580368 112849 580396 443226
rect 580448 441652 580500 441658
rect 580448 441594 580500 441600
rect 580460 152697 580488 441594
rect 580552 232393 580580 443634
rect 580644 325281 580672 443702
rect 580630 325272 580686 325281
rect 580630 325207 580686 325216
rect 580538 232384 580594 232393
rect 580538 232319 580594 232328
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580354 112840 580410 112849
rect 580354 112775 580410 112784
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 573916 3664 573968 3670
rect 573916 3606 573968 3612
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572732 480 572760 3470
rect 573928 480 573956 3606
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 581012 480 581040 443770
rect 582194 4856 582250 4865
rect 582194 4791 582250 4800
rect 582208 480 582236 4791
rect 583392 3596 583444 3602
rect 583392 3538 583444 3544
rect 583404 480 583432 3538
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3422 671200 3478 671256
rect 2778 658144 2834 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3238 566888 3294 566944
rect 2778 553832 2834 553888
rect 2962 527856 3018 527912
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3146 449520 3202 449576
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 579944 3570 580000
rect 3514 514800 3570 514856
rect 3606 501744 3662 501800
rect 217874 516840 217930 516896
rect 217782 515888 217838 515944
rect 217690 513712 217746 513768
rect 217598 489912 217654 489968
rect 217322 488280 217378 488336
rect 217506 488008 217562 488064
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 2870 397432 2926 397488
rect 2870 371320 2926 371376
rect 3330 358400 3386 358456
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 267144 3386 267200
rect 2870 254088 2926 254144
rect 3146 110608 3202 110664
rect 3974 345344 4030 345400
rect 3882 293120 3938 293176
rect 3790 241032 3846 241088
rect 3698 201864 3754 201920
rect 3606 188808 3662 188864
rect 3606 149776 3662 149832
rect 3514 136720 3570 136776
rect 3514 97588 3516 97608
rect 3516 97588 3568 97608
rect 3568 97588 3570 97608
rect 3514 97552 3570 97588
rect 3422 84632 3478 84688
rect 75182 308352 75238 308408
rect 219070 512760 219126 512816
rect 219346 510992 219402 511048
rect 219254 509904 219310 509960
rect 219162 508136 219218 508192
rect 247038 476584 247094 476640
rect 210882 303320 210938 303376
rect 211894 303184 211950 303240
rect 210974 300056 211030 300112
rect 210974 155216 211030 155272
rect 208582 3304 208638 3360
rect 212078 302912 212134 302968
rect 212262 302776 212318 302832
rect 213366 155760 213422 155816
rect 213274 155488 213330 155544
rect 213366 3440 213422 3496
rect 214746 300192 214802 300248
rect 214654 158616 214710 158672
rect 214470 3440 214526 3496
rect 214930 3984 214986 4040
rect 215022 3848 215078 3904
rect 215114 3712 215170 3768
rect 216218 158072 216274 158128
rect 216034 155624 216090 155680
rect 215666 3440 215722 3496
rect 214838 3168 214894 3224
rect 217046 193704 217102 193760
rect 216678 192752 216734 192808
rect 216678 188128 216734 188184
rect 217506 196832 217562 196888
rect 217414 195880 217470 195936
rect 217230 169904 217286 169960
rect 216862 3576 216918 3632
rect 216586 3304 216642 3360
rect 217690 168272 217746 168328
rect 217598 168000 217654 168056
rect 218794 300328 218850 300384
rect 218426 243480 218482 243536
rect 218518 190984 218574 191040
rect 217966 155896 218022 155952
rect 217782 155352 217838 155408
rect 218702 189896 218758 189952
rect 218978 158636 219034 158672
rect 218978 158616 218980 158636
rect 218980 158616 219032 158636
rect 219032 158616 219034 158636
rect 235906 476176 235962 476232
rect 237470 476312 237526 476368
rect 237562 476176 237618 476232
rect 240138 476176 240194 476232
rect 241426 476176 241482 476232
rect 244278 476468 244334 476504
rect 244278 476448 244280 476468
rect 244280 476448 244332 476468
rect 244332 476448 244334 476468
rect 242898 476332 242954 476368
rect 242898 476312 242900 476332
rect 242900 476312 242952 476332
rect 242952 476312 242954 476332
rect 244278 476312 244334 476368
rect 242806 476196 242862 476232
rect 242806 476176 242808 476196
rect 242808 476176 242860 476196
rect 242860 476176 242862 476196
rect 245658 476176 245714 476232
rect 247222 476176 247278 476232
rect 249798 476584 249854 476640
rect 249798 476176 249854 476232
rect 251086 476196 251142 476232
rect 251086 476176 251088 476196
rect 251088 476176 251140 476196
rect 251140 476176 251142 476196
rect 277766 476992 277822 477048
rect 304998 476992 305054 477048
rect 307758 476992 307814 477048
rect 253846 476856 253902 476912
rect 256606 476856 256662 476912
rect 270498 476856 270554 476912
rect 252558 476604 252614 476640
rect 252558 476584 252560 476604
rect 252560 476584 252612 476604
rect 252612 476584 252614 476604
rect 252374 476312 252430 476368
rect 255410 476720 255466 476776
rect 252466 476176 252522 476232
rect 257986 476312 258042 476368
rect 255962 476176 256018 476232
rect 258262 476332 258318 476368
rect 258262 476312 258264 476332
rect 258264 476312 258316 476332
rect 258316 476312 258318 476332
rect 258170 476196 258226 476232
rect 258170 476176 258172 476196
rect 258172 476176 258224 476196
rect 258224 476176 258226 476196
rect 263598 476604 263654 476640
rect 263598 476584 263600 476604
rect 263600 476584 263652 476604
rect 263652 476584 263654 476604
rect 264978 476584 265034 476640
rect 260746 476448 260802 476504
rect 267830 476468 267886 476504
rect 267830 476448 267832 476468
rect 267832 476448 267884 476468
rect 267884 476448 267886 476468
rect 273166 476584 273222 476640
rect 260838 476312 260894 476368
rect 260746 476176 260802 476232
rect 267646 476312 267702 476368
rect 262126 476176 262182 476232
rect 263506 476176 263562 476232
rect 264886 476176 264942 476232
rect 266266 476176 266322 476232
rect 267554 476176 267610 476232
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476176 271842 476232
rect 273258 476448 273314 476504
rect 274546 476312 274602 476368
rect 276018 476312 276074 476368
rect 274454 476176 274510 476232
rect 275926 476176 275982 476232
rect 302238 476740 302294 476776
rect 302238 476720 302240 476740
rect 302240 476720 302292 476740
rect 302292 476720 302294 476740
rect 277306 476176 277362 476232
rect 278686 476176 278742 476232
rect 280158 476312 280214 476368
rect 280066 476176 280122 476232
rect 283010 476176 283066 476232
rect 310518 476856 310574 476912
rect 285862 476176 285918 476232
rect 287242 476176 287298 476232
rect 289818 476176 289874 476232
rect 292670 476176 292726 476232
rect 295338 476176 295394 476232
rect 298098 476176 298154 476232
rect 300858 476176 300914 476232
rect 295982 444760 296038 444816
rect 294418 444624 294474 444680
rect 295154 444488 295210 444544
rect 299754 443264 299810 443320
rect 322938 476856 322994 476912
rect 313278 476468 313334 476504
rect 313278 476448 313280 476468
rect 313280 476448 313332 476468
rect 313332 476448 313334 476468
rect 314658 476448 314714 476504
rect 317418 476332 317474 476368
rect 317418 476312 317420 476332
rect 317420 476312 317472 476332
rect 317472 476312 317474 476332
rect 320178 476312 320234 476368
rect 325790 476176 325846 476232
rect 342258 444624 342314 444680
rect 345294 443128 345350 443184
rect 347594 442992 347650 443048
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 617480 580226 617536
rect 579802 564304 579858 564360
rect 579618 537784 579674 537840
rect 580170 484608 580226 484664
rect 580354 630808 580410 630864
rect 580446 590960 580502 591016
rect 580538 577632 580594 577688
rect 538862 444760 538918 444816
rect 307022 442176 307078 442232
rect 361210 442176 361266 442232
rect 361946 442176 362002 442232
rect 218794 3984 218850 4040
rect 218794 3576 218850 3632
rect 218058 3440 218114 3496
rect 233238 308352 233294 308408
rect 272154 273808 272210 273864
rect 275190 308896 275246 308952
rect 275006 306040 275062 306096
rect 275926 308624 275982 308680
rect 275650 306176 275706 306232
rect 276570 308760 276626 308816
rect 274730 303320 274786 303376
rect 277214 308488 277270 308544
rect 277490 305904 277546 305960
rect 277030 303184 277086 303240
rect 278410 303048 278466 303104
rect 277674 302912 277730 302968
rect 279054 302776 279110 302832
rect 280894 305768 280950 305824
rect 280710 305632 280766 305688
rect 283286 300328 283342 300384
rect 283102 300192 283158 300248
rect 284574 300056 284630 300112
rect 273626 275168 273682 275224
rect 273534 267008 273590 267064
rect 273442 262792 273498 262848
rect 273350 249056 273406 249112
rect 294418 308624 294474 308680
rect 295338 244976 295394 245032
rect 296718 245384 296774 245440
rect 298466 308760 298522 308816
rect 299570 248104 299626 248160
rect 299478 245520 299534 245576
rect 298098 245248 298154 245304
rect 296902 245112 296958 245168
rect 295522 244840 295578 244896
rect 299846 250824 299902 250880
rect 301318 264152 301374 264208
rect 302330 265512 302386 265568
rect 302238 254632 302294 254688
rect 302698 283464 302754 283520
rect 302606 282104 302662 282160
rect 303986 297336 304042 297392
rect 303710 269728 303766 269784
rect 302422 254496 302478 254552
rect 305642 301416 305698 301472
rect 307206 302912 307262 302968
rect 307850 303184 307906 303240
rect 308586 303048 308642 303104
rect 309782 304136 309838 304192
rect 306378 250688 306434 250744
rect 311346 306040 311402 306096
rect 312634 302776 312690 302832
rect 313646 305904 313702 305960
rect 316038 250552 316094 250608
rect 321558 247968 321614 248024
rect 323674 308352 323730 308408
rect 323122 247832 323178 247888
rect 322938 247696 322994 247752
rect 301042 246200 301098 246256
rect 325054 308488 325110 308544
rect 326066 305632 326122 305688
rect 330206 305768 330262 305824
rect 336830 250416 336886 250472
rect 332598 247560 332654 247616
rect 345110 309032 345166 309088
rect 346030 308896 346086 308952
rect 348146 306176 348202 306232
rect 299662 244704 299718 244760
rect 356334 245248 356390 245304
rect 356610 245112 356666 245168
rect 356334 244568 356390 244624
rect 356610 244432 356666 244488
rect 355506 243888 355562 243944
rect 277030 159840 277086 159896
rect 278134 159840 278190 159896
rect 279238 159840 279294 159896
rect 285954 159840 286010 159896
rect 256054 159568 256110 159624
rect 227718 158616 227774 158672
rect 238114 158652 238116 158672
rect 238116 158652 238168 158672
rect 238168 158652 238170 158672
rect 224314 158208 224370 158264
rect 224958 157800 225014 157856
rect 224314 157664 224370 157720
rect 219346 3440 219402 3496
rect 219346 3168 219402 3224
rect 222750 3848 222806 3904
rect 238114 158616 238170 158652
rect 239586 158616 239642 158672
rect 242438 158616 242494 158672
rect 244278 158616 244334 158672
rect 248326 158616 248382 158672
rect 250902 158616 250958 158672
rect 252098 158616 252154 158672
rect 231858 158480 231914 158536
rect 227534 3712 227590 3768
rect 226338 3576 226394 3632
rect 233238 158344 233294 158400
rect 237378 158208 237434 158264
rect 240598 158344 240654 158400
rect 237010 3440 237066 3496
rect 240506 3304 240562 3360
rect 245566 157800 245622 157856
rect 246762 158072 246818 158128
rect 247774 157800 247830 157856
rect 249798 158208 249854 158264
rect 248694 157800 248750 157856
rect 250718 157800 250774 157856
rect 251178 157936 251234 157992
rect 253478 157800 253534 157856
rect 271050 159568 271106 159624
rect 275834 159568 275890 159624
rect 257342 158616 257398 158672
rect 259918 158616 259974 158672
rect 261758 158616 261814 158672
rect 264334 158616 264390 158672
rect 265898 158616 265954 158672
rect 268382 158652 268384 158672
rect 268384 158652 268436 158672
rect 268436 158652 268438 158672
rect 268382 158616 268438 158652
rect 268750 158636 268806 158672
rect 268750 158616 268752 158636
rect 268752 158616 268804 158636
rect 268804 158616 268806 158636
rect 261206 157528 261262 157584
rect 260838 155760 260894 155816
rect 263690 157528 263746 157584
rect 263598 155624 263654 155680
rect 269854 158616 269910 158672
rect 266634 157664 266690 157720
rect 265990 157528 266046 157584
rect 264978 155896 265034 155952
rect 271142 158616 271198 158672
rect 272246 158616 272302 158672
rect 273350 158616 273406 158672
rect 274454 158616 274510 158672
rect 276110 158616 276166 158672
rect 281078 158616 281134 158672
rect 273718 157664 273774 157720
rect 267738 155488 267794 155544
rect 278502 157664 278558 157720
rect 274638 155352 274694 155408
rect 267830 155216 267886 155272
rect 283654 158616 283710 158672
rect 291014 159568 291070 159624
rect 293590 158616 293646 158672
rect 295982 158616 296038 158672
rect 298558 158616 298614 158672
rect 301042 158616 301098 158672
rect 303526 158616 303582 158672
rect 306102 158616 306158 158672
rect 288254 157528 288310 157584
rect 308678 158616 308734 158672
rect 311070 158616 311126 158672
rect 313462 158616 313518 158672
rect 315854 158616 315910 158672
rect 318614 158616 318670 158672
rect 321006 158616 321062 158672
rect 323398 158616 323454 158672
rect 325974 158616 326030 158672
rect 355506 157800 355562 157856
rect 319718 8880 319774 8936
rect 350446 6704 350502 6760
rect 348054 6568 348110 6624
rect 344558 6432 344614 6488
rect 340970 6296 341026 6352
rect 337474 6160 337530 6216
rect 327998 3304 328054 3360
rect 331586 3440 331642 3496
rect 335082 3576 335138 3632
rect 338670 3712 338726 3768
rect 345754 3984 345810 4040
rect 349250 3168 349306 3224
rect 351642 3848 351698 3904
rect 356242 3712 356298 3768
rect 356886 245520 356942 245576
rect 357438 245556 357440 245576
rect 357440 245556 357492 245576
rect 357492 245556 357494 245576
rect 357438 245520 357494 245556
rect 356886 245112 356942 245168
rect 357438 158752 357494 158808
rect 356242 3168 356298 3224
rect 358174 245384 358230 245440
rect 358634 306312 358690 306368
rect 360106 306312 360162 306368
rect 358726 3576 358782 3632
rect 357530 3440 357586 3496
rect 359922 3440 359978 3496
rect 361118 3440 361174 3496
rect 362406 308760 362462 308816
rect 363694 309032 363750 309088
rect 362314 3440 362370 3496
rect 363418 243888 363474 243944
rect 363326 6704 363382 6760
rect 363786 308896 363842 308952
rect 365810 308624 365866 308680
rect 363786 158480 363842 158536
rect 363694 157392 363750 157448
rect 363234 6160 363290 6216
rect 364706 6296 364762 6352
rect 365258 159568 365314 159624
rect 364614 3576 364670 3632
rect 363510 3440 363566 3496
rect 365810 3576 365866 3632
rect 366362 159160 366418 159216
rect 366454 159024 366510 159080
rect 366546 158752 366602 158808
rect 366270 158072 366326 158128
rect 365994 8880 366050 8936
rect 367834 159296 367890 159352
rect 367190 6568 367246 6624
rect 367098 6432 367154 6488
rect 369030 306176 369086 306232
rect 431222 308488 431278 308544
rect 369214 157936 369270 157992
rect 370410 158344 370466 158400
rect 370686 158888 370742 158944
rect 368202 3576 368258 3632
rect 369398 3576 369454 3632
rect 370594 3576 370650 3632
rect 373170 158208 373226 158264
rect 407118 306040 407174 306096
rect 386418 302912 386474 302968
rect 379978 3848 380034 3904
rect 385038 250688 385094 250744
rect 390650 3440 390706 3496
rect 394238 3576 394294 3632
rect 397734 3304 397790 3360
rect 418158 305904 418214 305960
rect 415398 302776 415454 302832
rect 471978 308352 472034 308408
rect 442262 305768 442318 305824
rect 434718 250552 434774 250608
rect 465170 247968 465226 248024
rect 469218 247832 469274 247888
rect 483018 305632 483074 305688
rect 473450 247696 473506 247752
rect 523130 247560 523186 247616
rect 580170 431568 580226 431624
rect 579618 378392 579674 378448
rect 546498 250416 546554 250472
rect 579618 272176 579674 272232
rect 580630 325216 580686 325272
rect 580538 232328 580594 232384
rect 580446 152632 580502 152688
rect 580354 112784 580410 112840
rect 580262 33088 580318 33144
rect 582194 4800 582250 4856
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 580533 577690 580599 577693
rect 583520 577690 584960 577780
rect 580533 577688 584960 577690
rect 580533 577632 580538 577688
rect 580594 577632 584960 577688
rect 580533 577630 584960 577632
rect 580533 577627 580599 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579613 537842 579679 537845
rect 583520 537842 584960 537932
rect 579613 537840 584960 537842
rect 579613 537784 579618 537840
rect 579674 537784 584960 537840
rect 579613 537782 584960 537784
rect 579613 537779 579679 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 583520 524364 584960 524604
rect 217869 516898 217935 516901
rect 219390 516898 220064 516924
rect 217869 516896 220064 516898
rect 217869 516840 217874 516896
rect 217930 516864 220064 516896
rect 217930 516840 219450 516864
rect 217869 516838 219450 516840
rect 217869 516835 217935 516838
rect 217777 515946 217843 515949
rect 219390 515946 220064 515972
rect 217777 515944 220064 515946
rect 217777 515888 217782 515944
rect 217838 515912 220064 515944
rect 217838 515888 219450 515912
rect 217777 515886 219450 515888
rect 217777 515883 217843 515886
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 217685 513770 217751 513773
rect 219390 513770 220064 513796
rect 217685 513768 220064 513770
rect 217685 513712 217690 513768
rect 217746 513736 220064 513768
rect 217746 513712 219450 513736
rect 217685 513710 219450 513712
rect 217685 513707 217751 513710
rect 219065 512818 219131 512821
rect 219390 512818 220064 512844
rect 219065 512816 220064 512818
rect 219065 512760 219070 512816
rect 219126 512784 220064 512816
rect 219126 512760 219450 512784
rect 219065 512758 219450 512760
rect 219065 512755 219131 512758
rect 583520 511172 584960 511412
rect 219390 511053 220064 511076
rect 219341 511048 220064 511053
rect 219341 510992 219346 511048
rect 219402 511016 220064 511048
rect 219402 510992 219450 511016
rect 219341 510990 219450 510992
rect 219341 510987 219407 510990
rect 219249 509962 219315 509965
rect 219390 509962 220064 509988
rect 219249 509960 220064 509962
rect 219249 509904 219254 509960
rect 219310 509928 220064 509960
rect 219310 509904 219450 509928
rect 219249 509902 219450 509904
rect 219249 509899 219315 509902
rect 219157 508194 219223 508197
rect 219390 508194 220064 508220
rect 219157 508192 220064 508194
rect 219157 508136 219162 508192
rect 219218 508160 220064 508192
rect 219218 508136 219450 508160
rect 219157 508134 219450 508136
rect 219157 508131 219223 508134
rect -960 501802 480 501892
rect 3601 501802 3667 501805
rect -960 501800 3667 501802
rect -960 501744 3606 501800
rect 3662 501744 3667 501800
rect -960 501742 3667 501744
rect -960 501652 480 501742
rect 3601 501739 3667 501742
rect 583520 497844 584960 498084
rect 217593 489970 217659 489973
rect 219390 489970 220064 489996
rect 217593 489968 220064 489970
rect 217593 489912 217598 489968
rect 217654 489936 220064 489968
rect 217654 489912 219450 489936
rect 217593 489910 219450 489912
rect 217593 489907 217659 489910
rect -960 488596 480 488836
rect 217317 488338 217383 488341
rect 219390 488338 220064 488364
rect 217317 488336 220064 488338
rect 217317 488280 217322 488336
rect 217378 488304 220064 488336
rect 217378 488280 219450 488304
rect 217317 488278 219450 488280
rect 217317 488275 217383 488278
rect 217501 488066 217567 488069
rect 219390 488066 220064 488092
rect 217501 488064 220064 488066
rect 217501 488008 217506 488064
rect 217562 488032 220064 488064
rect 217562 488008 219450 488032
rect 217501 488006 219450 488008
rect 217501 488003 217567 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 277761 477050 277827 477053
rect 278446 477050 278452 477052
rect 277761 477048 278452 477050
rect 277761 476992 277766 477048
rect 277822 476992 278452 477048
rect 277761 476990 278452 476992
rect 277761 476987 277827 476990
rect 278446 476988 278452 476990
rect 278516 476988 278522 477052
rect 304993 477050 305059 477053
rect 305862 477050 305868 477052
rect 304993 477048 305868 477050
rect 304993 476992 304998 477048
rect 305054 476992 305868 477048
rect 304993 476990 305868 476992
rect 304993 476987 305059 476990
rect 305862 476988 305868 476990
rect 305932 476988 305938 477052
rect 307753 477050 307819 477053
rect 308438 477050 308444 477052
rect 307753 477048 308444 477050
rect 307753 476992 307758 477048
rect 307814 476992 308444 477048
rect 307753 476990 308444 476992
rect 307753 476987 307819 476990
rect 308438 476988 308444 476990
rect 308508 476988 308514 477052
rect 253422 476852 253428 476916
rect 253492 476914 253498 476916
rect 253841 476914 253907 476917
rect 253492 476912 253907 476914
rect 253492 476856 253846 476912
rect 253902 476856 253907 476912
rect 253492 476854 253907 476856
rect 253492 476852 253498 476854
rect 253841 476851 253907 476854
rect 255814 476852 255820 476916
rect 255884 476914 255890 476916
rect 256601 476914 256667 476917
rect 255884 476912 256667 476914
rect 255884 476856 256606 476912
rect 256662 476856 256667 476912
rect 255884 476854 256667 476856
rect 255884 476852 255890 476854
rect 256601 476851 256667 476854
rect 270493 476914 270559 476917
rect 270902 476914 270908 476916
rect 270493 476912 270908 476914
rect 270493 476856 270498 476912
rect 270554 476856 270908 476912
rect 270493 476854 270908 476856
rect 270493 476851 270559 476854
rect 270902 476852 270908 476854
rect 270972 476852 270978 476916
rect 310513 476914 310579 476917
rect 311014 476914 311020 476916
rect 310513 476912 311020 476914
rect 310513 476856 310518 476912
rect 310574 476856 311020 476912
rect 310513 476854 311020 476856
rect 310513 476851 310579 476854
rect 311014 476852 311020 476854
rect 311084 476852 311090 476916
rect 322933 476914 322999 476917
rect 323342 476914 323348 476916
rect 322933 476912 323348 476914
rect 322933 476856 322938 476912
rect 322994 476856 323348 476912
rect 322933 476854 323348 476856
rect 322933 476851 322999 476854
rect 323342 476852 323348 476854
rect 323412 476852 323418 476916
rect 255405 476778 255471 476781
rect 256182 476778 256188 476780
rect 255405 476776 256188 476778
rect 255405 476720 255410 476776
rect 255466 476720 256188 476776
rect 255405 476718 256188 476720
rect 255405 476715 255471 476718
rect 256182 476716 256188 476718
rect 256252 476716 256258 476780
rect 302233 476778 302299 476781
rect 303470 476778 303476 476780
rect 302233 476776 303476 476778
rect 302233 476720 302238 476776
rect 302294 476720 303476 476776
rect 302233 476718 303476 476720
rect 302233 476715 302299 476718
rect 303470 476716 303476 476718
rect 303540 476716 303546 476780
rect 247033 476642 247099 476645
rect 248270 476642 248276 476644
rect 247033 476640 248276 476642
rect 247033 476584 247038 476640
rect 247094 476584 248276 476640
rect 247033 476582 248276 476584
rect 247033 476579 247099 476582
rect 248270 476580 248276 476582
rect 248340 476580 248346 476644
rect 249793 476642 249859 476645
rect 250662 476642 250668 476644
rect 249793 476640 250668 476642
rect 249793 476584 249798 476640
rect 249854 476584 250668 476640
rect 249793 476582 250668 476584
rect 249793 476579 249859 476582
rect 250662 476580 250668 476582
rect 250732 476580 250738 476644
rect 252553 476642 252619 476645
rect 263593 476644 263659 476645
rect 253606 476642 253612 476644
rect 252553 476640 253612 476642
rect 252553 476584 252558 476640
rect 252614 476584 253612 476640
rect 252553 476582 253612 476584
rect 252553 476579 252619 476582
rect 253606 476580 253612 476582
rect 253676 476580 253682 476644
rect 263542 476580 263548 476644
rect 263612 476642 263659 476644
rect 264973 476642 265039 476645
rect 265934 476642 265940 476644
rect 263612 476640 263704 476642
rect 263654 476584 263704 476640
rect 263612 476582 263704 476584
rect 264973 476640 265940 476642
rect 264973 476584 264978 476640
rect 265034 476584 265940 476640
rect 264973 476582 265940 476584
rect 263612 476580 263659 476582
rect 263593 476579 263659 476580
rect 264973 476579 265039 476582
rect 265934 476580 265940 476582
rect 266004 476580 266010 476644
rect 272190 476580 272196 476644
rect 272260 476642 272266 476644
rect 273161 476642 273227 476645
rect 272260 476640 273227 476642
rect 272260 476584 273166 476640
rect 273222 476584 273227 476640
rect 272260 476582 273227 476584
rect 272260 476580 272266 476582
rect 273161 476579 273227 476582
rect 244273 476508 244339 476509
rect 244222 476444 244228 476508
rect 244292 476506 244339 476508
rect 244292 476504 244384 476506
rect 244334 476448 244384 476504
rect 244292 476446 244384 476448
rect 244292 476444 244339 476446
rect 260598 476444 260604 476508
rect 260668 476506 260674 476508
rect 260741 476506 260807 476509
rect 260668 476504 260807 476506
rect 260668 476448 260746 476504
rect 260802 476448 260807 476504
rect 260668 476446 260807 476448
rect 260668 476444 260674 476446
rect 244273 476443 244339 476444
rect 260741 476443 260807 476446
rect 267825 476506 267891 476509
rect 268326 476506 268332 476508
rect 267825 476504 268332 476506
rect 267825 476448 267830 476504
rect 267886 476448 268332 476504
rect 267825 476446 268332 476448
rect 267825 476443 267891 476446
rect 268326 476444 268332 476446
rect 268396 476444 268402 476508
rect 273253 476506 273319 476509
rect 273478 476506 273484 476508
rect 273253 476504 273484 476506
rect 273253 476448 273258 476504
rect 273314 476448 273484 476504
rect 273253 476446 273484 476448
rect 273253 476443 273319 476446
rect 273478 476444 273484 476446
rect 273548 476444 273554 476508
rect 313273 476506 313339 476509
rect 313406 476506 313412 476508
rect 313273 476504 313412 476506
rect 313273 476448 313278 476504
rect 313334 476448 313412 476504
rect 313273 476446 313412 476448
rect 313273 476443 313339 476446
rect 313406 476444 313412 476446
rect 313476 476444 313482 476508
rect 314653 476506 314719 476509
rect 315798 476506 315804 476508
rect 314653 476504 315804 476506
rect 314653 476448 314658 476504
rect 314714 476448 315804 476504
rect 314653 476446 315804 476448
rect 314653 476443 314719 476446
rect 315798 476444 315804 476446
rect 315868 476444 315874 476508
rect 237465 476370 237531 476373
rect 238150 476370 238156 476372
rect 237465 476368 238156 476370
rect 237465 476312 237470 476368
rect 237526 476312 238156 476368
rect 237465 476310 238156 476312
rect 237465 476307 237531 476310
rect 238150 476308 238156 476310
rect 238220 476308 238226 476372
rect 242893 476370 242959 476373
rect 243118 476370 243124 476372
rect 242893 476368 243124 476370
rect 242893 476312 242898 476368
rect 242954 476312 243124 476368
rect 242893 476310 243124 476312
rect 242893 476307 242959 476310
rect 243118 476308 243124 476310
rect 243188 476308 243194 476372
rect 244273 476370 244339 476373
rect 245326 476370 245332 476372
rect 244273 476368 245332 476370
rect 244273 476312 244278 476368
rect 244334 476312 245332 476368
rect 244273 476310 245332 476312
rect 244273 476307 244339 476310
rect 245326 476308 245332 476310
rect 245396 476308 245402 476372
rect 251398 476308 251404 476372
rect 251468 476370 251474 476372
rect 252369 476370 252435 476373
rect 251468 476368 252435 476370
rect 251468 476312 252374 476368
rect 252430 476312 252435 476368
rect 251468 476310 252435 476312
rect 251468 476308 251474 476310
rect 252369 476307 252435 476310
rect 257102 476308 257108 476372
rect 257172 476370 257178 476372
rect 257981 476370 258047 476373
rect 257172 476368 258047 476370
rect 257172 476312 257986 476368
rect 258042 476312 258047 476368
rect 257172 476310 258047 476312
rect 257172 476308 257178 476310
rect 257981 476307 258047 476310
rect 258257 476370 258323 476373
rect 258390 476370 258396 476372
rect 258257 476368 258396 476370
rect 258257 476312 258262 476368
rect 258318 476312 258396 476368
rect 258257 476310 258396 476312
rect 258257 476307 258323 476310
rect 258390 476308 258396 476310
rect 258460 476308 258466 476372
rect 260833 476370 260899 476373
rect 260966 476370 260972 476372
rect 260833 476368 260972 476370
rect 260833 476312 260838 476368
rect 260894 476312 260972 476368
rect 260833 476310 260972 476312
rect 260833 476307 260899 476310
rect 260966 476308 260972 476310
rect 261036 476308 261042 476372
rect 266486 476308 266492 476372
rect 266556 476370 266562 476372
rect 267641 476370 267707 476373
rect 266556 476368 267707 476370
rect 266556 476312 267646 476368
rect 267702 476312 267707 476368
rect 266556 476310 267707 476312
rect 266556 476308 266562 476310
rect 267641 476307 267707 476310
rect 273294 476308 273300 476372
rect 273364 476370 273370 476372
rect 274541 476370 274607 476373
rect 276013 476372 276079 476373
rect 276013 476370 276060 476372
rect 273364 476368 274607 476370
rect 273364 476312 274546 476368
rect 274602 476312 274607 476368
rect 273364 476310 274607 476312
rect 275968 476368 276060 476370
rect 275968 476312 276018 476368
rect 275968 476310 276060 476312
rect 273364 476308 273370 476310
rect 274541 476307 274607 476310
rect 276013 476308 276060 476310
rect 276124 476308 276130 476372
rect 280153 476370 280219 476373
rect 280838 476370 280844 476372
rect 280153 476368 280844 476370
rect 280153 476312 280158 476368
rect 280214 476312 280844 476368
rect 280153 476310 280844 476312
rect 276013 476307 276079 476308
rect 280153 476307 280219 476310
rect 280838 476308 280844 476310
rect 280908 476308 280914 476372
rect 317413 476370 317479 476373
rect 318374 476370 318380 476372
rect 317413 476368 318380 476370
rect 317413 476312 317418 476368
rect 317474 476312 318380 476368
rect 317413 476310 318380 476312
rect 317413 476307 317479 476310
rect 318374 476308 318380 476310
rect 318444 476308 318450 476372
rect 320173 476370 320239 476373
rect 320950 476370 320956 476372
rect 320173 476368 320956 476370
rect 320173 476312 320178 476368
rect 320234 476312 320956 476368
rect 320173 476310 320956 476312
rect 320173 476307 320239 476310
rect 320950 476308 320956 476310
rect 321020 476308 321026 476372
rect 235901 476236 235967 476237
rect 235901 476234 235948 476236
rect 235856 476232 235948 476234
rect 235856 476176 235906 476232
rect 235856 476174 235948 476176
rect 235901 476172 235948 476174
rect 236012 476172 236018 476236
rect 237230 476172 237236 476236
rect 237300 476234 237306 476236
rect 237557 476234 237623 476237
rect 237300 476232 237623 476234
rect 237300 476176 237562 476232
rect 237618 476176 237623 476232
rect 237300 476174 237623 476176
rect 237300 476172 237306 476174
rect 235901 476171 235967 476172
rect 237557 476171 237623 476174
rect 239622 476172 239628 476236
rect 239692 476234 239698 476236
rect 240133 476234 240199 476237
rect 239692 476232 240199 476234
rect 239692 476176 240138 476232
rect 240194 476176 240199 476232
rect 239692 476174 240199 476176
rect 239692 476172 239698 476174
rect 240133 476171 240199 476174
rect 240542 476172 240548 476236
rect 240612 476234 240618 476236
rect 241421 476234 241487 476237
rect 240612 476232 241487 476234
rect 240612 476176 241426 476232
rect 241482 476176 241487 476232
rect 240612 476174 241487 476176
rect 240612 476172 240618 476174
rect 241421 476171 241487 476174
rect 241830 476172 241836 476236
rect 241900 476234 241906 476236
rect 242801 476234 242867 476237
rect 241900 476232 242867 476234
rect 241900 476176 242806 476232
rect 242862 476176 242867 476232
rect 241900 476174 242867 476176
rect 241900 476172 241906 476174
rect 242801 476171 242867 476174
rect 245653 476234 245719 476237
rect 246430 476234 246436 476236
rect 245653 476232 246436 476234
rect 245653 476176 245658 476232
rect 245714 476176 246436 476232
rect 245653 476174 246436 476176
rect 245653 476171 245719 476174
rect 246430 476172 246436 476174
rect 246500 476172 246506 476236
rect 247217 476234 247283 476237
rect 247534 476234 247540 476236
rect 247217 476232 247540 476234
rect 247217 476176 247222 476232
rect 247278 476176 247540 476232
rect 247217 476174 247540 476176
rect 247217 476171 247283 476174
rect 247534 476172 247540 476174
rect 247604 476172 247610 476236
rect 248638 476172 248644 476236
rect 248708 476234 248714 476236
rect 249793 476234 249859 476237
rect 248708 476232 249859 476234
rect 248708 476176 249798 476232
rect 249854 476176 249859 476232
rect 248708 476174 249859 476176
rect 248708 476172 248714 476174
rect 249793 476171 249859 476174
rect 250110 476172 250116 476236
rect 250180 476234 250186 476236
rect 251081 476234 251147 476237
rect 250180 476232 251147 476234
rect 250180 476176 251086 476232
rect 251142 476176 251147 476232
rect 250180 476174 251147 476176
rect 250180 476172 250186 476174
rect 251081 476171 251147 476174
rect 252318 476172 252324 476236
rect 252388 476234 252394 476236
rect 252461 476234 252527 476237
rect 252388 476232 252527 476234
rect 252388 476176 252466 476232
rect 252522 476176 252527 476232
rect 252388 476174 252527 476176
rect 252388 476172 252394 476174
rect 252461 476171 252527 476174
rect 254526 476172 254532 476236
rect 254596 476234 254602 476236
rect 255957 476234 256023 476237
rect 254596 476232 256023 476234
rect 254596 476176 255962 476232
rect 256018 476176 256023 476232
rect 254596 476174 256023 476176
rect 254596 476172 254602 476174
rect 255957 476171 256023 476174
rect 258022 476172 258028 476236
rect 258092 476234 258098 476236
rect 258165 476234 258231 476237
rect 258092 476232 258231 476234
rect 258092 476176 258170 476232
rect 258226 476176 258231 476232
rect 258092 476174 258231 476176
rect 258092 476172 258098 476174
rect 258165 476171 258231 476174
rect 259494 476172 259500 476236
rect 259564 476234 259570 476236
rect 260741 476234 260807 476237
rect 259564 476232 260807 476234
rect 259564 476176 260746 476232
rect 260802 476176 260807 476232
rect 259564 476174 260807 476176
rect 259564 476172 259570 476174
rect 260741 476171 260807 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262121 476234 262187 476237
rect 261772 476232 262187 476234
rect 261772 476176 262126 476232
rect 262182 476176 262187 476232
rect 261772 476174 262187 476176
rect 261772 476172 261778 476174
rect 262121 476171 262187 476174
rect 262806 476172 262812 476236
rect 262876 476234 262882 476236
rect 263501 476234 263567 476237
rect 262876 476232 263567 476234
rect 262876 476176 263506 476232
rect 263562 476176 263567 476232
rect 262876 476174 263567 476176
rect 262876 476172 262882 476174
rect 263501 476171 263567 476174
rect 263910 476172 263916 476236
rect 263980 476234 263986 476236
rect 264881 476234 264947 476237
rect 263980 476232 264947 476234
rect 263980 476176 264886 476232
rect 264942 476176 264947 476232
rect 263980 476174 264947 476176
rect 263980 476172 263986 476174
rect 264881 476171 264947 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266261 476234 266327 476237
rect 267549 476236 267615 476237
rect 267549 476234 267596 476236
rect 265452 476232 266327 476234
rect 265452 476176 266266 476232
rect 266322 476176 266327 476232
rect 265452 476174 266327 476176
rect 267504 476232 267596 476234
rect 267504 476176 267554 476232
rect 267504 476174 267596 476176
rect 265452 476172 265458 476174
rect 266261 476171 266327 476174
rect 267549 476172 267596 476174
rect 267660 476172 267666 476236
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 267549 476171 267615 476172
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271781 476234 271847 476237
rect 274449 476236 274515 476237
rect 275921 476236 275987 476237
rect 271340 476232 271847 476234
rect 271340 476176 271786 476232
rect 271842 476176 271847 476232
rect 271340 476174 271847 476176
rect 271340 476172 271346 476174
rect 271781 476171 271847 476174
rect 274398 476172 274404 476236
rect 274468 476234 274515 476236
rect 274468 476232 274560 476234
rect 274510 476176 274560 476232
rect 274468 476174 274560 476176
rect 274468 476172 274515 476174
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277301 476234 277367 476237
rect 277044 476232 277367 476234
rect 277044 476176 277306 476232
rect 277362 476176 277367 476232
rect 277044 476174 277367 476176
rect 277044 476172 277050 476174
rect 274449 476171 274515 476172
rect 275921 476171 275987 476172
rect 277301 476171 277367 476174
rect 278078 476172 278084 476236
rect 278148 476234 278154 476236
rect 278681 476234 278747 476237
rect 278148 476232 278747 476234
rect 278148 476176 278686 476232
rect 278742 476176 278747 476232
rect 278148 476174 278747 476176
rect 278148 476172 278154 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 283005 476234 283071 476237
rect 283414 476234 283420 476236
rect 283005 476232 283420 476234
rect 283005 476176 283010 476232
rect 283066 476176 283420 476232
rect 283005 476174 283420 476176
rect 283005 476171 283071 476174
rect 283414 476172 283420 476174
rect 283484 476172 283490 476236
rect 285857 476234 285923 476237
rect 285990 476234 285996 476236
rect 285857 476232 285996 476234
rect 285857 476176 285862 476232
rect 285918 476176 285996 476232
rect 285857 476174 285996 476176
rect 285857 476171 285923 476174
rect 285990 476172 285996 476174
rect 286060 476172 286066 476236
rect 287237 476234 287303 476237
rect 288198 476234 288204 476236
rect 287237 476232 288204 476234
rect 287237 476176 287242 476232
rect 287298 476176 288204 476232
rect 287237 476174 288204 476176
rect 287237 476171 287303 476174
rect 288198 476172 288204 476174
rect 288268 476172 288274 476236
rect 289813 476234 289879 476237
rect 290958 476234 290964 476236
rect 289813 476232 290964 476234
rect 289813 476176 289818 476232
rect 289874 476176 290964 476232
rect 289813 476174 290964 476176
rect 289813 476171 289879 476174
rect 290958 476172 290964 476174
rect 291028 476172 291034 476236
rect 292665 476234 292731 476237
rect 293350 476234 293356 476236
rect 292665 476232 293356 476234
rect 292665 476176 292670 476232
rect 292726 476176 293356 476232
rect 292665 476174 293356 476176
rect 292665 476171 292731 476174
rect 293350 476172 293356 476174
rect 293420 476172 293426 476236
rect 295333 476234 295399 476237
rect 295926 476234 295932 476236
rect 295333 476232 295932 476234
rect 295333 476176 295338 476232
rect 295394 476176 295932 476232
rect 295333 476174 295932 476176
rect 295333 476171 295399 476174
rect 295926 476172 295932 476174
rect 295996 476172 296002 476236
rect 298093 476234 298159 476237
rect 300853 476236 300919 476237
rect 298502 476234 298508 476236
rect 298093 476232 298508 476234
rect 298093 476176 298098 476232
rect 298154 476176 298508 476232
rect 298093 476174 298508 476176
rect 298093 476171 298159 476174
rect 298502 476172 298508 476174
rect 298572 476172 298578 476236
rect 300853 476234 300900 476236
rect 300808 476232 300900 476234
rect 300808 476176 300858 476232
rect 300808 476174 300900 476176
rect 300853 476172 300900 476174
rect 300964 476172 300970 476236
rect 325785 476234 325851 476237
rect 325918 476234 325924 476236
rect 325785 476232 325924 476234
rect 325785 476176 325790 476232
rect 325846 476176 325924 476232
rect 325785 476174 325924 476176
rect 300853 476171 300919 476172
rect 325785 476171 325851 476174
rect 325918 476172 325924 476174
rect 325988 476172 325994 476236
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 583520 471324 584960 471564
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 295977 444818 296043 444821
rect 538857 444818 538923 444821
rect 295977 444816 538923 444818
rect 295977 444760 295982 444816
rect 296038 444760 538862 444816
rect 538918 444760 538923 444816
rect 295977 444758 538923 444760
rect 295977 444755 296043 444758
rect 538857 444755 538923 444758
rect 294413 444682 294479 444685
rect 342253 444682 342319 444685
rect 294413 444680 342319 444682
rect 294413 444624 294418 444680
rect 294474 444624 342258 444680
rect 342314 444624 342319 444680
rect 583520 444668 584960 444908
rect 294413 444622 342319 444624
rect 294413 444619 294479 444622
rect 342253 444619 342319 444622
rect 295149 444546 295215 444549
rect 368974 444546 368980 444548
rect 295149 444544 368980 444546
rect 295149 444488 295154 444544
rect 295210 444488 368980 444544
rect 295149 444486 368980 444488
rect 295149 444483 295215 444486
rect 368974 444484 368980 444486
rect 369044 444484 369050 444548
rect 299749 443322 299815 443325
rect 363454 443322 363460 443324
rect 299749 443320 363460 443322
rect 299749 443264 299754 443320
rect 299810 443264 363460 443320
rect 299749 443262 363460 443264
rect 299749 443259 299815 443262
rect 363454 443260 363460 443262
rect 363524 443260 363530 443324
rect 214598 443124 214604 443188
rect 214668 443186 214674 443188
rect 345289 443186 345355 443189
rect 214668 443184 345355 443186
rect 214668 443128 345294 443184
rect 345350 443128 345355 443184
rect 214668 443126 345355 443128
rect 214668 443124 214674 443126
rect 345289 443123 345355 443126
rect 215886 442988 215892 443052
rect 215956 443050 215962 443052
rect 347589 443050 347655 443053
rect 215956 443048 347655 443050
rect 215956 442992 347594 443048
rect 347650 442992 347655 443048
rect 215956 442990 347655 442992
rect 215956 442988 215962 442990
rect 347589 442987 347655 442990
rect 307017 442234 307083 442237
rect 307017 442232 311910 442234
rect 307017 442176 307022 442232
rect 307078 442176 311910 442232
rect 307017 442174 311910 442176
rect 307017 442171 307083 442174
rect 311850 441690 311910 442174
rect 360326 442172 360332 442236
rect 360396 442234 360402 442236
rect 361205 442234 361271 442237
rect 360396 442232 361271 442234
rect 360396 442176 361210 442232
rect 361266 442176 361271 442232
rect 360396 442174 361271 442176
rect 360396 442172 360402 442174
rect 361205 442171 361271 442174
rect 361614 442172 361620 442236
rect 361684 442234 361690 442236
rect 361941 442234 362007 442237
rect 361684 442232 362007 442234
rect 361684 442176 361946 442232
rect 362002 442176 362007 442232
rect 361684 442174 362007 442176
rect 361684 442172 361690 442174
rect 361941 442171 362007 442174
rect 363822 441690 363828 441692
rect 311850 441630 363828 441690
rect 363822 441628 363828 441630
rect 363892 441628 363898 441692
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 2865 397490 2931 397493
rect -960 397488 2931 397490
rect -960 397432 2870 397488
rect 2926 397432 2931 397488
rect -960 397430 2931 397432
rect -960 397340 480 397430
rect 2865 397427 2931 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2865 371378 2931 371381
rect -960 371376 2931 371378
rect -960 371320 2870 371376
rect 2926 371320 2931 371376
rect -960 371318 2931 371320
rect -960 371228 480 371318
rect 2865 371315 2931 371318
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3969 345402 4035 345405
rect -960 345400 4035 345402
rect -960 345344 3974 345400
rect 4030 345344 4035 345400
rect -960 345342 4035 345344
rect -960 345252 480 345342
rect 3969 345339 4035 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580625 325274 580691 325277
rect 583520 325274 584960 325364
rect 580625 325272 584960 325274
rect 580625 325216 580630 325272
rect 580686 325216 584960 325272
rect 580625 325214 584960 325216
rect 580625 325211 580691 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 583520 311932 584960 312172
rect 345105 309090 345171 309093
rect 363689 309090 363755 309093
rect 345105 309088 363755 309090
rect 345105 309032 345110 309088
rect 345166 309032 363694 309088
rect 363750 309032 363755 309088
rect 345105 309030 363755 309032
rect 345105 309027 345171 309030
rect 363689 309027 363755 309030
rect 219014 308892 219020 308956
rect 219084 308954 219090 308956
rect 275185 308954 275251 308957
rect 219084 308952 275251 308954
rect 219084 308896 275190 308952
rect 275246 308896 275251 308952
rect 219084 308894 275251 308896
rect 219084 308892 219090 308894
rect 275185 308891 275251 308894
rect 346025 308954 346091 308957
rect 363781 308954 363847 308957
rect 346025 308952 363847 308954
rect 346025 308896 346030 308952
rect 346086 308896 363786 308952
rect 363842 308896 363847 308952
rect 346025 308894 363847 308896
rect 346025 308891 346091 308894
rect 363781 308891 363847 308894
rect 218830 308756 218836 308820
rect 218900 308818 218906 308820
rect 276565 308818 276631 308821
rect 218900 308816 276631 308818
rect 218900 308760 276570 308816
rect 276626 308760 276631 308816
rect 218900 308758 276631 308760
rect 218900 308756 218906 308758
rect 276565 308755 276631 308758
rect 298461 308818 298527 308821
rect 362401 308818 362467 308821
rect 298461 308816 362467 308818
rect 298461 308760 298466 308816
rect 298522 308760 362406 308816
rect 362462 308760 362467 308816
rect 298461 308758 362467 308760
rect 298461 308755 298527 308758
rect 362401 308755 362467 308758
rect 217358 308620 217364 308684
rect 217428 308682 217434 308684
rect 275921 308682 275987 308685
rect 217428 308680 275987 308682
rect 217428 308624 275926 308680
rect 275982 308624 275987 308680
rect 217428 308622 275987 308624
rect 217428 308620 217434 308622
rect 275921 308619 275987 308622
rect 294413 308682 294479 308685
rect 365805 308682 365871 308685
rect 294413 308680 365871 308682
rect 294413 308624 294418 308680
rect 294474 308624 365810 308680
rect 365866 308624 365871 308680
rect 294413 308622 365871 308624
rect 294413 308619 294479 308622
rect 365805 308619 365871 308622
rect 217542 308484 217548 308548
rect 217612 308546 217618 308548
rect 277209 308546 277275 308549
rect 217612 308544 277275 308546
rect 217612 308488 277214 308544
rect 277270 308488 277275 308544
rect 217612 308486 277275 308488
rect 217612 308484 217618 308486
rect 277209 308483 277275 308486
rect 325049 308546 325115 308549
rect 431217 308546 431283 308549
rect 325049 308544 431283 308546
rect 325049 308488 325054 308544
rect 325110 308488 431222 308544
rect 431278 308488 431283 308544
rect 325049 308486 431283 308488
rect 325049 308483 325115 308486
rect 431217 308483 431283 308486
rect 75177 308410 75243 308413
rect 233233 308410 233299 308413
rect 75177 308408 233299 308410
rect 75177 308352 75182 308408
rect 75238 308352 233238 308408
rect 233294 308352 233299 308408
rect 75177 308350 233299 308352
rect 75177 308347 75243 308350
rect 233233 308347 233299 308350
rect 323669 308410 323735 308413
rect 471973 308410 472039 308413
rect 323669 308408 472039 308410
rect 323669 308352 323674 308408
rect 323730 308352 471978 308408
rect 472034 308352 472039 308408
rect 323669 308350 472039 308352
rect 323669 308347 323735 308350
rect 471973 308347 472039 308350
rect 358629 306370 358695 306373
rect 360101 306370 360167 306373
rect 358629 306368 360167 306370
rect -960 306234 480 306324
rect 358629 306312 358634 306368
rect 358690 306312 360106 306368
rect 360162 306312 360167 306368
rect 358629 306310 360167 306312
rect 358629 306307 358695 306310
rect 360101 306307 360167 306310
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 216070 306172 216076 306236
rect 216140 306234 216146 306236
rect 275645 306234 275711 306237
rect 216140 306232 275711 306234
rect 216140 306176 275650 306232
rect 275706 306176 275711 306232
rect 216140 306174 275711 306176
rect 216140 306172 216146 306174
rect 275645 306171 275711 306174
rect 348141 306234 348207 306237
rect 369025 306234 369091 306237
rect 348141 306232 369091 306234
rect 348141 306176 348146 306232
rect 348202 306176 369030 306232
rect 369086 306176 369091 306232
rect 348141 306174 369091 306176
rect 348141 306171 348207 306174
rect 369025 306171 369091 306174
rect 214966 306036 214972 306100
rect 215036 306098 215042 306100
rect 275001 306098 275067 306101
rect 215036 306096 275067 306098
rect 215036 306040 275006 306096
rect 275062 306040 275067 306096
rect 215036 306038 275067 306040
rect 215036 306036 215042 306038
rect 275001 306035 275067 306038
rect 311341 306098 311407 306101
rect 407113 306098 407179 306101
rect 311341 306096 407179 306098
rect 311341 306040 311346 306096
rect 311402 306040 407118 306096
rect 407174 306040 407179 306096
rect 311341 306038 407179 306040
rect 311341 306035 311407 306038
rect 407113 306035 407179 306038
rect 216254 305900 216260 305964
rect 216324 305962 216330 305964
rect 277485 305962 277551 305965
rect 216324 305960 277551 305962
rect 216324 305904 277490 305960
rect 277546 305904 277551 305960
rect 216324 305902 277551 305904
rect 216324 305900 216330 305902
rect 277485 305899 277551 305902
rect 313641 305962 313707 305965
rect 418153 305962 418219 305965
rect 313641 305960 418219 305962
rect 313641 305904 313646 305960
rect 313702 305904 418158 305960
rect 418214 305904 418219 305960
rect 313641 305902 418219 305904
rect 313641 305899 313707 305902
rect 418153 305899 418219 305902
rect 216990 305764 216996 305828
rect 217060 305826 217066 305828
rect 280889 305826 280955 305829
rect 217060 305824 280955 305826
rect 217060 305768 280894 305824
rect 280950 305768 280955 305824
rect 217060 305766 280955 305768
rect 217060 305764 217066 305766
rect 280889 305763 280955 305766
rect 330201 305826 330267 305829
rect 442257 305826 442323 305829
rect 330201 305824 442323 305826
rect 330201 305768 330206 305824
rect 330262 305768 442262 305824
rect 442318 305768 442323 305824
rect 330201 305766 442323 305768
rect 330201 305763 330267 305766
rect 442257 305763 442323 305766
rect 217174 305628 217180 305692
rect 217244 305690 217250 305692
rect 280705 305690 280771 305693
rect 217244 305688 280771 305690
rect 217244 305632 280710 305688
rect 280766 305632 280771 305688
rect 217244 305630 280771 305632
rect 217244 305628 217250 305630
rect 280705 305627 280771 305630
rect 326061 305690 326127 305693
rect 483013 305690 483079 305693
rect 326061 305688 483079 305690
rect 326061 305632 326066 305688
rect 326122 305632 483018 305688
rect 483074 305632 483079 305688
rect 326061 305630 483079 305632
rect 326061 305627 326127 305630
rect 483013 305627 483079 305630
rect 309777 304194 309843 304197
rect 369158 304194 369164 304196
rect 309777 304192 369164 304194
rect 309777 304136 309782 304192
rect 309838 304136 369164 304192
rect 309777 304134 369164 304136
rect 309777 304131 309843 304134
rect 369158 304132 369164 304134
rect 369228 304132 369234 304196
rect 210877 303378 210943 303381
rect 274725 303378 274791 303381
rect 210877 303376 274791 303378
rect 210877 303320 210882 303376
rect 210938 303320 274730 303376
rect 274786 303320 274791 303376
rect 210877 303318 274791 303320
rect 210877 303315 210943 303318
rect 274725 303315 274791 303318
rect 211889 303242 211955 303245
rect 277025 303242 277091 303245
rect 211889 303240 277091 303242
rect 211889 303184 211894 303240
rect 211950 303184 277030 303240
rect 277086 303184 277091 303240
rect 211889 303182 277091 303184
rect 211889 303179 211955 303182
rect 277025 303179 277091 303182
rect 307845 303242 307911 303245
rect 363638 303242 363644 303244
rect 307845 303240 363644 303242
rect 307845 303184 307850 303240
rect 307906 303184 363644 303240
rect 307845 303182 363644 303184
rect 307845 303179 307911 303182
rect 363638 303180 363644 303182
rect 363708 303180 363714 303244
rect 212942 303044 212948 303108
rect 213012 303106 213018 303108
rect 278405 303106 278471 303109
rect 213012 303104 278471 303106
rect 213012 303048 278410 303104
rect 278466 303048 278471 303104
rect 213012 303046 278471 303048
rect 213012 303044 213018 303046
rect 278405 303043 278471 303046
rect 308581 303106 308647 303109
rect 367686 303106 367692 303108
rect 308581 303104 367692 303106
rect 308581 303048 308586 303104
rect 308642 303048 367692 303104
rect 308581 303046 367692 303048
rect 308581 303043 308647 303046
rect 367686 303044 367692 303046
rect 367756 303044 367762 303108
rect 212073 302970 212139 302973
rect 277669 302970 277735 302973
rect 212073 302968 277735 302970
rect 212073 302912 212078 302968
rect 212134 302912 277674 302968
rect 277730 302912 277735 302968
rect 212073 302910 277735 302912
rect 212073 302907 212139 302910
rect 277669 302907 277735 302910
rect 307201 302970 307267 302973
rect 386413 302970 386479 302973
rect 307201 302968 386479 302970
rect 307201 302912 307206 302968
rect 307262 302912 386418 302968
rect 386474 302912 386479 302968
rect 307201 302910 386479 302912
rect 307201 302907 307267 302910
rect 386413 302907 386479 302910
rect 212257 302834 212323 302837
rect 279049 302834 279115 302837
rect 212257 302832 279115 302834
rect 212257 302776 212262 302832
rect 212318 302776 279054 302832
rect 279110 302776 279115 302832
rect 212257 302774 279115 302776
rect 212257 302771 212323 302774
rect 279049 302771 279115 302774
rect 312629 302834 312695 302837
rect 415393 302834 415459 302837
rect 312629 302832 415459 302834
rect 312629 302776 312634 302832
rect 312690 302776 415398 302832
rect 415454 302776 415459 302832
rect 312629 302774 415459 302776
rect 312629 302771 312695 302774
rect 415393 302771 415459 302774
rect 305637 301474 305703 301477
rect 364926 301474 364932 301476
rect 305637 301472 364932 301474
rect 305637 301416 305642 301472
rect 305698 301416 364932 301472
rect 305637 301414 364932 301416
rect 305637 301411 305703 301414
rect 364926 301412 364932 301414
rect 364996 301412 365002 301476
rect 218789 300386 218855 300389
rect 283281 300386 283347 300389
rect 218789 300384 283347 300386
rect 218789 300328 218794 300384
rect 218850 300328 283286 300384
rect 283342 300328 283347 300384
rect 218789 300326 283347 300328
rect 218789 300323 218855 300326
rect 283281 300323 283347 300326
rect 214741 300250 214807 300253
rect 283097 300250 283163 300253
rect 214741 300248 283163 300250
rect 214741 300192 214746 300248
rect 214802 300192 283102 300248
rect 283158 300192 283163 300248
rect 214741 300190 283163 300192
rect 214741 300187 214807 300190
rect 283097 300187 283163 300190
rect 210969 300114 211035 300117
rect 284569 300114 284635 300117
rect 210969 300112 284635 300114
rect 210969 300056 210974 300112
rect 211030 300056 284574 300112
rect 284630 300056 284635 300112
rect 210969 300054 284635 300056
rect 210969 300051 211035 300054
rect 284569 300051 284635 300054
rect 583520 298604 584960 298844
rect 303981 297394 304047 297397
rect 368422 297394 368428 297396
rect 303981 297392 368428 297394
rect 303981 297336 303986 297392
rect 304042 297336 368428 297392
rect 303981 297334 368428 297336
rect 303981 297331 304047 297334
rect 368422 297332 368428 297334
rect 368492 297332 368498 297396
rect -960 293178 480 293268
rect 3877 293178 3943 293181
rect -960 293176 3943 293178
rect -960 293120 3882 293176
rect 3938 293120 3943 293176
rect -960 293118 3943 293120
rect -960 293028 480 293118
rect 3877 293115 3943 293118
rect 583520 285276 584960 285516
rect 302693 283522 302759 283525
rect 367134 283522 367140 283524
rect 302693 283520 367140 283522
rect 302693 283464 302698 283520
rect 302754 283464 367140 283520
rect 302693 283462 367140 283464
rect 302693 283459 302759 283462
rect 367134 283460 367140 283462
rect 367204 283460 367210 283524
rect 302601 282162 302667 282165
rect 364374 282162 364380 282164
rect 302601 282160 364380 282162
rect 302601 282104 302606 282160
rect 302662 282104 364380 282160
rect 302601 282102 364380 282104
rect 302601 282099 302667 282102
rect 364374 282100 364380 282102
rect 364444 282100 364450 282164
rect -960 279972 480 280212
rect 216438 275164 216444 275228
rect 216508 275226 216514 275228
rect 273621 275226 273687 275229
rect 216508 275224 273687 275226
rect 216508 275168 273626 275224
rect 273682 275168 273687 275224
rect 216508 275166 273687 275168
rect 216508 275164 216514 275166
rect 273621 275163 273687 275166
rect 214414 273804 214420 273868
rect 214484 273866 214490 273868
rect 272149 273866 272215 273869
rect 214484 273864 272215 273866
rect 214484 273808 272154 273864
rect 272210 273808 272215 273864
rect 214484 273806 272215 273808
rect 214484 273804 214490 273806
rect 272149 273803 272215 273806
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 303705 269786 303771 269789
rect 369894 269786 369900 269788
rect 303705 269784 369900 269786
rect 303705 269728 303710 269784
rect 303766 269728 369900 269784
rect 303705 269726 369900 269728
rect 303705 269723 303771 269726
rect 369894 269724 369900 269726
rect 369964 269724 369970 269788
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 215150 267004 215156 267068
rect 215220 267066 215226 267068
rect 273529 267066 273595 267069
rect 215220 267064 273595 267066
rect 215220 267008 273534 267064
rect 273590 267008 273595 267064
rect 215220 267006 273595 267008
rect 215220 267004 215226 267006
rect 273529 267003 273595 267006
rect 302325 265570 302391 265573
rect 362902 265570 362908 265572
rect 302325 265568 362908 265570
rect 302325 265512 302330 265568
rect 302386 265512 362908 265568
rect 302325 265510 362908 265512
rect 302325 265507 302391 265510
rect 362902 265508 362908 265510
rect 362972 265508 362978 265572
rect 301313 264210 301379 264213
rect 358854 264210 358860 264212
rect 301313 264208 358860 264210
rect 301313 264152 301318 264208
rect 301374 264152 358860 264208
rect 301313 264150 358860 264152
rect 301313 264147 301379 264150
rect 358854 264148 358860 264150
rect 358924 264148 358930 264212
rect 219198 262788 219204 262852
rect 219268 262850 219274 262852
rect 273437 262850 273503 262853
rect 219268 262848 273503 262850
rect 219268 262792 273442 262848
rect 273498 262792 273503 262848
rect 219268 262790 273503 262792
rect 219268 262788 219274 262790
rect 273437 262787 273503 262790
rect 583520 258756 584960 258996
rect 302233 254690 302299 254693
rect 362534 254690 362540 254692
rect 302233 254688 362540 254690
rect 302233 254632 302238 254688
rect 302294 254632 362540 254688
rect 302233 254630 362540 254632
rect 302233 254627 302299 254630
rect 362534 254628 362540 254630
rect 362604 254628 362610 254692
rect 302417 254554 302483 254557
rect 365662 254554 365668 254556
rect 302417 254552 365668 254554
rect 302417 254496 302422 254552
rect 302478 254496 365668 254552
rect 302417 254494 365668 254496
rect 302417 254491 302483 254494
rect 365662 254492 365668 254494
rect 365732 254492 365738 254556
rect -960 254146 480 254236
rect 2865 254146 2931 254149
rect -960 254144 2931 254146
rect -960 254088 2870 254144
rect 2926 254088 2931 254144
rect -960 254086 2931 254088
rect -960 253996 480 254086
rect 2865 254083 2931 254086
rect 299841 250882 299907 250885
rect 367318 250882 367324 250884
rect 299841 250880 367324 250882
rect 299841 250824 299846 250880
rect 299902 250824 367324 250880
rect 299841 250822 367324 250824
rect 299841 250819 299907 250822
rect 367318 250820 367324 250822
rect 367388 250820 367394 250884
rect 306373 250746 306439 250749
rect 385033 250746 385099 250749
rect 306373 250744 385099 250746
rect 306373 250688 306378 250744
rect 306434 250688 385038 250744
rect 385094 250688 385099 250744
rect 306373 250686 385099 250688
rect 306373 250683 306439 250686
rect 385033 250683 385099 250686
rect 316033 250610 316099 250613
rect 434713 250610 434779 250613
rect 316033 250608 434779 250610
rect 316033 250552 316038 250608
rect 316094 250552 434718 250608
rect 434774 250552 434779 250608
rect 316033 250550 434779 250552
rect 316033 250547 316099 250550
rect 434713 250547 434779 250550
rect 336825 250474 336891 250477
rect 546493 250474 546559 250477
rect 336825 250472 546559 250474
rect 336825 250416 336830 250472
rect 336886 250416 546498 250472
rect 546554 250416 546559 250472
rect 336825 250414 546559 250416
rect 336825 250411 336891 250414
rect 546493 250411 546559 250414
rect 213126 249052 213132 249116
rect 213196 249114 213202 249116
rect 273345 249114 273411 249117
rect 213196 249112 273411 249114
rect 213196 249056 273350 249112
rect 273406 249056 273411 249112
rect 213196 249054 273411 249056
rect 213196 249052 213202 249054
rect 273345 249051 273411 249054
rect 299565 248162 299631 248165
rect 364558 248162 364564 248164
rect 299565 248160 364564 248162
rect 299565 248104 299570 248160
rect 299626 248104 364564 248160
rect 299565 248102 364564 248104
rect 299565 248099 299631 248102
rect 364558 248100 364564 248102
rect 364628 248100 364634 248164
rect 321553 248026 321619 248029
rect 465165 248026 465231 248029
rect 321553 248024 465231 248026
rect 321553 247968 321558 248024
rect 321614 247968 465170 248024
rect 465226 247968 465231 248024
rect 321553 247966 465231 247968
rect 321553 247963 321619 247966
rect 465165 247963 465231 247966
rect 323117 247890 323183 247893
rect 469213 247890 469279 247893
rect 323117 247888 469279 247890
rect 323117 247832 323122 247888
rect 323178 247832 469218 247888
rect 469274 247832 469279 247888
rect 323117 247830 469279 247832
rect 323117 247827 323183 247830
rect 469213 247827 469279 247830
rect 322933 247754 322999 247757
rect 473445 247754 473511 247757
rect 322933 247752 473511 247754
rect 322933 247696 322938 247752
rect 322994 247696 473450 247752
rect 473506 247696 473511 247752
rect 322933 247694 473511 247696
rect 322933 247691 322999 247694
rect 473445 247691 473511 247694
rect 332593 247618 332659 247621
rect 523125 247618 523191 247621
rect 332593 247616 523191 247618
rect 332593 247560 332598 247616
rect 332654 247560 523130 247616
rect 523186 247560 523191 247616
rect 332593 247558 523191 247560
rect 332593 247555 332659 247558
rect 523125 247555 523191 247558
rect 301037 246258 301103 246261
rect 360142 246258 360148 246260
rect 301037 246256 360148 246258
rect 301037 246200 301042 246256
rect 301098 246200 360148 246256
rect 301037 246198 360148 246200
rect 301037 246195 301103 246198
rect 360142 246196 360148 246198
rect 360212 246196 360218 246260
rect 299473 245578 299539 245581
rect 356881 245578 356947 245581
rect 299473 245576 356947 245578
rect 299473 245520 299478 245576
rect 299534 245520 356886 245576
rect 356942 245520 356947 245576
rect 299473 245518 356947 245520
rect 299473 245515 299539 245518
rect 356881 245515 356947 245518
rect 357433 245578 357499 245581
rect 358118 245578 358124 245580
rect 357433 245576 358124 245578
rect 357433 245520 357438 245576
rect 357494 245520 358124 245576
rect 357433 245518 358124 245520
rect 357433 245515 357499 245518
rect 358118 245516 358124 245518
rect 358188 245516 358194 245580
rect 296713 245442 296779 245445
rect 358169 245442 358235 245445
rect 358302 245442 358308 245444
rect 296713 245440 356530 245442
rect 296713 245384 296718 245440
rect 296774 245384 356530 245440
rect 296713 245382 356530 245384
rect 296713 245379 296779 245382
rect 298093 245306 298159 245309
rect 356329 245306 356395 245309
rect 298093 245304 356395 245306
rect 298093 245248 298098 245304
rect 298154 245248 356334 245304
rect 356390 245248 356395 245304
rect 298093 245246 356395 245248
rect 356470 245306 356530 245382
rect 358169 245440 358308 245442
rect 358169 245384 358174 245440
rect 358230 245384 358308 245440
rect 358169 245382 358308 245384
rect 358169 245379 358235 245382
rect 358302 245380 358308 245382
rect 358372 245380 358378 245444
rect 583520 245428 584960 245668
rect 358486 245306 358492 245308
rect 356470 245246 358492 245306
rect 298093 245243 298159 245246
rect 356329 245243 356395 245246
rect 358486 245244 358492 245246
rect 358556 245244 358562 245308
rect 296897 245170 296963 245173
rect 356605 245170 356671 245173
rect 296897 245168 356671 245170
rect 296897 245112 296902 245168
rect 296958 245112 356610 245168
rect 356666 245112 356671 245168
rect 296897 245110 356671 245112
rect 296897 245107 296963 245110
rect 356605 245107 356671 245110
rect 356881 245170 356947 245173
rect 359038 245170 359044 245172
rect 356881 245168 359044 245170
rect 356881 245112 356886 245168
rect 356942 245112 359044 245168
rect 356881 245110 359044 245112
rect 356881 245107 356947 245110
rect 359038 245108 359044 245110
rect 359108 245108 359114 245172
rect 295333 245034 295399 245037
rect 359222 245034 359228 245036
rect 295333 245032 359228 245034
rect 295333 244976 295338 245032
rect 295394 244976 359228 245032
rect 295333 244974 359228 244976
rect 295333 244971 295399 244974
rect 359222 244972 359228 244974
rect 359292 244972 359298 245036
rect 295517 244898 295583 244901
rect 359406 244898 359412 244900
rect 295517 244896 359412 244898
rect 295517 244840 295522 244896
rect 295578 244840 359412 244896
rect 295517 244838 359412 244840
rect 295517 244835 295583 244838
rect 359406 244836 359412 244838
rect 359476 244836 359482 244900
rect 299657 244762 299723 244765
rect 357566 244762 357572 244764
rect 299657 244760 357572 244762
rect 299657 244704 299662 244760
rect 299718 244704 357572 244760
rect 299657 244702 357572 244704
rect 299657 244699 299723 244702
rect 357566 244700 357572 244702
rect 357636 244700 357642 244764
rect 356329 244626 356395 244629
rect 360510 244626 360516 244628
rect 356329 244624 360516 244626
rect 356329 244568 356334 244624
rect 356390 244568 360516 244624
rect 356329 244566 360516 244568
rect 356329 244563 356395 244566
rect 360510 244564 360516 244566
rect 360580 244564 360586 244628
rect 356605 244490 356671 244493
rect 360694 244490 360700 244492
rect 356605 244488 360700 244490
rect 356605 244432 356610 244488
rect 356666 244432 360700 244488
rect 356605 244430 360700 244432
rect 356605 244427 356671 244430
rect 360694 244428 360700 244430
rect 360764 244428 360770 244492
rect 355501 243946 355567 243949
rect 363413 243946 363479 243949
rect 355501 243944 363479 243946
rect 355501 243888 355506 243944
rect 355562 243888 363418 243944
rect 363474 243888 363479 243944
rect 355501 243886 363479 243888
rect 355501 243883 355567 243886
rect 363413 243883 363479 243886
rect 218421 243538 218487 243541
rect 218646 243538 218652 243540
rect 218421 243536 218652 243538
rect 218421 243480 218426 243536
rect 218482 243480 218652 243536
rect 218421 243478 218652 243480
rect 218421 243475 218487 243478
rect 218646 243476 218652 243478
rect 218716 243476 218722 243540
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 580533 232386 580599 232389
rect 583520 232386 584960 232476
rect 580533 232384 584960 232386
rect 580533 232328 580538 232384
rect 580594 232328 584960 232384
rect 580533 232326 584960 232328
rect 580533 232323 580599 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect -960 214918 674 214978
rect -960 214842 480 214918
rect 614 214842 674 214918
rect -960 214828 674 214842
rect 246 214782 674 214828
rect 246 214298 306 214782
rect 246 214238 6930 214298
rect 6870 214026 6930 214238
rect 214598 214026 214604 214028
rect 6870 213966 214604 214026
rect 214598 213964 214604 213966
rect 214668 213964 214674 214028
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 217501 196890 217567 196893
rect 219390 196890 220064 196924
rect 217501 196888 220064 196890
rect 217501 196832 217506 196888
rect 217562 196864 220064 196888
rect 217562 196832 219450 196864
rect 217501 196830 219450 196832
rect 217501 196827 217567 196830
rect 217409 195938 217475 195941
rect 219390 195938 220064 195972
rect 217409 195936 220064 195938
rect 217409 195880 217414 195936
rect 217470 195912 220064 195936
rect 217470 195880 219450 195912
rect 217409 195878 219450 195880
rect 217409 195875 217475 195878
rect 217041 193762 217107 193765
rect 219390 193762 220064 193796
rect 217041 193760 220064 193762
rect 217041 193704 217046 193760
rect 217102 193736 220064 193760
rect 217102 193704 219450 193736
rect 217041 193702 219450 193704
rect 217041 193699 217107 193702
rect 216673 192810 216739 192813
rect 219390 192810 220064 192844
rect 216673 192808 220064 192810
rect 216673 192752 216678 192808
rect 216734 192784 220064 192808
rect 216734 192752 219450 192784
rect 216673 192750 219450 192752
rect 216673 192747 216739 192750
rect 583520 192538 584960 192628
rect 583342 192478 584960 192538
rect 583342 192402 583402 192478
rect 583520 192402 584960 192478
rect 583342 192388 584960 192402
rect 583342 192342 583586 192388
rect 363822 191796 363828 191860
rect 363892 191858 363898 191860
rect 583526 191858 583586 192342
rect 363892 191798 583586 191858
rect 363892 191796 363898 191798
rect 218513 191042 218579 191045
rect 219390 191042 220064 191076
rect 218513 191040 220064 191042
rect 218513 190984 218518 191040
rect 218574 191016 220064 191040
rect 218574 190984 219450 191016
rect 218513 190982 219450 190984
rect 218513 190979 218579 190982
rect 218697 189954 218763 189957
rect 219390 189954 220064 189988
rect 218697 189952 220064 189954
rect 218697 189896 218702 189952
rect 218758 189928 220064 189952
rect 218758 189896 219450 189928
rect 218697 189894 219450 189896
rect 218697 189891 218763 189894
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 216673 188186 216739 188189
rect 219390 188186 220064 188220
rect 216673 188184 220064 188186
rect 216673 188128 216678 188184
rect 216734 188160 220064 188184
rect 216734 188128 219450 188160
rect 216673 188126 219450 188128
rect 216673 188123 216739 188126
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 217225 169962 217291 169965
rect 219390 169962 220064 169996
rect 217225 169960 220064 169962
rect 217225 169904 217230 169960
rect 217286 169936 220064 169960
rect 217286 169904 219450 169936
rect 217225 169902 219450 169904
rect 217225 169899 217291 169902
rect 217685 168330 217751 168333
rect 219390 168330 220064 168364
rect 217685 168328 220064 168330
rect 217685 168272 217690 168328
rect 217746 168304 220064 168328
rect 217746 168272 219450 168304
rect 217685 168270 219450 168272
rect 217685 168267 217751 168270
rect 217593 168058 217659 168061
rect 219390 168058 220064 168092
rect 217593 168056 220064 168058
rect 217593 168000 217598 168056
rect 217654 168032 220064 168056
rect 217654 168000 219450 168032
rect 217593 167998 219450 168000
rect 217593 167995 217659 167998
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 215886 162890 215892 162892
rect -960 162830 215892 162890
rect -960 162740 480 162830
rect 215886 162828 215892 162830
rect 215956 162828 215962 162892
rect 277025 159900 277091 159901
rect 278129 159900 278195 159901
rect 279233 159900 279299 159901
rect 276984 159898 276990 159900
rect 276934 159838 276990 159898
rect 277054 159896 277091 159900
rect 278072 159898 278078 159900
rect 277086 159840 277091 159896
rect 276984 159836 276990 159838
rect 277054 159836 277091 159840
rect 278038 159838 278078 159898
rect 278142 159896 278195 159900
rect 279160 159898 279166 159900
rect 278190 159840 278195 159896
rect 278072 159836 278078 159838
rect 278142 159836 278195 159840
rect 279142 159838 279166 159898
rect 279160 159836 279166 159838
rect 279230 159896 279299 159900
rect 279230 159840 279238 159896
rect 279294 159840 279299 159896
rect 279230 159836 279299 159840
rect 277025 159835 277091 159836
rect 278129 159835 278195 159836
rect 279233 159835 279299 159836
rect 285949 159900 286015 159901
rect 285949 159896 285966 159900
rect 286030 159898 286036 159900
rect 285949 159840 285954 159896
rect 285949 159836 285966 159840
rect 286030 159838 286106 159898
rect 286030 159836 286036 159838
rect 285949 159835 286015 159836
rect 256049 159628 256115 159629
rect 271045 159628 271111 159629
rect 275829 159628 275895 159629
rect 291009 159628 291075 159629
rect 256040 159626 256046 159628
rect 255958 159566 256046 159626
rect 256040 159564 256046 159566
rect 256110 159564 256116 159628
rect 271000 159626 271006 159628
rect 270954 159566 271006 159626
rect 271070 159624 271111 159628
rect 275760 159626 275766 159628
rect 271106 159568 271111 159624
rect 271000 159564 271006 159566
rect 271070 159564 271111 159568
rect 275738 159566 275766 159626
rect 275760 159564 275766 159566
rect 275830 159624 275895 159628
rect 290992 159626 290998 159628
rect 275830 159568 275834 159624
rect 275890 159568 275895 159624
rect 275830 159564 275895 159568
rect 290918 159566 290998 159626
rect 291062 159624 291075 159628
rect 291070 159568 291075 159624
rect 290992 159564 290998 159566
rect 291062 159564 291075 159568
rect 364558 159564 364564 159628
rect 364628 159626 364634 159628
rect 365253 159626 365319 159629
rect 364628 159624 365319 159626
rect 364628 159568 365258 159624
rect 365314 159568 365319 159624
rect 364628 159566 365319 159568
rect 364628 159564 364634 159566
rect 256049 159563 256115 159564
rect 271045 159563 271111 159564
rect 275829 159563 275895 159564
rect 291009 159563 291075 159564
rect 365253 159563 365319 159566
rect 262806 159292 262812 159356
rect 262876 159354 262882 159356
rect 367829 159354 367895 159357
rect 262876 159352 367895 159354
rect 262876 159296 367834 159352
rect 367890 159296 367895 159352
rect 262876 159294 367895 159296
rect 262876 159292 262882 159294
rect 367829 159291 367895 159294
rect 258206 159156 258212 159220
rect 258276 159218 258282 159220
rect 366357 159218 366423 159221
rect 258276 159216 366423 159218
rect 258276 159160 366362 159216
rect 366418 159160 366423 159216
rect 258276 159158 366423 159160
rect 258276 159156 258282 159158
rect 366357 159155 366423 159158
rect 255998 159020 256004 159084
rect 256068 159082 256074 159084
rect 366449 159082 366515 159085
rect 256068 159080 366515 159082
rect 256068 159024 366454 159080
rect 366510 159024 366515 159080
rect 256068 159022 366515 159024
rect 256068 159020 256074 159022
rect 366449 159019 366515 159022
rect 253606 158884 253612 158948
rect 253676 158946 253682 158948
rect 370681 158946 370747 158949
rect 253676 158944 370747 158946
rect 253676 158888 370686 158944
rect 370742 158888 370747 158944
rect 253676 158886 370747 158888
rect 253676 158884 253682 158886
rect 370681 158883 370747 158886
rect 243118 158748 243124 158812
rect 243188 158810 243194 158812
rect 357433 158810 357499 158813
rect 357566 158810 357572 158812
rect 243188 158750 357266 158810
rect 243188 158748 243194 158750
rect 214649 158674 214715 158677
rect 218973 158676 219039 158677
rect 214966 158674 214972 158676
rect 214649 158672 214972 158674
rect 214649 158616 214654 158672
rect 214710 158616 214972 158672
rect 214649 158614 214972 158616
rect 214649 158611 214715 158614
rect 214966 158612 214972 158614
rect 215036 158612 215042 158676
rect 218973 158672 219020 158676
rect 219084 158674 219090 158676
rect 227713 158674 227779 158677
rect 218973 158616 218978 158672
rect 218973 158612 219020 158616
rect 219084 158614 219130 158674
rect 219206 158672 227779 158674
rect 219206 158616 227718 158672
rect 227774 158616 227779 158672
rect 219206 158614 227779 158616
rect 219084 158612 219090 158614
rect 218973 158611 219039 158612
rect 218830 158476 218836 158540
rect 218900 158538 218906 158540
rect 219206 158538 219266 158614
rect 227713 158611 227779 158614
rect 238109 158676 238175 158677
rect 239581 158676 239647 158677
rect 238109 158672 238156 158676
rect 238220 158674 238226 158676
rect 238109 158616 238114 158672
rect 238109 158612 238156 158616
rect 238220 158614 238266 158674
rect 239581 158672 239628 158676
rect 239692 158674 239698 158676
rect 239581 158616 239586 158672
rect 238220 158612 238226 158614
rect 239581 158612 239628 158616
rect 239692 158614 239738 158674
rect 239692 158612 239698 158614
rect 241830 158612 241836 158676
rect 241900 158674 241906 158676
rect 242433 158674 242499 158677
rect 244273 158676 244339 158677
rect 248321 158676 248387 158677
rect 250897 158676 250963 158677
rect 244222 158674 244228 158676
rect 241900 158672 242499 158674
rect 241900 158616 242438 158672
rect 242494 158616 242499 158672
rect 241900 158614 242499 158616
rect 244182 158614 244228 158674
rect 244292 158672 244339 158676
rect 248270 158674 248276 158676
rect 244334 158616 244339 158672
rect 241900 158612 241906 158614
rect 238109 158611 238175 158612
rect 239581 158611 239647 158612
rect 242433 158611 242499 158614
rect 244222 158612 244228 158614
rect 244292 158612 244339 158616
rect 248230 158614 248276 158674
rect 248340 158672 248387 158676
rect 250846 158674 250852 158676
rect 248382 158616 248387 158672
rect 248270 158612 248276 158614
rect 248340 158612 248387 158616
rect 250806 158614 250852 158674
rect 250916 158672 250963 158676
rect 250958 158616 250963 158672
rect 250846 158612 250852 158614
rect 250916 158612 250963 158616
rect 251398 158612 251404 158676
rect 251468 158674 251474 158676
rect 252093 158674 252159 158677
rect 251468 158672 252159 158674
rect 251468 158616 252098 158672
rect 252154 158616 252159 158672
rect 251468 158614 252159 158616
rect 251468 158612 251474 158614
rect 244273 158611 244339 158612
rect 248321 158611 248387 158612
rect 250897 158611 250963 158612
rect 252093 158611 252159 158614
rect 257102 158612 257108 158676
rect 257172 158674 257178 158676
rect 257337 158674 257403 158677
rect 257172 158672 257403 158674
rect 257172 158616 257342 158672
rect 257398 158616 257403 158672
rect 257172 158614 257403 158616
rect 257172 158612 257178 158614
rect 257337 158611 257403 158614
rect 259494 158612 259500 158676
rect 259564 158674 259570 158676
rect 259913 158674 259979 158677
rect 261753 158676 261819 158677
rect 261702 158674 261708 158676
rect 259564 158672 259979 158674
rect 259564 158616 259918 158672
rect 259974 158616 259979 158672
rect 259564 158614 259979 158616
rect 261662 158614 261708 158674
rect 261772 158672 261819 158676
rect 261814 158616 261819 158672
rect 259564 158612 259570 158614
rect 259913 158611 259979 158614
rect 261702 158612 261708 158614
rect 261772 158612 261819 158616
rect 263910 158612 263916 158676
rect 263980 158674 263986 158676
rect 264329 158674 264395 158677
rect 263980 158672 264395 158674
rect 263980 158616 264334 158672
rect 264390 158616 264395 158672
rect 263980 158614 264395 158616
rect 263980 158612 263986 158614
rect 261753 158611 261819 158612
rect 264329 158611 264395 158614
rect 265382 158612 265388 158676
rect 265452 158674 265458 158676
rect 265893 158674 265959 158677
rect 268377 158676 268443 158677
rect 268745 158676 268811 158677
rect 269849 158676 269915 158677
rect 271137 158676 271203 158677
rect 272241 158676 272307 158677
rect 273345 158676 273411 158677
rect 274449 158676 274515 158677
rect 276105 158676 276171 158677
rect 281073 158676 281139 158677
rect 283649 158676 283715 158677
rect 293585 158676 293651 158677
rect 295977 158676 296043 158677
rect 298553 158676 298619 158677
rect 268326 158674 268332 158676
rect 265452 158672 265959 158674
rect 265452 158616 265898 158672
rect 265954 158616 265959 158672
rect 265452 158614 265959 158616
rect 268286 158614 268332 158674
rect 268396 158672 268443 158676
rect 268694 158674 268700 158676
rect 268438 158616 268443 158672
rect 265452 158612 265458 158614
rect 265893 158611 265959 158614
rect 268326 158612 268332 158614
rect 268396 158612 268443 158616
rect 268654 158614 268700 158674
rect 268764 158672 268811 158676
rect 269798 158674 269804 158676
rect 268806 158616 268811 158672
rect 268694 158612 268700 158614
rect 268764 158612 268811 158616
rect 269758 158614 269804 158674
rect 269868 158672 269915 158676
rect 271086 158674 271092 158676
rect 269910 158616 269915 158672
rect 269798 158612 269804 158614
rect 269868 158612 269915 158616
rect 271046 158614 271092 158674
rect 271156 158672 271203 158676
rect 272190 158674 272196 158676
rect 271198 158616 271203 158672
rect 271086 158612 271092 158614
rect 271156 158612 271203 158616
rect 272150 158614 272196 158674
rect 272260 158672 272307 158676
rect 273294 158674 273300 158676
rect 272302 158616 272307 158672
rect 272190 158612 272196 158614
rect 272260 158612 272307 158616
rect 273254 158614 273300 158674
rect 273364 158672 273411 158676
rect 274398 158674 274404 158676
rect 273406 158616 273411 158672
rect 273294 158612 273300 158614
rect 273364 158612 273411 158616
rect 274358 158614 274404 158674
rect 274468 158672 274515 158676
rect 276054 158674 276060 158676
rect 274510 158616 274515 158672
rect 274398 158612 274404 158614
rect 274468 158612 274515 158616
rect 276014 158614 276060 158674
rect 276124 158672 276171 158676
rect 281022 158674 281028 158676
rect 276166 158616 276171 158672
rect 276054 158612 276060 158614
rect 276124 158612 276171 158616
rect 280982 158614 281028 158674
rect 281092 158672 281139 158676
rect 283598 158674 283604 158676
rect 281134 158616 281139 158672
rect 281022 158612 281028 158614
rect 281092 158612 281139 158616
rect 283558 158614 283604 158674
rect 283668 158672 283715 158676
rect 293534 158674 293540 158676
rect 283710 158616 283715 158672
rect 283598 158612 283604 158614
rect 283668 158612 283715 158616
rect 293494 158614 293540 158674
rect 293604 158672 293651 158676
rect 295926 158674 295932 158676
rect 293646 158616 293651 158672
rect 293534 158612 293540 158614
rect 293604 158612 293651 158616
rect 295886 158614 295932 158674
rect 295996 158672 296043 158676
rect 298502 158674 298508 158676
rect 296038 158616 296043 158672
rect 295926 158612 295932 158614
rect 295996 158612 296043 158616
rect 298462 158614 298508 158674
rect 298572 158672 298619 158676
rect 298614 158616 298619 158672
rect 298502 158612 298508 158614
rect 298572 158612 298619 158616
rect 300894 158612 300900 158676
rect 300964 158674 300970 158676
rect 301037 158674 301103 158677
rect 303521 158676 303587 158677
rect 306097 158676 306163 158677
rect 308673 158676 308739 158677
rect 311065 158676 311131 158677
rect 313457 158676 313523 158677
rect 315849 158676 315915 158677
rect 318609 158676 318675 158677
rect 321001 158676 321067 158677
rect 323393 158676 323459 158677
rect 325969 158676 326035 158677
rect 303470 158674 303476 158676
rect 300964 158672 301103 158674
rect 300964 158616 301042 158672
rect 301098 158616 301103 158672
rect 300964 158614 301103 158616
rect 303430 158614 303476 158674
rect 303540 158672 303587 158676
rect 306046 158674 306052 158676
rect 303582 158616 303587 158672
rect 300964 158612 300970 158614
rect 268377 158611 268443 158612
rect 268745 158611 268811 158612
rect 269849 158611 269915 158612
rect 271137 158611 271203 158612
rect 272241 158611 272307 158612
rect 273345 158611 273411 158612
rect 274449 158611 274515 158612
rect 276105 158611 276171 158612
rect 281073 158611 281139 158612
rect 283649 158611 283715 158612
rect 293585 158611 293651 158612
rect 295977 158611 296043 158612
rect 298553 158611 298619 158612
rect 301037 158611 301103 158614
rect 303470 158612 303476 158614
rect 303540 158612 303587 158616
rect 306006 158614 306052 158674
rect 306116 158672 306163 158676
rect 308622 158674 308628 158676
rect 306158 158616 306163 158672
rect 306046 158612 306052 158614
rect 306116 158612 306163 158616
rect 308582 158614 308628 158674
rect 308692 158672 308739 158676
rect 311014 158674 311020 158676
rect 308734 158616 308739 158672
rect 308622 158612 308628 158614
rect 308692 158612 308739 158616
rect 310974 158614 311020 158674
rect 311084 158672 311131 158676
rect 313406 158674 313412 158676
rect 311126 158616 311131 158672
rect 311014 158612 311020 158614
rect 311084 158612 311131 158616
rect 313366 158614 313412 158674
rect 313476 158672 313523 158676
rect 315798 158674 315804 158676
rect 313518 158616 313523 158672
rect 313406 158612 313412 158614
rect 313476 158612 313523 158616
rect 315758 158614 315804 158674
rect 315868 158672 315915 158676
rect 318558 158674 318564 158676
rect 315910 158616 315915 158672
rect 315798 158612 315804 158614
rect 315868 158612 315915 158616
rect 318518 158614 318564 158674
rect 318628 158672 318675 158676
rect 320950 158674 320956 158676
rect 318670 158616 318675 158672
rect 318558 158612 318564 158614
rect 318628 158612 318675 158616
rect 320910 158614 320956 158674
rect 321020 158672 321067 158676
rect 323342 158674 323348 158676
rect 321062 158616 321067 158672
rect 320950 158612 320956 158614
rect 321020 158612 321067 158616
rect 323302 158614 323348 158674
rect 323412 158672 323459 158676
rect 325918 158674 325924 158676
rect 323454 158616 323459 158672
rect 323342 158612 323348 158614
rect 323412 158612 323459 158616
rect 325878 158614 325924 158674
rect 325988 158672 326035 158676
rect 326030 158616 326035 158672
rect 325918 158612 325924 158614
rect 325988 158612 326035 158616
rect 357206 158674 357266 158750
rect 357433 158808 357572 158810
rect 357433 158752 357438 158808
rect 357494 158752 357572 158808
rect 357433 158750 357572 158752
rect 357433 158747 357499 158750
rect 357566 158748 357572 158750
rect 357636 158748 357642 158812
rect 366541 158810 366607 158813
rect 357758 158750 364350 158810
rect 357758 158674 357818 158750
rect 357206 158614 357818 158674
rect 364290 158674 364350 158750
rect 364750 158808 366607 158810
rect 364750 158752 366546 158808
rect 366602 158752 366607 158808
rect 364750 158750 366607 158752
rect 364750 158674 364810 158750
rect 366541 158747 366607 158750
rect 364290 158614 364810 158674
rect 303521 158611 303587 158612
rect 306097 158611 306163 158612
rect 308673 158611 308739 158612
rect 311065 158611 311131 158612
rect 313457 158611 313523 158612
rect 315849 158611 315915 158612
rect 318609 158611 318675 158612
rect 321001 158611 321067 158612
rect 323393 158611 323459 158612
rect 325969 158611 326035 158612
rect 231853 158538 231919 158541
rect 218900 158478 219266 158538
rect 219390 158536 231919 158538
rect 219390 158480 231858 158536
rect 231914 158480 231919 158536
rect 219390 158478 231919 158480
rect 218900 158476 218906 158478
rect 217542 158340 217548 158404
rect 217612 158402 217618 158404
rect 219390 158402 219450 158478
rect 231853 158475 231919 158478
rect 237230 158476 237236 158540
rect 237300 158538 237306 158540
rect 363781 158538 363847 158541
rect 237300 158536 363847 158538
rect 237300 158480 363786 158536
rect 363842 158480 363847 158536
rect 237300 158478 363847 158480
rect 237300 158476 237306 158478
rect 363781 158475 363847 158478
rect 233233 158402 233299 158405
rect 240593 158404 240659 158405
rect 240542 158402 240548 158404
rect 217612 158342 219450 158402
rect 224174 158400 233299 158402
rect 224174 158344 233238 158400
rect 233294 158344 233299 158400
rect 224174 158342 233299 158344
rect 240502 158342 240548 158402
rect 240612 158400 240659 158404
rect 240654 158344 240659 158400
rect 217612 158340 217618 158342
rect 216254 158204 216260 158268
rect 216324 158266 216330 158268
rect 224174 158266 224234 158342
rect 233233 158339 233299 158342
rect 240542 158340 240548 158342
rect 240612 158340 240659 158344
rect 252318 158340 252324 158404
rect 252388 158402 252394 158404
rect 370405 158402 370471 158405
rect 252388 158400 370471 158402
rect 252388 158344 370410 158400
rect 370466 158344 370471 158400
rect 252388 158342 370471 158344
rect 252388 158340 252394 158342
rect 240593 158339 240659 158340
rect 370405 158339 370471 158342
rect 216324 158206 224234 158266
rect 224309 158266 224375 158269
rect 237373 158266 237439 158269
rect 249793 158266 249859 158269
rect 224309 158264 237439 158266
rect 224309 158208 224314 158264
rect 224370 158208 237378 158264
rect 237434 158208 237439 158264
rect 224309 158206 237439 158208
rect 216324 158204 216330 158206
rect 224309 158203 224375 158206
rect 237373 158203 237439 158206
rect 238710 158264 249859 158266
rect 238710 158208 249798 158264
rect 249854 158208 249859 158264
rect 238710 158206 249859 158208
rect 216070 158068 216076 158132
rect 216140 158130 216146 158132
rect 216213 158130 216279 158133
rect 216140 158128 216279 158130
rect 216140 158072 216218 158128
rect 216274 158072 216279 158128
rect 216140 158070 216279 158072
rect 216140 158068 216146 158070
rect 216213 158067 216279 158070
rect 217174 158068 217180 158132
rect 217244 158130 217250 158132
rect 238710 158130 238770 158206
rect 249793 158203 249859 158206
rect 258574 158204 258580 158268
rect 258644 158266 258650 158268
rect 373165 158266 373231 158269
rect 258644 158264 373231 158266
rect 258644 158208 373170 158264
rect 373226 158208 373231 158264
rect 258644 158206 373231 158208
rect 258644 158204 258650 158206
rect 373165 158203 373231 158206
rect 217244 158070 238770 158130
rect 217244 158068 217250 158070
rect 246614 158068 246620 158132
rect 246684 158130 246690 158132
rect 246757 158130 246823 158133
rect 246684 158128 246823 158130
rect 246684 158072 246762 158128
rect 246818 158072 246823 158128
rect 246684 158070 246823 158072
rect 246684 158068 246690 158070
rect 246757 158067 246823 158070
rect 254526 158068 254532 158132
rect 254596 158130 254602 158132
rect 366265 158130 366331 158133
rect 254596 158128 366331 158130
rect 254596 158072 366270 158128
rect 366326 158072 366331 158128
rect 254596 158070 366331 158072
rect 254596 158068 254602 158070
rect 366265 158067 366331 158070
rect 216990 157932 216996 157996
rect 217060 157994 217066 157996
rect 251173 157994 251239 157997
rect 217060 157992 251239 157994
rect 217060 157936 251178 157992
rect 251234 157936 251239 157992
rect 217060 157934 251239 157936
rect 217060 157932 217066 157934
rect 251173 157931 251239 157934
rect 260782 157932 260788 157996
rect 260852 157994 260858 157996
rect 369209 157994 369275 157997
rect 260852 157992 369275 157994
rect 260852 157936 369214 157992
rect 369270 157936 369275 157992
rect 260852 157934 369275 157936
rect 260852 157932 260858 157934
rect 369209 157931 369275 157934
rect 217358 157796 217364 157860
rect 217428 157858 217434 157860
rect 224953 157858 225019 157861
rect 245561 157860 245627 157861
rect 247769 157860 247835 157861
rect 248689 157860 248755 157861
rect 245510 157858 245516 157860
rect 217428 157856 225019 157858
rect 217428 157800 224958 157856
rect 225014 157800 225019 157856
rect 217428 157798 225019 157800
rect 245470 157798 245516 157858
rect 245580 157856 245627 157860
rect 247718 157858 247724 157860
rect 245622 157800 245627 157856
rect 217428 157796 217434 157798
rect 224953 157795 225019 157798
rect 245510 157796 245516 157798
rect 245580 157796 245627 157800
rect 247678 157798 247724 157858
rect 247788 157856 247835 157860
rect 248638 157858 248644 157860
rect 247830 157800 247835 157856
rect 247718 157796 247724 157798
rect 247788 157796 247835 157800
rect 248598 157798 248644 157858
rect 248708 157856 248755 157860
rect 248750 157800 248755 157856
rect 248638 157796 248644 157798
rect 248708 157796 248755 157800
rect 250110 157796 250116 157860
rect 250180 157858 250186 157860
rect 250713 157858 250779 157861
rect 253473 157860 253539 157861
rect 253422 157858 253428 157860
rect 250180 157856 250779 157858
rect 250180 157800 250718 157856
rect 250774 157800 250779 157856
rect 250180 157798 250779 157800
rect 253382 157798 253428 157858
rect 253492 157856 253539 157860
rect 253534 157800 253539 157856
rect 250180 157796 250186 157798
rect 245561 157795 245627 157796
rect 247769 157795 247835 157796
rect 248689 157795 248755 157796
rect 250713 157795 250779 157798
rect 253422 157796 253428 157798
rect 253492 157796 253539 157800
rect 267038 157796 267044 157860
rect 267108 157858 267114 157860
rect 355501 157858 355567 157861
rect 267108 157856 355567 157858
rect 267108 157800 355506 157856
rect 355562 157800 355567 157856
rect 267108 157798 355567 157800
rect 267108 157796 267114 157798
rect 253473 157795 253539 157796
rect 355501 157795 355567 157798
rect 212942 157660 212948 157724
rect 213012 157722 213018 157724
rect 224309 157722 224375 157725
rect 213012 157720 224375 157722
rect 213012 157664 224314 157720
rect 224370 157664 224375 157720
rect 213012 157662 224375 157664
rect 213012 157660 213018 157662
rect 224309 157659 224375 157662
rect 266486 157660 266492 157724
rect 266556 157722 266562 157724
rect 266629 157722 266695 157725
rect 273713 157724 273779 157725
rect 278497 157724 278563 157725
rect 273662 157722 273668 157724
rect 266556 157720 266695 157722
rect 266556 157664 266634 157720
rect 266690 157664 266695 157720
rect 266556 157662 266695 157664
rect 273622 157662 273668 157722
rect 273732 157720 273779 157724
rect 278446 157722 278452 157724
rect 273774 157664 273779 157720
rect 266556 157660 266562 157662
rect 266629 157659 266695 157662
rect 273662 157660 273668 157662
rect 273732 157660 273779 157664
rect 278406 157662 278452 157722
rect 278516 157720 278563 157724
rect 278558 157664 278563 157720
rect 278446 157660 278452 157662
rect 278516 157660 278563 157664
rect 273713 157659 273779 157660
rect 278497 157659 278563 157660
rect 261201 157588 261267 157589
rect 261150 157586 261156 157588
rect 261110 157526 261156 157586
rect 261220 157584 261267 157588
rect 261262 157528 261267 157584
rect 261150 157524 261156 157526
rect 261220 157524 261267 157528
rect 263542 157524 263548 157588
rect 263612 157586 263618 157588
rect 263685 157586 263751 157589
rect 265985 157588 266051 157589
rect 288249 157588 288315 157589
rect 265934 157586 265940 157588
rect 263612 157584 263751 157586
rect 263612 157528 263690 157584
rect 263746 157528 263751 157584
rect 263612 157526 263751 157528
rect 265894 157526 265940 157586
rect 266004 157584 266051 157588
rect 288198 157586 288204 157588
rect 266046 157528 266051 157584
rect 263612 157524 263618 157526
rect 261201 157523 261267 157524
rect 263685 157523 263751 157526
rect 265934 157524 265940 157526
rect 266004 157524 266051 157528
rect 288158 157526 288204 157586
rect 288268 157584 288315 157588
rect 288310 157528 288315 157584
rect 288198 157524 288204 157526
rect 288268 157524 288315 157528
rect 265985 157523 266051 157524
rect 288249 157523 288315 157524
rect 236494 157388 236500 157452
rect 236564 157450 236570 157452
rect 363689 157450 363755 157453
rect 236564 157448 363755 157450
rect 236564 157392 363694 157448
rect 363750 157392 363755 157448
rect 236564 157390 363755 157392
rect 236564 157388 236570 157390
rect 363689 157387 363755 157390
rect 217961 155954 218027 155957
rect 264973 155954 265039 155957
rect 217961 155952 265039 155954
rect 217961 155896 217966 155952
rect 218022 155896 264978 155952
rect 265034 155896 265039 155952
rect 217961 155894 265039 155896
rect 217961 155891 218027 155894
rect 264973 155891 265039 155894
rect 213361 155818 213427 155821
rect 260833 155818 260899 155821
rect 213361 155816 260899 155818
rect 213361 155760 213366 155816
rect 213422 155760 260838 155816
rect 260894 155760 260899 155816
rect 213361 155758 260899 155760
rect 213361 155755 213427 155758
rect 260833 155755 260899 155758
rect 216029 155682 216095 155685
rect 263593 155682 263659 155685
rect 216029 155680 263659 155682
rect 216029 155624 216034 155680
rect 216090 155624 263598 155680
rect 263654 155624 263659 155680
rect 216029 155622 263659 155624
rect 216029 155619 216095 155622
rect 263593 155619 263659 155622
rect 213269 155546 213335 155549
rect 267733 155546 267799 155549
rect 213269 155544 267799 155546
rect 213269 155488 213274 155544
rect 213330 155488 267738 155544
rect 267794 155488 267799 155544
rect 213269 155486 267799 155488
rect 213269 155483 213335 155486
rect 267733 155483 267799 155486
rect 217777 155410 217843 155413
rect 274633 155410 274699 155413
rect 217777 155408 274699 155410
rect 217777 155352 217782 155408
rect 217838 155352 274638 155408
rect 274694 155352 274699 155408
rect 217777 155350 274699 155352
rect 217777 155347 217843 155350
rect 274633 155347 274699 155350
rect 210969 155274 211035 155277
rect 267825 155274 267891 155277
rect 210969 155272 267891 155274
rect 210969 155216 210974 155272
rect 211030 155216 267830 155272
rect 267886 155216 267891 155272
rect 210969 155214 267891 155216
rect 210969 155211 211035 155214
rect 267825 155211 267891 155214
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580349 112842 580415 112845
rect 583520 112842 584960 112932
rect 580349 112840 584960 112842
rect 580349 112784 580354 112840
rect 580410 112784 584960 112840
rect 580349 112782 584960 112784
rect 580349 112779 580415 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 363454 71844 363460 71908
rect 363524 71906 363530 71908
rect 583526 71906 583586 72798
rect 363524 71846 583586 71906
rect 363524 71844 363530 71846
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 360326 44298 360332 44300
rect 6870 44238 360332 44298
rect 360326 44236 360332 44238
rect 360396 44236 360402 44300
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 319713 8938 319779 8941
rect 365989 8938 366055 8941
rect 319713 8936 366055 8938
rect 319713 8880 319718 8936
rect 319774 8880 365994 8936
rect 366050 8880 366055 8936
rect 319713 8878 366055 8880
rect 319713 8875 319779 8878
rect 365989 8875 366055 8878
rect 350441 6762 350507 6765
rect 363321 6762 363387 6765
rect 350441 6760 363387 6762
rect 350441 6704 350446 6760
rect 350502 6704 363326 6760
rect 363382 6704 363387 6760
rect 350441 6702 363387 6704
rect 350441 6699 350507 6702
rect 363321 6699 363387 6702
rect 348049 6626 348115 6629
rect 367185 6626 367251 6629
rect 348049 6624 367251 6626
rect -960 6490 480 6580
rect 348049 6568 348054 6624
rect 348110 6568 367190 6624
rect 367246 6568 367251 6624
rect 348049 6566 367251 6568
rect 348049 6563 348115 6566
rect 367185 6563 367251 6566
rect 344553 6490 344619 6493
rect 367093 6490 367159 6493
rect -960 6430 674 6490
rect -960 6354 480 6430
rect 614 6354 674 6430
rect 344553 6488 367159 6490
rect 344553 6432 344558 6488
rect 344614 6432 367098 6488
rect 367154 6432 367159 6488
rect 583520 6476 584960 6716
rect 344553 6430 367159 6432
rect 344553 6427 344619 6430
rect 367093 6427 367159 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 340965 6354 341031 6357
rect 364701 6354 364767 6357
rect 340965 6352 364767 6354
rect 340965 6296 340970 6352
rect 341026 6296 364706 6352
rect 364762 6296 364767 6352
rect 340965 6294 364767 6296
rect 246 5810 306 6294
rect 340965 6291 341031 6294
rect 364701 6291 364767 6294
rect 337469 6218 337535 6221
rect 363229 6218 363295 6221
rect 337469 6216 363295 6218
rect 337469 6160 337474 6216
rect 337530 6160 363234 6216
rect 363290 6160 363295 6216
rect 337469 6158 363295 6160
rect 337469 6155 337535 6158
rect 363229 6155 363295 6158
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 361614 5674 361620 5676
rect 6870 5614 361620 5674
rect 361614 5612 361620 5614
rect 361684 5612 361690 5676
rect 368974 4796 368980 4860
rect 369044 4858 369050 4860
rect 582189 4858 582255 4861
rect 369044 4856 582255 4858
rect 369044 4800 582194 4856
rect 582250 4800 582255 4856
rect 369044 4798 582255 4800
rect 369044 4796 369050 4798
rect 582189 4795 582255 4798
rect 214925 4042 214991 4045
rect 218789 4042 218855 4045
rect 214925 4040 218855 4042
rect 214925 3984 214930 4040
rect 214986 3984 218794 4040
rect 218850 3984 218855 4040
rect 214925 3982 218855 3984
rect 214925 3979 214991 3982
rect 218789 3979 218855 3982
rect 345749 4042 345815 4045
rect 360510 4042 360516 4044
rect 345749 4040 360516 4042
rect 345749 3984 345754 4040
rect 345810 3984 360516 4040
rect 345749 3982 360516 3984
rect 345749 3979 345815 3982
rect 360510 3980 360516 3982
rect 360580 3980 360586 4044
rect 367318 4042 367324 4044
rect 364290 3982 367324 4042
rect 215017 3906 215083 3909
rect 222745 3906 222811 3909
rect 215017 3904 222811 3906
rect 215017 3848 215022 3904
rect 215078 3848 222750 3904
rect 222806 3848 222811 3904
rect 215017 3846 222811 3848
rect 215017 3843 215083 3846
rect 222745 3843 222811 3846
rect 351637 3906 351703 3909
rect 364290 3906 364350 3982
rect 367318 3980 367324 3982
rect 367388 3980 367394 4044
rect 351637 3904 364350 3906
rect 351637 3848 351642 3904
rect 351698 3848 364350 3904
rect 351637 3846 364350 3848
rect 351637 3843 351703 3846
rect 364926 3844 364932 3908
rect 364996 3906 365002 3908
rect 379973 3906 380039 3909
rect 364996 3904 380039 3906
rect 364996 3848 379978 3904
rect 380034 3848 380039 3904
rect 364996 3846 380039 3848
rect 364996 3844 365002 3846
rect 379973 3843 380039 3846
rect 215109 3770 215175 3773
rect 227529 3770 227595 3773
rect 215109 3768 227595 3770
rect 215109 3712 215114 3768
rect 215170 3712 227534 3768
rect 227590 3712 227595 3768
rect 215109 3710 227595 3712
rect 215109 3707 215175 3710
rect 227529 3707 227595 3710
rect 338665 3770 338731 3773
rect 356237 3770 356303 3773
rect 358486 3770 358492 3772
rect 338665 3768 356303 3770
rect 338665 3712 338670 3768
rect 338726 3712 356242 3768
rect 356298 3712 356303 3768
rect 338665 3710 356303 3712
rect 338665 3707 338731 3710
rect 356237 3707 356303 3710
rect 356470 3710 358492 3770
rect 216857 3634 216923 3637
rect 218646 3634 218652 3636
rect 216857 3632 218652 3634
rect 216857 3576 216862 3632
rect 216918 3576 218652 3632
rect 216857 3574 218652 3576
rect 216857 3571 216923 3574
rect 218646 3572 218652 3574
rect 218716 3572 218722 3636
rect 218789 3634 218855 3637
rect 226333 3634 226399 3637
rect 218789 3632 226399 3634
rect 218789 3576 218794 3632
rect 218850 3576 226338 3632
rect 226394 3576 226399 3632
rect 218789 3574 226399 3576
rect 218789 3571 218855 3574
rect 226333 3571 226399 3574
rect 335077 3634 335143 3637
rect 356470 3634 356530 3710
rect 358486 3708 358492 3710
rect 358556 3708 358562 3772
rect 367686 3708 367692 3772
rect 367756 3770 367762 3772
rect 367756 3710 370882 3770
rect 367756 3708 367762 3710
rect 335077 3632 356530 3634
rect 335077 3576 335082 3632
rect 335138 3576 356530 3632
rect 335077 3574 356530 3576
rect 335077 3571 335143 3574
rect 358118 3572 358124 3636
rect 358188 3634 358194 3636
rect 358721 3634 358787 3637
rect 358188 3632 358787 3634
rect 358188 3576 358726 3632
rect 358782 3576 358787 3632
rect 358188 3574 358787 3576
rect 358188 3572 358194 3574
rect 358721 3571 358787 3574
rect 364374 3572 364380 3636
rect 364444 3634 364450 3636
rect 364609 3634 364675 3637
rect 364444 3632 364675 3634
rect 364444 3576 364614 3632
rect 364670 3576 364675 3632
rect 364444 3574 364675 3576
rect 364444 3572 364450 3574
rect 364609 3571 364675 3574
rect 365662 3572 365668 3636
rect 365732 3634 365738 3636
rect 365805 3634 365871 3637
rect 365732 3632 365871 3634
rect 365732 3576 365810 3632
rect 365866 3576 365871 3632
rect 365732 3574 365871 3576
rect 365732 3572 365738 3574
rect 365805 3571 365871 3574
rect 367134 3572 367140 3636
rect 367204 3634 367210 3636
rect 368197 3634 368263 3637
rect 367204 3632 368263 3634
rect 367204 3576 368202 3632
rect 368258 3576 368263 3632
rect 367204 3574 368263 3576
rect 367204 3572 367210 3574
rect 368197 3571 368263 3574
rect 368422 3572 368428 3636
rect 368492 3634 368498 3636
rect 369393 3634 369459 3637
rect 368492 3632 369459 3634
rect 368492 3576 369398 3632
rect 369454 3576 369459 3632
rect 368492 3574 369459 3576
rect 368492 3572 368498 3574
rect 369393 3571 369459 3574
rect 369894 3572 369900 3636
rect 369964 3634 369970 3636
rect 370589 3634 370655 3637
rect 369964 3632 370655 3634
rect 369964 3576 370594 3632
rect 370650 3576 370655 3632
rect 369964 3574 370655 3576
rect 370822 3634 370882 3710
rect 394233 3634 394299 3637
rect 370822 3632 394299 3634
rect 370822 3576 394238 3632
rect 394294 3576 394299 3632
rect 370822 3574 394299 3576
rect 369964 3572 369970 3574
rect 370589 3571 370655 3574
rect 394233 3571 394299 3574
rect 213126 3436 213132 3500
rect 213196 3498 213202 3500
rect 213361 3498 213427 3501
rect 213196 3496 213427 3498
rect 213196 3440 213366 3496
rect 213422 3440 213427 3496
rect 213196 3438 213427 3440
rect 213196 3436 213202 3438
rect 213361 3435 213427 3438
rect 214465 3498 214531 3501
rect 215150 3498 215156 3500
rect 214465 3496 215156 3498
rect 214465 3440 214470 3496
rect 214526 3440 215156 3496
rect 214465 3438 215156 3440
rect 214465 3435 214531 3438
rect 215150 3436 215156 3438
rect 215220 3436 215226 3500
rect 215661 3498 215727 3501
rect 216438 3498 216444 3500
rect 215661 3496 216444 3498
rect 215661 3440 215666 3496
rect 215722 3440 216444 3496
rect 215661 3438 216444 3440
rect 215661 3435 215727 3438
rect 216438 3436 216444 3438
rect 216508 3436 216514 3500
rect 218053 3498 218119 3501
rect 219198 3498 219204 3500
rect 218053 3496 219204 3498
rect 218053 3440 218058 3496
rect 218114 3440 219204 3496
rect 218053 3438 219204 3440
rect 218053 3435 218119 3438
rect 219198 3436 219204 3438
rect 219268 3436 219274 3500
rect 219341 3498 219407 3501
rect 237005 3498 237071 3501
rect 219341 3496 237071 3498
rect 219341 3440 219346 3496
rect 219402 3440 237010 3496
rect 237066 3440 237071 3496
rect 219341 3438 237071 3440
rect 219341 3435 219407 3438
rect 237005 3435 237071 3438
rect 331581 3498 331647 3501
rect 357525 3498 357591 3501
rect 358302 3498 358308 3500
rect 331581 3496 357082 3498
rect 331581 3440 331586 3496
rect 331642 3440 357082 3496
rect 331581 3438 357082 3440
rect 331581 3435 331647 3438
rect 208577 3362 208643 3365
rect 214414 3362 214420 3364
rect 208577 3360 214420 3362
rect 208577 3304 208582 3360
rect 208638 3304 214420 3360
rect 208577 3302 214420 3304
rect 208577 3299 208643 3302
rect 214414 3300 214420 3302
rect 214484 3300 214490 3364
rect 216581 3362 216647 3365
rect 240501 3362 240567 3365
rect 216581 3360 240567 3362
rect 216581 3304 216586 3360
rect 216642 3304 240506 3360
rect 240562 3304 240567 3360
rect 216581 3302 240567 3304
rect 216581 3299 216647 3302
rect 240501 3299 240567 3302
rect 327993 3362 328059 3365
rect 357022 3362 357082 3438
rect 357525 3496 358308 3498
rect 357525 3440 357530 3496
rect 357586 3440 358308 3496
rect 357525 3438 358308 3440
rect 357525 3435 357591 3438
rect 358302 3436 358308 3438
rect 358372 3436 358378 3500
rect 358854 3436 358860 3500
rect 358924 3498 358930 3500
rect 359917 3498 359983 3501
rect 358924 3496 359983 3498
rect 358924 3440 359922 3496
rect 359978 3440 359983 3496
rect 358924 3438 359983 3440
rect 358924 3436 358930 3438
rect 359917 3435 359983 3438
rect 360142 3436 360148 3500
rect 360212 3498 360218 3500
rect 361113 3498 361179 3501
rect 360212 3496 361179 3498
rect 360212 3440 361118 3496
rect 361174 3440 361179 3496
rect 360212 3438 361179 3440
rect 360212 3436 360218 3438
rect 361113 3435 361179 3438
rect 362309 3498 362375 3501
rect 362534 3498 362540 3500
rect 362309 3496 362540 3498
rect 362309 3440 362314 3496
rect 362370 3440 362540 3496
rect 362309 3438 362540 3440
rect 362309 3435 362375 3438
rect 362534 3436 362540 3438
rect 362604 3436 362610 3500
rect 362902 3436 362908 3500
rect 362972 3498 362978 3500
rect 363505 3498 363571 3501
rect 362972 3496 363571 3498
rect 362972 3440 363510 3496
rect 363566 3440 363571 3496
rect 362972 3438 363571 3440
rect 362972 3436 362978 3438
rect 363505 3435 363571 3438
rect 363638 3436 363644 3500
rect 363708 3498 363714 3500
rect 390645 3498 390711 3501
rect 363708 3496 390711 3498
rect 363708 3440 390650 3496
rect 390706 3440 390711 3496
rect 363708 3438 390711 3440
rect 363708 3436 363714 3438
rect 390645 3435 390711 3438
rect 359406 3362 359412 3364
rect 327993 3360 356162 3362
rect 327993 3304 327998 3360
rect 328054 3304 356162 3360
rect 327993 3302 356162 3304
rect 357022 3302 359412 3362
rect 327993 3299 328059 3302
rect 214833 3226 214899 3229
rect 219341 3226 219407 3229
rect 214833 3224 219407 3226
rect 214833 3168 214838 3224
rect 214894 3168 219346 3224
rect 219402 3168 219407 3224
rect 214833 3166 219407 3168
rect 214833 3163 214899 3166
rect 219341 3163 219407 3166
rect 349245 3226 349311 3229
rect 349245 3224 354690 3226
rect 349245 3168 349250 3224
rect 349306 3168 354690 3224
rect 349245 3166 354690 3168
rect 349245 3163 349311 3166
rect 354630 2954 354690 3166
rect 356102 3090 356162 3302
rect 359406 3300 359412 3302
rect 359476 3300 359482 3364
rect 369158 3300 369164 3364
rect 369228 3362 369234 3364
rect 397729 3362 397795 3365
rect 369228 3360 397795 3362
rect 369228 3304 397734 3360
rect 397790 3304 397795 3360
rect 369228 3302 397795 3304
rect 369228 3300 369234 3302
rect 397729 3299 397795 3302
rect 356237 3226 356303 3229
rect 360694 3226 360700 3228
rect 356237 3224 360700 3226
rect 356237 3168 356242 3224
rect 356298 3168 360700 3224
rect 356237 3166 360700 3168
rect 356237 3163 356303 3166
rect 360694 3164 360700 3166
rect 360764 3164 360770 3228
rect 359222 3090 359228 3092
rect 356102 3030 359228 3090
rect 359222 3028 359228 3030
rect 359292 3028 359298 3092
rect 359038 2954 359044 2956
rect 354630 2894 359044 2954
rect 359038 2892 359044 2894
rect 359108 2892 359114 2956
<< via3 >>
rect 278452 476988 278516 477052
rect 305868 476988 305932 477052
rect 308444 476988 308508 477052
rect 253428 476852 253492 476916
rect 255820 476852 255884 476916
rect 270908 476852 270972 476916
rect 311020 476852 311084 476916
rect 323348 476852 323412 476916
rect 256188 476716 256252 476780
rect 303476 476716 303540 476780
rect 248276 476580 248340 476644
rect 250668 476580 250732 476644
rect 253612 476580 253676 476644
rect 263548 476640 263612 476644
rect 263548 476584 263598 476640
rect 263598 476584 263612 476640
rect 263548 476580 263612 476584
rect 265940 476580 266004 476644
rect 272196 476580 272260 476644
rect 244228 476504 244292 476508
rect 244228 476448 244278 476504
rect 244278 476448 244292 476504
rect 244228 476444 244292 476448
rect 260604 476444 260668 476508
rect 268332 476444 268396 476508
rect 273484 476444 273548 476508
rect 313412 476444 313476 476508
rect 315804 476444 315868 476508
rect 238156 476308 238220 476372
rect 243124 476308 243188 476372
rect 245332 476308 245396 476372
rect 251404 476308 251468 476372
rect 257108 476308 257172 476372
rect 258396 476308 258460 476372
rect 260972 476308 261036 476372
rect 266492 476308 266556 476372
rect 273300 476308 273364 476372
rect 276060 476368 276124 476372
rect 276060 476312 276074 476368
rect 276074 476312 276124 476368
rect 276060 476308 276124 476312
rect 280844 476308 280908 476372
rect 318380 476308 318444 476372
rect 320956 476308 321020 476372
rect 235948 476232 236012 476236
rect 235948 476176 235962 476232
rect 235962 476176 236012 476232
rect 235948 476172 236012 476176
rect 237236 476172 237300 476236
rect 239628 476172 239692 476236
rect 240548 476172 240612 476236
rect 241836 476172 241900 476236
rect 246436 476172 246500 476236
rect 247540 476172 247604 476236
rect 248644 476172 248708 476236
rect 250116 476172 250180 476236
rect 252324 476172 252388 476236
rect 254532 476172 254596 476236
rect 258028 476172 258092 476236
rect 259500 476172 259564 476236
rect 261708 476172 261772 476236
rect 262812 476172 262876 476236
rect 263916 476172 263980 476236
rect 265388 476172 265452 476236
rect 267596 476232 267660 476236
rect 267596 476176 267610 476232
rect 267610 476176 267660 476232
rect 267596 476172 267660 476176
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 274404 476232 274468 476236
rect 274404 476176 274454 476232
rect 274454 476176 274468 476232
rect 274404 476172 274468 476176
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278084 476172 278148 476236
rect 279188 476172 279252 476236
rect 283420 476172 283484 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293356 476172 293420 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476232 300964 476236
rect 300900 476176 300914 476232
rect 300914 476176 300964 476232
rect 300900 476172 300964 476176
rect 325924 476172 325988 476236
rect 368980 444484 369044 444548
rect 363460 443260 363524 443324
rect 214604 443124 214668 443188
rect 215892 442988 215956 443052
rect 360332 442172 360396 442236
rect 361620 442172 361684 442236
rect 363828 441628 363892 441692
rect 219020 308892 219084 308956
rect 218836 308756 218900 308820
rect 217364 308620 217428 308684
rect 217548 308484 217612 308548
rect 216076 306172 216140 306236
rect 214972 306036 215036 306100
rect 216260 305900 216324 305964
rect 216996 305764 217060 305828
rect 217180 305628 217244 305692
rect 369164 304132 369228 304196
rect 363644 303180 363708 303244
rect 212948 303044 213012 303108
rect 367692 303044 367756 303108
rect 364932 301412 364996 301476
rect 368428 297332 368492 297396
rect 367140 283460 367204 283524
rect 364380 282100 364444 282164
rect 216444 275164 216508 275228
rect 214420 273804 214484 273868
rect 369900 269724 369964 269788
rect 215156 267004 215220 267068
rect 362908 265508 362972 265572
rect 358860 264148 358924 264212
rect 219204 262788 219268 262852
rect 362540 254628 362604 254692
rect 365668 254492 365732 254556
rect 367324 250820 367388 250884
rect 213132 249052 213196 249116
rect 364564 248100 364628 248164
rect 360148 246196 360212 246260
rect 358124 245516 358188 245580
rect 358308 245380 358372 245444
rect 358492 245244 358556 245308
rect 359044 245108 359108 245172
rect 359228 244972 359292 245036
rect 359412 244836 359476 244900
rect 357572 244700 357636 244764
rect 360516 244564 360580 244628
rect 360700 244428 360764 244492
rect 218652 243476 218716 243540
rect 214604 213964 214668 214028
rect 363828 191796 363892 191860
rect 215892 162828 215956 162892
rect 276990 159896 277054 159900
rect 276990 159840 277030 159896
rect 277030 159840 277054 159896
rect 276990 159836 277054 159840
rect 278078 159896 278142 159900
rect 278078 159840 278134 159896
rect 278134 159840 278142 159896
rect 278078 159836 278142 159840
rect 279166 159836 279230 159900
rect 285966 159896 286030 159900
rect 285966 159840 286010 159896
rect 286010 159840 286030 159896
rect 285966 159836 286030 159840
rect 256046 159624 256110 159628
rect 256046 159568 256054 159624
rect 256054 159568 256110 159624
rect 256046 159564 256110 159568
rect 271006 159624 271070 159628
rect 271006 159568 271050 159624
rect 271050 159568 271070 159624
rect 271006 159564 271070 159568
rect 275766 159564 275830 159628
rect 290998 159624 291062 159628
rect 290998 159568 291014 159624
rect 291014 159568 291062 159624
rect 290998 159564 291062 159568
rect 364564 159564 364628 159628
rect 262812 159292 262876 159356
rect 258212 159156 258276 159220
rect 256004 159020 256068 159084
rect 253612 158884 253676 158948
rect 243124 158748 243188 158812
rect 214972 158612 215036 158676
rect 219020 158672 219084 158676
rect 219020 158616 219034 158672
rect 219034 158616 219084 158672
rect 219020 158612 219084 158616
rect 218836 158476 218900 158540
rect 238156 158672 238220 158676
rect 238156 158616 238170 158672
rect 238170 158616 238220 158672
rect 238156 158612 238220 158616
rect 239628 158672 239692 158676
rect 239628 158616 239642 158672
rect 239642 158616 239692 158672
rect 239628 158612 239692 158616
rect 241836 158612 241900 158676
rect 244228 158672 244292 158676
rect 244228 158616 244278 158672
rect 244278 158616 244292 158672
rect 244228 158612 244292 158616
rect 248276 158672 248340 158676
rect 248276 158616 248326 158672
rect 248326 158616 248340 158672
rect 248276 158612 248340 158616
rect 250852 158672 250916 158676
rect 250852 158616 250902 158672
rect 250902 158616 250916 158672
rect 250852 158612 250916 158616
rect 251404 158612 251468 158676
rect 257108 158612 257172 158676
rect 259500 158612 259564 158676
rect 261708 158672 261772 158676
rect 261708 158616 261758 158672
rect 261758 158616 261772 158672
rect 261708 158612 261772 158616
rect 263916 158612 263980 158676
rect 265388 158612 265452 158676
rect 268332 158672 268396 158676
rect 268332 158616 268382 158672
rect 268382 158616 268396 158672
rect 268332 158612 268396 158616
rect 268700 158672 268764 158676
rect 268700 158616 268750 158672
rect 268750 158616 268764 158672
rect 268700 158612 268764 158616
rect 269804 158672 269868 158676
rect 269804 158616 269854 158672
rect 269854 158616 269868 158672
rect 269804 158612 269868 158616
rect 271092 158672 271156 158676
rect 271092 158616 271142 158672
rect 271142 158616 271156 158672
rect 271092 158612 271156 158616
rect 272196 158672 272260 158676
rect 272196 158616 272246 158672
rect 272246 158616 272260 158672
rect 272196 158612 272260 158616
rect 273300 158672 273364 158676
rect 273300 158616 273350 158672
rect 273350 158616 273364 158672
rect 273300 158612 273364 158616
rect 274404 158672 274468 158676
rect 274404 158616 274454 158672
rect 274454 158616 274468 158672
rect 274404 158612 274468 158616
rect 276060 158672 276124 158676
rect 276060 158616 276110 158672
rect 276110 158616 276124 158672
rect 276060 158612 276124 158616
rect 281028 158672 281092 158676
rect 281028 158616 281078 158672
rect 281078 158616 281092 158672
rect 281028 158612 281092 158616
rect 283604 158672 283668 158676
rect 283604 158616 283654 158672
rect 283654 158616 283668 158672
rect 283604 158612 283668 158616
rect 293540 158672 293604 158676
rect 293540 158616 293590 158672
rect 293590 158616 293604 158672
rect 293540 158612 293604 158616
rect 295932 158672 295996 158676
rect 295932 158616 295982 158672
rect 295982 158616 295996 158672
rect 295932 158612 295996 158616
rect 298508 158672 298572 158676
rect 298508 158616 298558 158672
rect 298558 158616 298572 158672
rect 298508 158612 298572 158616
rect 300900 158612 300964 158676
rect 303476 158672 303540 158676
rect 303476 158616 303526 158672
rect 303526 158616 303540 158672
rect 303476 158612 303540 158616
rect 306052 158672 306116 158676
rect 306052 158616 306102 158672
rect 306102 158616 306116 158672
rect 306052 158612 306116 158616
rect 308628 158672 308692 158676
rect 308628 158616 308678 158672
rect 308678 158616 308692 158672
rect 308628 158612 308692 158616
rect 311020 158672 311084 158676
rect 311020 158616 311070 158672
rect 311070 158616 311084 158672
rect 311020 158612 311084 158616
rect 313412 158672 313476 158676
rect 313412 158616 313462 158672
rect 313462 158616 313476 158672
rect 313412 158612 313476 158616
rect 315804 158672 315868 158676
rect 315804 158616 315854 158672
rect 315854 158616 315868 158672
rect 315804 158612 315868 158616
rect 318564 158672 318628 158676
rect 318564 158616 318614 158672
rect 318614 158616 318628 158672
rect 318564 158612 318628 158616
rect 320956 158672 321020 158676
rect 320956 158616 321006 158672
rect 321006 158616 321020 158672
rect 320956 158612 321020 158616
rect 323348 158672 323412 158676
rect 323348 158616 323398 158672
rect 323398 158616 323412 158672
rect 323348 158612 323412 158616
rect 325924 158672 325988 158676
rect 325924 158616 325974 158672
rect 325974 158616 325988 158672
rect 325924 158612 325988 158616
rect 357572 158748 357636 158812
rect 217548 158340 217612 158404
rect 237236 158476 237300 158540
rect 240548 158400 240612 158404
rect 240548 158344 240598 158400
rect 240598 158344 240612 158400
rect 216260 158204 216324 158268
rect 240548 158340 240612 158344
rect 252324 158340 252388 158404
rect 216076 158068 216140 158132
rect 217180 158068 217244 158132
rect 258580 158204 258644 158268
rect 246620 158068 246684 158132
rect 254532 158068 254596 158132
rect 216996 157932 217060 157996
rect 260788 157932 260852 157996
rect 217364 157796 217428 157860
rect 245516 157856 245580 157860
rect 245516 157800 245566 157856
rect 245566 157800 245580 157856
rect 245516 157796 245580 157800
rect 247724 157856 247788 157860
rect 247724 157800 247774 157856
rect 247774 157800 247788 157856
rect 247724 157796 247788 157800
rect 248644 157856 248708 157860
rect 248644 157800 248694 157856
rect 248694 157800 248708 157856
rect 248644 157796 248708 157800
rect 250116 157796 250180 157860
rect 253428 157856 253492 157860
rect 253428 157800 253478 157856
rect 253478 157800 253492 157856
rect 253428 157796 253492 157800
rect 267044 157796 267108 157860
rect 212948 157660 213012 157724
rect 266492 157660 266556 157724
rect 273668 157720 273732 157724
rect 273668 157664 273718 157720
rect 273718 157664 273732 157720
rect 273668 157660 273732 157664
rect 278452 157720 278516 157724
rect 278452 157664 278502 157720
rect 278502 157664 278516 157720
rect 278452 157660 278516 157664
rect 261156 157584 261220 157588
rect 261156 157528 261206 157584
rect 261206 157528 261220 157584
rect 261156 157524 261220 157528
rect 263548 157524 263612 157588
rect 265940 157584 266004 157588
rect 265940 157528 265990 157584
rect 265990 157528 266004 157584
rect 265940 157524 266004 157528
rect 288204 157584 288268 157588
rect 288204 157528 288254 157584
rect 288254 157528 288268 157584
rect 288204 157524 288268 157528
rect 236500 157388 236564 157452
rect 363460 71844 363524 71908
rect 360332 44236 360396 44300
rect 361620 5612 361684 5676
rect 368980 4796 369044 4860
rect 360516 3980 360580 4044
rect 367324 3980 367388 4044
rect 364932 3844 364996 3908
rect 218652 3572 218716 3636
rect 358492 3708 358556 3772
rect 367692 3708 367756 3772
rect 358124 3572 358188 3636
rect 364380 3572 364444 3636
rect 365668 3572 365732 3636
rect 367140 3572 367204 3636
rect 368428 3572 368492 3636
rect 369900 3572 369964 3636
rect 213132 3436 213196 3500
rect 215156 3436 215220 3500
rect 216444 3436 216508 3500
rect 219204 3436 219268 3500
rect 214420 3300 214484 3364
rect 358308 3436 358372 3500
rect 358860 3436 358924 3500
rect 360148 3436 360212 3500
rect 362540 3436 362604 3500
rect 362908 3436 362972 3500
rect 363644 3436 363708 3500
rect 359412 3300 359476 3364
rect 369164 3300 369228 3364
rect 360700 3164 360764 3228
rect 359228 3028 359292 3092
rect 359044 2892 359108 2956
<< metal4 >>
rect -9036 711868 -8416 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 -8416 711868
rect -9036 711548 -8416 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 -8416 711548
rect -9036 682954 -8416 711312
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 -8416 682954
rect -9036 682634 -8416 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 -8416 682634
rect -9036 646954 -8416 682398
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 -8416 646954
rect -9036 646634 -8416 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 -8416 646634
rect -9036 610954 -8416 646398
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 -8416 610954
rect -9036 610634 -8416 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 -8416 610634
rect -9036 574954 -8416 610398
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 -8416 574954
rect -9036 574634 -8416 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 -8416 574634
rect -9036 538954 -8416 574398
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 -8416 538954
rect -9036 538634 -8416 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 -8416 538634
rect -9036 502954 -8416 538398
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 -8416 502954
rect -9036 502634 -8416 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 -8416 502634
rect -9036 466954 -8416 502398
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 -8416 466954
rect -9036 466634 -8416 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 -8416 466634
rect -9036 430954 -8416 466398
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 -8416 430954
rect -9036 430634 -8416 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 -8416 430634
rect -9036 394954 -8416 430398
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 -8416 394954
rect -9036 394634 -8416 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 -8416 394634
rect -9036 358954 -8416 394398
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 -8416 358954
rect -9036 358634 -8416 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 -8416 358634
rect -9036 322954 -8416 358398
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 -8416 322954
rect -9036 322634 -8416 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 -8416 322634
rect -9036 286954 -8416 322398
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 -8416 286954
rect -9036 286634 -8416 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 -8416 286634
rect -9036 250954 -8416 286398
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 -8416 250954
rect -9036 250634 -8416 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 -8416 250634
rect -9036 214954 -8416 250398
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 -8416 214954
rect -9036 214634 -8416 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 -8416 214634
rect -9036 178954 -8416 214398
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 -8416 178954
rect -9036 178634 -8416 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 -8416 178634
rect -9036 142954 -8416 178398
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 -8416 142954
rect -9036 142634 -8416 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 -8416 142634
rect -9036 106954 -8416 142398
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 -8416 106954
rect -9036 106634 -8416 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 -8416 106634
rect -9036 70954 -8416 106398
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 -8416 70954
rect -9036 70634 -8416 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 -8416 70634
rect -9036 34954 -8416 70398
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 -8416 34954
rect -9036 34634 -8416 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 -8416 34634
rect -9036 -7376 -8416 34398
rect -8076 710908 -7456 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 -7456 710908
rect -8076 710588 -7456 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 -7456 710588
rect -8076 678454 -7456 710352
rect -8076 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 -7456 678454
rect -8076 678134 -7456 678218
rect -8076 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 -7456 678134
rect -8076 642454 -7456 677898
rect -8076 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 -7456 642454
rect -8076 642134 -7456 642218
rect -8076 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 -7456 642134
rect -8076 606454 -7456 641898
rect -8076 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 -7456 606454
rect -8076 606134 -7456 606218
rect -8076 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 -7456 606134
rect -8076 570454 -7456 605898
rect -8076 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 -7456 570454
rect -8076 570134 -7456 570218
rect -8076 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 -7456 570134
rect -8076 534454 -7456 569898
rect -8076 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 -7456 534454
rect -8076 534134 -7456 534218
rect -8076 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 -7456 534134
rect -8076 498454 -7456 533898
rect -8076 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 -7456 498454
rect -8076 498134 -7456 498218
rect -8076 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 -7456 498134
rect -8076 462454 -7456 497898
rect -8076 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 -7456 462454
rect -8076 462134 -7456 462218
rect -8076 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 -7456 462134
rect -8076 426454 -7456 461898
rect -8076 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 -7456 426454
rect -8076 426134 -7456 426218
rect -8076 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 -7456 426134
rect -8076 390454 -7456 425898
rect -8076 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 -7456 390454
rect -8076 390134 -7456 390218
rect -8076 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 -7456 390134
rect -8076 354454 -7456 389898
rect -8076 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 -7456 354454
rect -8076 354134 -7456 354218
rect -8076 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 -7456 354134
rect -8076 318454 -7456 353898
rect -8076 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 -7456 318454
rect -8076 318134 -7456 318218
rect -8076 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 -7456 318134
rect -8076 282454 -7456 317898
rect -8076 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 -7456 282454
rect -8076 282134 -7456 282218
rect -8076 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 -7456 282134
rect -8076 246454 -7456 281898
rect -8076 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 -7456 246454
rect -8076 246134 -7456 246218
rect -8076 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 -7456 246134
rect -8076 210454 -7456 245898
rect -8076 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 -7456 210454
rect -8076 210134 -7456 210218
rect -8076 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 -7456 210134
rect -8076 174454 -7456 209898
rect -8076 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 -7456 174454
rect -8076 174134 -7456 174218
rect -8076 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 -7456 174134
rect -8076 138454 -7456 173898
rect -8076 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 -7456 138454
rect -8076 138134 -7456 138218
rect -8076 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 -7456 138134
rect -8076 102454 -7456 137898
rect -8076 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 -7456 102454
rect -8076 102134 -7456 102218
rect -8076 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 -7456 102134
rect -8076 66454 -7456 101898
rect -8076 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 -7456 66454
rect -8076 66134 -7456 66218
rect -8076 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 -7456 66134
rect -8076 30454 -7456 65898
rect -8076 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 -7456 30454
rect -8076 30134 -7456 30218
rect -8076 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 -7456 30134
rect -8076 -6416 -7456 29898
rect -7116 709948 -6496 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 -6496 709948
rect -7116 709628 -6496 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 -6496 709628
rect -7116 673954 -6496 709392
rect -7116 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 -6496 673954
rect -7116 673634 -6496 673718
rect -7116 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 -6496 673634
rect -7116 637954 -6496 673398
rect -7116 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 -6496 637954
rect -7116 637634 -6496 637718
rect -7116 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 -6496 637634
rect -7116 601954 -6496 637398
rect -7116 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 -6496 601954
rect -7116 601634 -6496 601718
rect -7116 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 -6496 601634
rect -7116 565954 -6496 601398
rect -7116 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 -6496 565954
rect -7116 565634 -6496 565718
rect -7116 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 -6496 565634
rect -7116 529954 -6496 565398
rect -7116 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 -6496 529954
rect -7116 529634 -6496 529718
rect -7116 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 -6496 529634
rect -7116 493954 -6496 529398
rect -7116 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 -6496 493954
rect -7116 493634 -6496 493718
rect -7116 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 -6496 493634
rect -7116 457954 -6496 493398
rect -7116 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 -6496 457954
rect -7116 457634 -6496 457718
rect -7116 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 -6496 457634
rect -7116 421954 -6496 457398
rect -7116 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 -6496 421954
rect -7116 421634 -6496 421718
rect -7116 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 -6496 421634
rect -7116 385954 -6496 421398
rect -7116 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 -6496 385954
rect -7116 385634 -6496 385718
rect -7116 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 -6496 385634
rect -7116 349954 -6496 385398
rect -7116 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 -6496 349954
rect -7116 349634 -6496 349718
rect -7116 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 -6496 349634
rect -7116 313954 -6496 349398
rect -7116 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 -6496 313954
rect -7116 313634 -6496 313718
rect -7116 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 -6496 313634
rect -7116 277954 -6496 313398
rect -7116 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 -6496 277954
rect -7116 277634 -6496 277718
rect -7116 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 -6496 277634
rect -7116 241954 -6496 277398
rect -7116 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 -6496 241954
rect -7116 241634 -6496 241718
rect -7116 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 -6496 241634
rect -7116 205954 -6496 241398
rect -7116 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 -6496 205954
rect -7116 205634 -6496 205718
rect -7116 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 -6496 205634
rect -7116 169954 -6496 205398
rect -7116 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 -6496 169954
rect -7116 169634 -6496 169718
rect -7116 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 -6496 169634
rect -7116 133954 -6496 169398
rect -7116 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 -6496 133954
rect -7116 133634 -6496 133718
rect -7116 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 -6496 133634
rect -7116 97954 -6496 133398
rect -7116 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 -6496 97954
rect -7116 97634 -6496 97718
rect -7116 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 -6496 97634
rect -7116 61954 -6496 97398
rect -7116 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 -6496 61954
rect -7116 61634 -6496 61718
rect -7116 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 -6496 61634
rect -7116 25954 -6496 61398
rect -7116 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 -6496 25954
rect -7116 25634 -6496 25718
rect -7116 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 -6496 25634
rect -7116 -5456 -6496 25398
rect -6156 708988 -5536 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 -5536 708988
rect -6156 708668 -5536 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 -5536 708668
rect -6156 669454 -5536 708432
rect -6156 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 -5536 669454
rect -6156 669134 -5536 669218
rect -6156 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 -5536 669134
rect -6156 633454 -5536 668898
rect -6156 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 -5536 633454
rect -6156 633134 -5536 633218
rect -6156 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 -5536 633134
rect -6156 597454 -5536 632898
rect -6156 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 -5536 597454
rect -6156 597134 -5536 597218
rect -6156 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 -5536 597134
rect -6156 561454 -5536 596898
rect -6156 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 -5536 561454
rect -6156 561134 -5536 561218
rect -6156 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 -5536 561134
rect -6156 525454 -5536 560898
rect -6156 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 -5536 525454
rect -6156 525134 -5536 525218
rect -6156 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 -5536 525134
rect -6156 489454 -5536 524898
rect -6156 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 -5536 489454
rect -6156 489134 -5536 489218
rect -6156 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 -5536 489134
rect -6156 453454 -5536 488898
rect -6156 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 -5536 453454
rect -6156 453134 -5536 453218
rect -6156 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 -5536 453134
rect -6156 417454 -5536 452898
rect -6156 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 -5536 417454
rect -6156 417134 -5536 417218
rect -6156 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 -5536 417134
rect -6156 381454 -5536 416898
rect -6156 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 -5536 381454
rect -6156 381134 -5536 381218
rect -6156 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 -5536 381134
rect -6156 345454 -5536 380898
rect -6156 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 -5536 345454
rect -6156 345134 -5536 345218
rect -6156 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 -5536 345134
rect -6156 309454 -5536 344898
rect -6156 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 -5536 309454
rect -6156 309134 -5536 309218
rect -6156 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 -5536 309134
rect -6156 273454 -5536 308898
rect -6156 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 -5536 273454
rect -6156 273134 -5536 273218
rect -6156 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 -5536 273134
rect -6156 237454 -5536 272898
rect -6156 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 -5536 237454
rect -6156 237134 -5536 237218
rect -6156 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 -5536 237134
rect -6156 201454 -5536 236898
rect -6156 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 -5536 201454
rect -6156 201134 -5536 201218
rect -6156 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 -5536 201134
rect -6156 165454 -5536 200898
rect -6156 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 -5536 165454
rect -6156 165134 -5536 165218
rect -6156 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 -5536 165134
rect -6156 129454 -5536 164898
rect -6156 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 -5536 129454
rect -6156 129134 -5536 129218
rect -6156 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 -5536 129134
rect -6156 93454 -5536 128898
rect -6156 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 -5536 93454
rect -6156 93134 -5536 93218
rect -6156 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 -5536 93134
rect -6156 57454 -5536 92898
rect -6156 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 -5536 57454
rect -6156 57134 -5536 57218
rect -6156 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 -5536 57134
rect -6156 21454 -5536 56898
rect -6156 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 -5536 21454
rect -6156 21134 -5536 21218
rect -6156 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 -5536 21134
rect -6156 -4496 -5536 20898
rect -5196 708028 -4576 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 -4576 708028
rect -5196 707708 -4576 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 -4576 707708
rect -5196 700954 -4576 707472
rect -5196 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 -4576 700954
rect -5196 700634 -4576 700718
rect -5196 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 -4576 700634
rect -5196 664954 -4576 700398
rect -5196 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 -4576 664954
rect -5196 664634 -4576 664718
rect -5196 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 -4576 664634
rect -5196 628954 -4576 664398
rect -5196 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 -4576 628954
rect -5196 628634 -4576 628718
rect -5196 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 -4576 628634
rect -5196 592954 -4576 628398
rect -5196 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 -4576 592954
rect -5196 592634 -4576 592718
rect -5196 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 -4576 592634
rect -5196 556954 -4576 592398
rect -5196 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 -4576 556954
rect -5196 556634 -4576 556718
rect -5196 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 -4576 556634
rect -5196 520954 -4576 556398
rect -5196 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 -4576 520954
rect -5196 520634 -4576 520718
rect -5196 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 -4576 520634
rect -5196 484954 -4576 520398
rect -5196 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 -4576 484954
rect -5196 484634 -4576 484718
rect -5196 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 -4576 484634
rect -5196 448954 -4576 484398
rect -5196 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 -4576 448954
rect -5196 448634 -4576 448718
rect -5196 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 -4576 448634
rect -5196 412954 -4576 448398
rect -5196 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 -4576 412954
rect -5196 412634 -4576 412718
rect -5196 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 -4576 412634
rect -5196 376954 -4576 412398
rect -5196 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 -4576 376954
rect -5196 376634 -4576 376718
rect -5196 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 -4576 376634
rect -5196 340954 -4576 376398
rect -5196 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 -4576 340954
rect -5196 340634 -4576 340718
rect -5196 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 -4576 340634
rect -5196 304954 -4576 340398
rect -5196 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 -4576 304954
rect -5196 304634 -4576 304718
rect -5196 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 -4576 304634
rect -5196 268954 -4576 304398
rect -5196 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 -4576 268954
rect -5196 268634 -4576 268718
rect -5196 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 -4576 268634
rect -5196 232954 -4576 268398
rect -5196 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 -4576 232954
rect -5196 232634 -4576 232718
rect -5196 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 -4576 232634
rect -5196 196954 -4576 232398
rect -5196 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 -4576 196954
rect -5196 196634 -4576 196718
rect -5196 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 -4576 196634
rect -5196 160954 -4576 196398
rect -5196 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 -4576 160954
rect -5196 160634 -4576 160718
rect -5196 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 -4576 160634
rect -5196 124954 -4576 160398
rect -5196 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 -4576 124954
rect -5196 124634 -4576 124718
rect -5196 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 -4576 124634
rect -5196 88954 -4576 124398
rect -5196 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 -4576 88954
rect -5196 88634 -4576 88718
rect -5196 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 -4576 88634
rect -5196 52954 -4576 88398
rect -5196 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 -4576 52954
rect -5196 52634 -4576 52718
rect -5196 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 -4576 52634
rect -5196 16954 -4576 52398
rect -5196 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 -4576 16954
rect -5196 16634 -4576 16718
rect -5196 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 -4576 16634
rect -5196 -3536 -4576 16398
rect -4236 707068 -3616 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 -3616 707068
rect -4236 706748 -3616 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 -3616 706748
rect -4236 696454 -3616 706512
rect -4236 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 -3616 696454
rect -4236 696134 -3616 696218
rect -4236 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 -3616 696134
rect -4236 660454 -3616 695898
rect -4236 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 -3616 660454
rect -4236 660134 -3616 660218
rect -4236 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 -3616 660134
rect -4236 624454 -3616 659898
rect -4236 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 -3616 624454
rect -4236 624134 -3616 624218
rect -4236 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 -3616 624134
rect -4236 588454 -3616 623898
rect -4236 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 -3616 588454
rect -4236 588134 -3616 588218
rect -4236 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 -3616 588134
rect -4236 552454 -3616 587898
rect -4236 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 -3616 552454
rect -4236 552134 -3616 552218
rect -4236 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 -3616 552134
rect -4236 516454 -3616 551898
rect -4236 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 -3616 516454
rect -4236 516134 -3616 516218
rect -4236 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 -3616 516134
rect -4236 480454 -3616 515898
rect -4236 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 -3616 480454
rect -4236 480134 -3616 480218
rect -4236 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 -3616 480134
rect -4236 444454 -3616 479898
rect -4236 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 -3616 444454
rect -4236 444134 -3616 444218
rect -4236 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 -3616 444134
rect -4236 408454 -3616 443898
rect -4236 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 -3616 408454
rect -4236 408134 -3616 408218
rect -4236 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 -3616 408134
rect -4236 372454 -3616 407898
rect -4236 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 -3616 372454
rect -4236 372134 -3616 372218
rect -4236 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 -3616 372134
rect -4236 336454 -3616 371898
rect -4236 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 -3616 336454
rect -4236 336134 -3616 336218
rect -4236 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 -3616 336134
rect -4236 300454 -3616 335898
rect -4236 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 -3616 300454
rect -4236 300134 -3616 300218
rect -4236 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 -3616 300134
rect -4236 264454 -3616 299898
rect -4236 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 -3616 264454
rect -4236 264134 -3616 264218
rect -4236 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 -3616 264134
rect -4236 228454 -3616 263898
rect -4236 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 -3616 228454
rect -4236 228134 -3616 228218
rect -4236 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 -3616 228134
rect -4236 192454 -3616 227898
rect -4236 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 -3616 192454
rect -4236 192134 -3616 192218
rect -4236 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 -3616 192134
rect -4236 156454 -3616 191898
rect -4236 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 -3616 156454
rect -4236 156134 -3616 156218
rect -4236 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 -3616 156134
rect -4236 120454 -3616 155898
rect -4236 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 -3616 120454
rect -4236 120134 -3616 120218
rect -4236 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 -3616 120134
rect -4236 84454 -3616 119898
rect -4236 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 -3616 84454
rect -4236 84134 -3616 84218
rect -4236 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 -3616 84134
rect -4236 48454 -3616 83898
rect -4236 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 -3616 48454
rect -4236 48134 -3616 48218
rect -4236 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 -3616 48134
rect -4236 12454 -3616 47898
rect -4236 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 -3616 12454
rect -4236 12134 -3616 12218
rect -4236 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 -3616 12134
rect -4236 -2576 -3616 11898
rect -3276 706108 -2656 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 -2656 706108
rect -3276 705788 -2656 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 -2656 705788
rect -3276 691954 -2656 705552
rect -3276 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 -2656 691954
rect -3276 691634 -2656 691718
rect -3276 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 -2656 691634
rect -3276 655954 -2656 691398
rect -3276 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 -2656 655954
rect -3276 655634 -2656 655718
rect -3276 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 -2656 655634
rect -3276 619954 -2656 655398
rect -3276 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 -2656 619954
rect -3276 619634 -2656 619718
rect -3276 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 -2656 619634
rect -3276 583954 -2656 619398
rect -3276 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 -2656 583954
rect -3276 583634 -2656 583718
rect -3276 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 -2656 583634
rect -3276 547954 -2656 583398
rect -3276 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 -2656 547954
rect -3276 547634 -2656 547718
rect -3276 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 -2656 547634
rect -3276 511954 -2656 547398
rect -3276 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 -2656 511954
rect -3276 511634 -2656 511718
rect -3276 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 -2656 511634
rect -3276 475954 -2656 511398
rect -3276 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 -2656 475954
rect -3276 475634 -2656 475718
rect -3276 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 -2656 475634
rect -3276 439954 -2656 475398
rect -3276 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 -2656 439954
rect -3276 439634 -2656 439718
rect -3276 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 -2656 439634
rect -3276 403954 -2656 439398
rect -3276 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 -2656 403954
rect -3276 403634 -2656 403718
rect -3276 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 -2656 403634
rect -3276 367954 -2656 403398
rect -3276 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 -2656 367954
rect -3276 367634 -2656 367718
rect -3276 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 -2656 367634
rect -3276 331954 -2656 367398
rect -3276 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 -2656 331954
rect -3276 331634 -2656 331718
rect -3276 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 -2656 331634
rect -3276 295954 -2656 331398
rect -3276 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 -2656 295954
rect -3276 295634 -2656 295718
rect -3276 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 -2656 295634
rect -3276 259954 -2656 295398
rect -3276 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 -2656 259954
rect -3276 259634 -2656 259718
rect -3276 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 -2656 259634
rect -3276 223954 -2656 259398
rect -3276 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 -2656 223954
rect -3276 223634 -2656 223718
rect -3276 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 -2656 223634
rect -3276 187954 -2656 223398
rect -3276 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 -2656 187954
rect -3276 187634 -2656 187718
rect -3276 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 -2656 187634
rect -3276 151954 -2656 187398
rect -3276 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 -2656 151954
rect -3276 151634 -2656 151718
rect -3276 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 -2656 151634
rect -3276 115954 -2656 151398
rect -3276 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 -2656 115954
rect -3276 115634 -2656 115718
rect -3276 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 -2656 115634
rect -3276 79954 -2656 115398
rect -3276 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 -2656 79954
rect -3276 79634 -2656 79718
rect -3276 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 -2656 79634
rect -3276 43954 -2656 79398
rect -3276 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 -2656 43954
rect -3276 43634 -2656 43718
rect -3276 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 -2656 43634
rect -3276 7954 -2656 43398
rect -3276 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 -2656 7954
rect -3276 7634 -2656 7718
rect -3276 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 -2656 7634
rect -3276 -1616 -2656 7398
rect -2316 705148 -1696 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 -1696 705148
rect -2316 704828 -1696 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 -1696 704828
rect -2316 687454 -1696 704592
rect -2316 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 -1696 687454
rect -2316 687134 -1696 687218
rect -2316 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 -1696 687134
rect -2316 651454 -1696 686898
rect -2316 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 -1696 651454
rect -2316 651134 -1696 651218
rect -2316 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 -1696 651134
rect -2316 615454 -1696 650898
rect -2316 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 -1696 615454
rect -2316 615134 -1696 615218
rect -2316 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 -1696 615134
rect -2316 579454 -1696 614898
rect -2316 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 -1696 579454
rect -2316 579134 -1696 579218
rect -2316 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 -1696 579134
rect -2316 543454 -1696 578898
rect -2316 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 -1696 543454
rect -2316 543134 -1696 543218
rect -2316 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 -1696 543134
rect -2316 507454 -1696 542898
rect -2316 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 -1696 507454
rect -2316 507134 -1696 507218
rect -2316 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 -1696 507134
rect -2316 471454 -1696 506898
rect -2316 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 -1696 471454
rect -2316 471134 -1696 471218
rect -2316 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 -1696 471134
rect -2316 435454 -1696 470898
rect -2316 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 -1696 435454
rect -2316 435134 -1696 435218
rect -2316 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 -1696 435134
rect -2316 399454 -1696 434898
rect -2316 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 -1696 399454
rect -2316 399134 -1696 399218
rect -2316 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 -1696 399134
rect -2316 363454 -1696 398898
rect -2316 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 -1696 363454
rect -2316 363134 -1696 363218
rect -2316 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 -1696 363134
rect -2316 327454 -1696 362898
rect -2316 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 -1696 327454
rect -2316 327134 -1696 327218
rect -2316 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 -1696 327134
rect -2316 291454 -1696 326898
rect -2316 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 -1696 291454
rect -2316 291134 -1696 291218
rect -2316 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 -1696 291134
rect -2316 255454 -1696 290898
rect -2316 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 -1696 255454
rect -2316 255134 -1696 255218
rect -2316 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 -1696 255134
rect -2316 219454 -1696 254898
rect -2316 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 -1696 219454
rect -2316 219134 -1696 219218
rect -2316 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 -1696 219134
rect -2316 183454 -1696 218898
rect -2316 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 -1696 183454
rect -2316 183134 -1696 183218
rect -2316 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 -1696 183134
rect -2316 147454 -1696 182898
rect -2316 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 -1696 147454
rect -2316 147134 -1696 147218
rect -2316 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 -1696 147134
rect -2316 111454 -1696 146898
rect -2316 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 -1696 111454
rect -2316 111134 -1696 111218
rect -2316 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 -1696 111134
rect -2316 75454 -1696 110898
rect -2316 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 -1696 75454
rect -2316 75134 -1696 75218
rect -2316 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 -1696 75134
rect -2316 39454 -1696 74898
rect -2316 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 -1696 39454
rect -2316 39134 -1696 39218
rect -2316 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 -1696 39134
rect -2316 3454 -1696 38898
rect -2316 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 -1696 3454
rect -2316 3134 -1696 3218
rect -2316 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 -1696 3134
rect -2316 -656 -1696 2898
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 -1696 -656
rect -2316 -976 -1696 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 -1696 -976
rect -2316 -1244 -1696 -1212
rect 1794 705148 2414 711900
rect 1794 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 2414 705148
rect 1794 704828 2414 704912
rect 1794 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 2414 704828
rect 1794 687454 2414 704592
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -656 2414 2898
rect 1794 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 2414 -656
rect 1794 -976 2414 -892
rect 1794 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 2414 -976
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 -2656 -1616
rect -3276 -1936 -2656 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 -2656 -1936
rect -3276 -2204 -2656 -2172
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 -3616 -2576
rect -4236 -2896 -3616 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 -3616 -2896
rect -4236 -3164 -3616 -3132
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 -4576 -3536
rect -5196 -3856 -4576 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 -4576 -3856
rect -5196 -4124 -4576 -4092
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 -5536 -4496
rect -6156 -4816 -5536 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 -5536 -4816
rect -6156 -5084 -5536 -5052
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 -6496 -5456
rect -7116 -5776 -6496 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 -6496 -5776
rect -7116 -6044 -6496 -6012
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 -7456 -6416
rect -8076 -6736 -7456 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 -7456 -6736
rect -8076 -7004 -7456 -6972
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 -8416 -7376
rect -9036 -7696 -8416 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 -8416 -7696
rect -9036 -7964 -8416 -7932
rect 1794 -7964 2414 -1212
rect 6294 706108 6914 711900
rect 6294 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 6914 706108
rect 6294 705788 6914 705872
rect 6294 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 6914 705788
rect 6294 691954 6914 705552
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1616 6914 7398
rect 6294 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 6914 -1616
rect 6294 -1936 6914 -1852
rect 6294 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 6914 -1936
rect 6294 -7964 6914 -2172
rect 10794 707068 11414 711900
rect 10794 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 11414 707068
rect 10794 706748 11414 706832
rect 10794 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 11414 706748
rect 10794 696454 11414 706512
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2576 11414 11898
rect 10794 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 11414 -2576
rect 10794 -2896 11414 -2812
rect 10794 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 11414 -2896
rect 10794 -7964 11414 -3132
rect 15294 708028 15914 711900
rect 15294 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 15914 708028
rect 15294 707708 15914 707792
rect 15294 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 15914 707708
rect 15294 700954 15914 707472
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3536 15914 16398
rect 15294 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 15914 -3536
rect 15294 -3856 15914 -3772
rect 15294 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 15914 -3856
rect 15294 -7964 15914 -4092
rect 19794 708988 20414 711900
rect 19794 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 20414 708988
rect 19794 708668 20414 708752
rect 19794 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 20414 708668
rect 19794 669454 20414 708432
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4496 20414 20898
rect 19794 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 20414 -4496
rect 19794 -4816 20414 -4732
rect 19794 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 20414 -4816
rect 19794 -7964 20414 -5052
rect 24294 709948 24914 711900
rect 24294 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 24914 709948
rect 24294 709628 24914 709712
rect 24294 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 24914 709628
rect 24294 673954 24914 709392
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5456 24914 25398
rect 24294 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 24914 -5456
rect 24294 -5776 24914 -5692
rect 24294 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 24914 -5776
rect 24294 -7964 24914 -6012
rect 28794 710908 29414 711900
rect 28794 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 29414 710908
rect 28794 710588 29414 710672
rect 28794 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 29414 710588
rect 28794 678454 29414 710352
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6416 29414 29898
rect 28794 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 29414 -6416
rect 28794 -6736 29414 -6652
rect 28794 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 29414 -6736
rect 28794 -7964 29414 -6972
rect 33294 711868 33914 711900
rect 33294 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 33914 711868
rect 33294 711548 33914 711632
rect 33294 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 33914 711548
rect 33294 682954 33914 711312
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7376 33914 34398
rect 33294 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 33914 -7376
rect 33294 -7696 33914 -7612
rect 33294 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 33914 -7696
rect 33294 -7964 33914 -7932
rect 37794 705148 38414 711900
rect 37794 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 38414 705148
rect 37794 704828 38414 704912
rect 37794 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 38414 704828
rect 37794 687454 38414 704592
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -656 38414 2898
rect 37794 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 38414 -656
rect 37794 -976 38414 -892
rect 37794 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 38414 -976
rect 37794 -7964 38414 -1212
rect 42294 706108 42914 711900
rect 42294 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 42914 706108
rect 42294 705788 42914 705872
rect 42294 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 42914 705788
rect 42294 691954 42914 705552
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1616 42914 7398
rect 42294 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 42914 -1616
rect 42294 -1936 42914 -1852
rect 42294 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 42914 -1936
rect 42294 -7964 42914 -2172
rect 46794 707068 47414 711900
rect 46794 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 47414 707068
rect 46794 706748 47414 706832
rect 46794 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 47414 706748
rect 46794 696454 47414 706512
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2576 47414 11898
rect 46794 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 47414 -2576
rect 46794 -2896 47414 -2812
rect 46794 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 47414 -2896
rect 46794 -7964 47414 -3132
rect 51294 708028 51914 711900
rect 51294 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 51914 708028
rect 51294 707708 51914 707792
rect 51294 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 51914 707708
rect 51294 700954 51914 707472
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3536 51914 16398
rect 51294 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 51914 -3536
rect 51294 -3856 51914 -3772
rect 51294 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 51914 -3856
rect 51294 -7964 51914 -4092
rect 55794 708988 56414 711900
rect 55794 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 56414 708988
rect 55794 708668 56414 708752
rect 55794 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 56414 708668
rect 55794 669454 56414 708432
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4496 56414 20898
rect 55794 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 56414 -4496
rect 55794 -4816 56414 -4732
rect 55794 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 56414 -4816
rect 55794 -7964 56414 -5052
rect 60294 709948 60914 711900
rect 60294 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 60914 709948
rect 60294 709628 60914 709712
rect 60294 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 60914 709628
rect 60294 673954 60914 709392
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5456 60914 25398
rect 60294 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 60914 -5456
rect 60294 -5776 60914 -5692
rect 60294 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 60914 -5776
rect 60294 -7964 60914 -6012
rect 64794 710908 65414 711900
rect 64794 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 65414 710908
rect 64794 710588 65414 710672
rect 64794 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 65414 710588
rect 64794 678454 65414 710352
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6416 65414 29898
rect 64794 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 65414 -6416
rect 64794 -6736 65414 -6652
rect 64794 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 65414 -6736
rect 64794 -7964 65414 -6972
rect 69294 711868 69914 711900
rect 69294 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 69914 711868
rect 69294 711548 69914 711632
rect 69294 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 69914 711548
rect 69294 682954 69914 711312
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7376 69914 34398
rect 69294 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 69914 -7376
rect 69294 -7696 69914 -7612
rect 69294 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 69914 -7696
rect 69294 -7964 69914 -7932
rect 73794 705148 74414 711900
rect 73794 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 74414 705148
rect 73794 704828 74414 704912
rect 73794 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 74414 704828
rect 73794 687454 74414 704592
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -656 74414 2898
rect 73794 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 74414 -656
rect 73794 -976 74414 -892
rect 73794 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 74414 -976
rect 73794 -7964 74414 -1212
rect 78294 706108 78914 711900
rect 78294 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 78914 706108
rect 78294 705788 78914 705872
rect 78294 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 78914 705788
rect 78294 691954 78914 705552
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1616 78914 7398
rect 78294 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 78914 -1616
rect 78294 -1936 78914 -1852
rect 78294 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 78914 -1936
rect 78294 -7964 78914 -2172
rect 82794 707068 83414 711900
rect 82794 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 83414 707068
rect 82794 706748 83414 706832
rect 82794 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 83414 706748
rect 82794 696454 83414 706512
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2576 83414 11898
rect 82794 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 83414 -2576
rect 82794 -2896 83414 -2812
rect 82794 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 83414 -2896
rect 82794 -7964 83414 -3132
rect 87294 708028 87914 711900
rect 87294 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 87914 708028
rect 87294 707708 87914 707792
rect 87294 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 87914 707708
rect 87294 700954 87914 707472
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3536 87914 16398
rect 87294 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 87914 -3536
rect 87294 -3856 87914 -3772
rect 87294 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 87914 -3856
rect 87294 -7964 87914 -4092
rect 91794 708988 92414 711900
rect 91794 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 92414 708988
rect 91794 708668 92414 708752
rect 91794 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 92414 708668
rect 91794 669454 92414 708432
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4496 92414 20898
rect 91794 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 92414 -4496
rect 91794 -4816 92414 -4732
rect 91794 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 92414 -4816
rect 91794 -7964 92414 -5052
rect 96294 709948 96914 711900
rect 96294 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 96914 709948
rect 96294 709628 96914 709712
rect 96294 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 96914 709628
rect 96294 673954 96914 709392
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5456 96914 25398
rect 96294 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 96914 -5456
rect 96294 -5776 96914 -5692
rect 96294 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 96914 -5776
rect 96294 -7964 96914 -6012
rect 100794 710908 101414 711900
rect 100794 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 101414 710908
rect 100794 710588 101414 710672
rect 100794 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 101414 710588
rect 100794 678454 101414 710352
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6416 101414 29898
rect 100794 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 101414 -6416
rect 100794 -6736 101414 -6652
rect 100794 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 101414 -6736
rect 100794 -7964 101414 -6972
rect 105294 711868 105914 711900
rect 105294 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 105914 711868
rect 105294 711548 105914 711632
rect 105294 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 105914 711548
rect 105294 682954 105914 711312
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7376 105914 34398
rect 105294 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 105914 -7376
rect 105294 -7696 105914 -7612
rect 105294 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 105914 -7696
rect 105294 -7964 105914 -7932
rect 109794 705148 110414 711900
rect 109794 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 110414 705148
rect 109794 704828 110414 704912
rect 109794 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 110414 704828
rect 109794 687454 110414 704592
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -656 110414 2898
rect 109794 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 110414 -656
rect 109794 -976 110414 -892
rect 109794 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 110414 -976
rect 109794 -7964 110414 -1212
rect 114294 706108 114914 711900
rect 114294 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 114914 706108
rect 114294 705788 114914 705872
rect 114294 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 114914 705788
rect 114294 691954 114914 705552
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1616 114914 7398
rect 114294 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 114914 -1616
rect 114294 -1936 114914 -1852
rect 114294 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 114914 -1936
rect 114294 -7964 114914 -2172
rect 118794 707068 119414 711900
rect 118794 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 119414 707068
rect 118794 706748 119414 706832
rect 118794 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 119414 706748
rect 118794 696454 119414 706512
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2576 119414 11898
rect 118794 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 119414 -2576
rect 118794 -2896 119414 -2812
rect 118794 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 119414 -2896
rect 118794 -7964 119414 -3132
rect 123294 708028 123914 711900
rect 123294 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 123914 708028
rect 123294 707708 123914 707792
rect 123294 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 123914 707708
rect 123294 700954 123914 707472
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3536 123914 16398
rect 123294 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 123914 -3536
rect 123294 -3856 123914 -3772
rect 123294 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 123914 -3856
rect 123294 -7964 123914 -4092
rect 127794 708988 128414 711900
rect 127794 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 128414 708988
rect 127794 708668 128414 708752
rect 127794 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 128414 708668
rect 127794 669454 128414 708432
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4496 128414 20898
rect 127794 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 128414 -4496
rect 127794 -4816 128414 -4732
rect 127794 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 128414 -4816
rect 127794 -7964 128414 -5052
rect 132294 709948 132914 711900
rect 132294 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 132914 709948
rect 132294 709628 132914 709712
rect 132294 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 132914 709628
rect 132294 673954 132914 709392
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5456 132914 25398
rect 132294 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 132914 -5456
rect 132294 -5776 132914 -5692
rect 132294 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 132914 -5776
rect 132294 -7964 132914 -6012
rect 136794 710908 137414 711900
rect 136794 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 137414 710908
rect 136794 710588 137414 710672
rect 136794 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 137414 710588
rect 136794 678454 137414 710352
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6416 137414 29898
rect 136794 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 137414 -6416
rect 136794 -6736 137414 -6652
rect 136794 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 137414 -6736
rect 136794 -7964 137414 -6972
rect 141294 711868 141914 711900
rect 141294 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 141914 711868
rect 141294 711548 141914 711632
rect 141294 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 141914 711548
rect 141294 682954 141914 711312
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7376 141914 34398
rect 141294 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 141914 -7376
rect 141294 -7696 141914 -7612
rect 141294 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 141914 -7696
rect 141294 -7964 141914 -7932
rect 145794 705148 146414 711900
rect 145794 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 146414 705148
rect 145794 704828 146414 704912
rect 145794 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 146414 704828
rect 145794 687454 146414 704592
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -656 146414 2898
rect 145794 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 146414 -656
rect 145794 -976 146414 -892
rect 145794 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 146414 -976
rect 145794 -7964 146414 -1212
rect 150294 706108 150914 711900
rect 150294 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 150914 706108
rect 150294 705788 150914 705872
rect 150294 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 150914 705788
rect 150294 691954 150914 705552
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1616 150914 7398
rect 150294 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 150914 -1616
rect 150294 -1936 150914 -1852
rect 150294 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 150914 -1936
rect 150294 -7964 150914 -2172
rect 154794 707068 155414 711900
rect 154794 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 155414 707068
rect 154794 706748 155414 706832
rect 154794 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 155414 706748
rect 154794 696454 155414 706512
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2576 155414 11898
rect 154794 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 155414 -2576
rect 154794 -2896 155414 -2812
rect 154794 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 155414 -2896
rect 154794 -7964 155414 -3132
rect 159294 708028 159914 711900
rect 159294 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 159914 708028
rect 159294 707708 159914 707792
rect 159294 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 159914 707708
rect 159294 700954 159914 707472
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3536 159914 16398
rect 159294 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 159914 -3536
rect 159294 -3856 159914 -3772
rect 159294 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 159914 -3856
rect 159294 -7964 159914 -4092
rect 163794 708988 164414 711900
rect 163794 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 164414 708988
rect 163794 708668 164414 708752
rect 163794 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 164414 708668
rect 163794 669454 164414 708432
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4496 164414 20898
rect 163794 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 164414 -4496
rect 163794 -4816 164414 -4732
rect 163794 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 164414 -4816
rect 163794 -7964 164414 -5052
rect 168294 709948 168914 711900
rect 168294 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 168914 709948
rect 168294 709628 168914 709712
rect 168294 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 168914 709628
rect 168294 673954 168914 709392
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5456 168914 25398
rect 168294 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 168914 -5456
rect 168294 -5776 168914 -5692
rect 168294 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 168914 -5776
rect 168294 -7964 168914 -6012
rect 172794 710908 173414 711900
rect 172794 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 173414 710908
rect 172794 710588 173414 710672
rect 172794 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 173414 710588
rect 172794 678454 173414 710352
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6416 173414 29898
rect 172794 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 173414 -6416
rect 172794 -6736 173414 -6652
rect 172794 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 173414 -6736
rect 172794 -7964 173414 -6972
rect 177294 711868 177914 711900
rect 177294 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 177914 711868
rect 177294 711548 177914 711632
rect 177294 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 177914 711548
rect 177294 682954 177914 711312
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7376 177914 34398
rect 177294 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 177914 -7376
rect 177294 -7696 177914 -7612
rect 177294 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 177914 -7696
rect 177294 -7964 177914 -7932
rect 181794 705148 182414 711900
rect 181794 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 182414 705148
rect 181794 704828 182414 704912
rect 181794 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 182414 704828
rect 181794 687454 182414 704592
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -656 182414 2898
rect 181794 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 182414 -656
rect 181794 -976 182414 -892
rect 181794 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 182414 -976
rect 181794 -7964 182414 -1212
rect 186294 706108 186914 711900
rect 186294 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 186914 706108
rect 186294 705788 186914 705872
rect 186294 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 186914 705788
rect 186294 691954 186914 705552
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1616 186914 7398
rect 186294 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 186914 -1616
rect 186294 -1936 186914 -1852
rect 186294 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 186914 -1936
rect 186294 -7964 186914 -2172
rect 190794 707068 191414 711900
rect 190794 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 191414 707068
rect 190794 706748 191414 706832
rect 190794 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 191414 706748
rect 190794 696454 191414 706512
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2576 191414 11898
rect 190794 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 191414 -2576
rect 190794 -2896 191414 -2812
rect 190794 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 191414 -2896
rect 190794 -7964 191414 -3132
rect 195294 708028 195914 711900
rect 195294 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 195914 708028
rect 195294 707708 195914 707792
rect 195294 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 195914 707708
rect 195294 700954 195914 707472
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3536 195914 16398
rect 195294 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 195914 -3536
rect 195294 -3856 195914 -3772
rect 195294 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 195914 -3856
rect 195294 -7964 195914 -4092
rect 199794 708988 200414 711900
rect 199794 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 200414 708988
rect 199794 708668 200414 708752
rect 199794 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 200414 708668
rect 199794 669454 200414 708432
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4496 200414 20898
rect 199794 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 200414 -4496
rect 199794 -4816 200414 -4732
rect 199794 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 200414 -4816
rect 199794 -7964 200414 -5052
rect 204294 709948 204914 711900
rect 204294 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 204914 709948
rect 204294 709628 204914 709712
rect 204294 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 204914 709628
rect 204294 673954 204914 709392
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5456 204914 25398
rect 204294 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 204914 -5456
rect 204294 -5776 204914 -5692
rect 204294 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 204914 -5776
rect 204294 -7964 204914 -6012
rect 208794 710908 209414 711900
rect 208794 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 209414 710908
rect 208794 710588 209414 710672
rect 208794 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 209414 710588
rect 208794 678454 209414 710352
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 213294 711868 213914 711900
rect 213294 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 213914 711868
rect 213294 711548 213914 711632
rect 213294 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 213914 711548
rect 213294 682954 213914 711312
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 705148 218414 711900
rect 217794 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 218414 705148
rect 217794 704828 218414 704912
rect 217794 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 218414 704828
rect 217794 687454 218414 704592
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 706108 222914 711900
rect 222294 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 222914 706108
rect 222294 705788 222914 705872
rect 222294 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 222914 705788
rect 222294 691954 222914 705552
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 707068 227414 711900
rect 226794 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 227414 707068
rect 226794 706748 227414 706832
rect 226794 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 227414 706748
rect 226794 696454 227414 706512
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 708028 231914 711900
rect 231294 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 231914 708028
rect 231294 707708 231914 707792
rect 231294 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 231914 707708
rect 231294 700954 231914 707472
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708988 236414 711900
rect 235794 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 236414 708988
rect 235794 708668 236414 708752
rect 235794 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 236414 708668
rect 235794 669454 236414 708432
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709948 240914 711900
rect 240294 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 240914 709948
rect 240294 709628 240914 709712
rect 240294 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 240914 709628
rect 240294 673954 240914 709392
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710908 245414 711900
rect 244794 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 245414 710908
rect 244794 710588 245414 710672
rect 244794 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 245414 710588
rect 244794 678454 245414 710352
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711868 249914 711900
rect 249294 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 249914 711868
rect 249294 711548 249914 711632
rect 249294 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 249914 711548
rect 249294 682954 249914 711312
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 705148 254414 711900
rect 253794 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 254414 705148
rect 253794 704828 254414 704912
rect 253794 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 254414 704828
rect 253794 687454 254414 704592
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 706108 258914 711900
rect 258294 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 258914 706108
rect 258294 705788 258914 705872
rect 258294 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 258914 705788
rect 258294 691954 258914 705552
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 707068 263414 711900
rect 262794 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 263414 707068
rect 262794 706748 263414 706832
rect 262794 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 263414 706748
rect 262794 696454 263414 706512
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 708028 267914 711900
rect 267294 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 267914 708028
rect 267294 707708 267914 707792
rect 267294 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 267914 707708
rect 267294 700954 267914 707472
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708988 272414 711900
rect 271794 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 272414 708988
rect 271794 708668 272414 708752
rect 271794 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 272414 708668
rect 271794 669454 272414 708432
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709948 276914 711900
rect 276294 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 276914 709948
rect 276294 709628 276914 709712
rect 276294 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 276914 709628
rect 276294 673954 276914 709392
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710908 281414 711900
rect 280794 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 281414 710908
rect 280794 710588 281414 710672
rect 280794 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 281414 710588
rect 280794 678454 281414 710352
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711868 285914 711900
rect 285294 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 285914 711868
rect 285294 711548 285914 711632
rect 285294 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 285914 711548
rect 285294 682954 285914 711312
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 705148 290414 711900
rect 289794 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 290414 705148
rect 289794 704828 290414 704912
rect 289794 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 290414 704828
rect 289794 687454 290414 704592
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 706108 294914 711900
rect 294294 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 294914 706108
rect 294294 705788 294914 705872
rect 294294 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 294914 705788
rect 294294 691954 294914 705552
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 707068 299414 711900
rect 298794 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 299414 707068
rect 298794 706748 299414 706832
rect 298794 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 299414 706748
rect 298794 696454 299414 706512
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 708028 303914 711900
rect 303294 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 303914 708028
rect 303294 707708 303914 707792
rect 303294 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 303914 707708
rect 303294 700954 303914 707472
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708988 308414 711900
rect 307794 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 308414 708988
rect 307794 708668 308414 708752
rect 307794 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 308414 708668
rect 307794 669454 308414 708432
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709948 312914 711900
rect 312294 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 312914 709948
rect 312294 709628 312914 709712
rect 312294 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 312914 709628
rect 312294 673954 312914 709392
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710908 317414 711900
rect 316794 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 317414 710908
rect 316794 710588 317414 710672
rect 316794 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 317414 710588
rect 316794 678454 317414 710352
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711868 321914 711900
rect 321294 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 321914 711868
rect 321294 711548 321914 711632
rect 321294 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 321914 711548
rect 321294 682954 321914 711312
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 705148 326414 711900
rect 325794 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 326414 705148
rect 325794 704828 326414 704912
rect 325794 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 326414 704828
rect 325794 687454 326414 704592
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 706108 330914 711900
rect 330294 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 330914 706108
rect 330294 705788 330914 705872
rect 330294 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 330914 705788
rect 330294 691954 330914 705552
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 707068 335414 711900
rect 334794 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 335414 707068
rect 334794 706748 335414 706832
rect 334794 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 335414 706748
rect 334794 696454 335414 706512
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 708028 339914 711900
rect 339294 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 339914 708028
rect 339294 707708 339914 707792
rect 339294 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 339914 707708
rect 339294 700954 339914 707472
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708988 344414 711900
rect 343794 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 344414 708988
rect 343794 708668 344414 708752
rect 343794 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 344414 708668
rect 343794 669454 344414 708432
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709948 348914 711900
rect 348294 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 348914 709948
rect 348294 709628 348914 709712
rect 348294 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 348914 709628
rect 348294 673954 348914 709392
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710908 353414 711900
rect 352794 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 353414 710908
rect 352794 710588 353414 710672
rect 352794 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 353414 710588
rect 352794 678454 353414 710352
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711868 357914 711900
rect 357294 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 357914 711868
rect 357294 711548 357914 711632
rect 357294 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 357914 711548
rect 357294 682954 357914 711312
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 705148 362414 711900
rect 361794 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 362414 705148
rect 361794 704828 362414 704912
rect 361794 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 362414 704828
rect 361794 687454 362414 704592
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 235950 479710 236116 479770
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 237144 479710 237298 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 214603 443188 214669 443189
rect 214603 443124 214604 443188
rect 214668 443124 214669 443188
rect 214603 443123 214669 443124
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 212947 303108 213013 303109
rect 212947 303044 212948 303108
rect 213012 303044 213013 303108
rect 212947 303043 213013 303044
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 212950 157725 213010 303043
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 214419 273868 214485 273869
rect 214419 273804 214420 273868
rect 214484 273804 214485 273868
rect 214419 273803 214485 273804
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213131 249116 213197 249117
rect 213131 249052 213132 249116
rect 213196 249052 213197 249116
rect 213131 249051 213197 249052
rect 212947 157724 213013 157725
rect 212947 157660 212948 157724
rect 213012 157660 213013 157724
rect 212947 157659 213013 157660
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6416 209414 29898
rect 213134 3501 213194 249051
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213131 3500 213197 3501
rect 213131 3436 213132 3500
rect 213196 3436 213197 3500
rect 213131 3435 213197 3436
rect 208794 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 209414 -6416
rect 208794 -6736 209414 -6652
rect 208794 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 209414 -6736
rect 208794 -7964 209414 -6972
rect 213294 -7376 213914 34398
rect 214422 3365 214482 273803
rect 214606 214029 214666 443123
rect 215891 443052 215957 443053
rect 215891 442988 215892 443052
rect 215956 442988 215957 443052
rect 215891 442987 215957 442988
rect 214971 306100 215037 306101
rect 214971 306036 214972 306100
rect 215036 306036 215037 306100
rect 214971 306035 215037 306036
rect 214603 214028 214669 214029
rect 214603 213964 214604 214028
rect 214668 213964 214669 214028
rect 214603 213963 214669 213964
rect 214974 158677 215034 306035
rect 215155 267068 215221 267069
rect 215155 267004 215156 267068
rect 215220 267004 215221 267068
rect 215155 267003 215221 267004
rect 214971 158676 215037 158677
rect 214971 158612 214972 158676
rect 215036 158612 215037 158676
rect 214971 158611 215037 158612
rect 215158 3501 215218 267003
rect 215894 162893 215954 442987
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217363 308684 217429 308685
rect 217363 308620 217364 308684
rect 217428 308620 217429 308684
rect 217363 308619 217429 308620
rect 216075 306236 216141 306237
rect 216075 306172 216076 306236
rect 216140 306172 216141 306236
rect 216075 306171 216141 306172
rect 215891 162892 215957 162893
rect 215891 162828 215892 162892
rect 215956 162828 215957 162892
rect 215891 162827 215957 162828
rect 216078 158133 216138 306171
rect 216259 305964 216325 305965
rect 216259 305900 216260 305964
rect 216324 305900 216325 305964
rect 216259 305899 216325 305900
rect 216262 158269 216322 305899
rect 216995 305828 217061 305829
rect 216995 305764 216996 305828
rect 217060 305764 217061 305828
rect 216995 305763 217061 305764
rect 216443 275228 216509 275229
rect 216443 275164 216444 275228
rect 216508 275164 216509 275228
rect 216443 275163 216509 275164
rect 216259 158268 216325 158269
rect 216259 158204 216260 158268
rect 216324 158204 216325 158268
rect 216259 158203 216325 158204
rect 216075 158132 216141 158133
rect 216075 158068 216076 158132
rect 216140 158068 216141 158132
rect 216075 158067 216141 158068
rect 216446 3501 216506 275163
rect 216998 157997 217058 305763
rect 217179 305692 217245 305693
rect 217179 305628 217180 305692
rect 217244 305628 217245 305692
rect 217179 305627 217245 305628
rect 217182 158133 217242 305627
rect 217179 158132 217245 158133
rect 217179 158068 217180 158132
rect 217244 158068 217245 158132
rect 217179 158067 217245 158068
rect 216995 157996 217061 157997
rect 216995 157932 216996 157996
rect 217060 157932 217061 157996
rect 216995 157931 217061 157932
rect 217366 157861 217426 308619
rect 217547 308548 217613 308549
rect 217547 308484 217548 308548
rect 217612 308484 217613 308548
rect 217547 308483 217613 308484
rect 217550 158405 217610 308483
rect 217794 291454 218414 326898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 219019 308956 219085 308957
rect 219019 308892 219020 308956
rect 219084 308892 219085 308956
rect 219019 308891 219085 308892
rect 218835 308820 218901 308821
rect 218835 308756 218836 308820
rect 218900 308756 218901 308820
rect 218835 308755 218901 308756
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 245308 218414 254898
rect 218651 243540 218717 243541
rect 218651 243476 218652 243540
rect 218716 243476 218717 243540
rect 218651 243475 218717 243476
rect 217547 158404 217613 158405
rect 217547 158340 217548 158404
rect 217612 158340 217613 158404
rect 217547 158339 217613 158340
rect 217363 157860 217429 157861
rect 217363 157796 217364 157860
rect 217428 157796 217429 157860
rect 217363 157795 217429 157796
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 215155 3500 215221 3501
rect 215155 3436 215156 3500
rect 215220 3436 215221 3500
rect 215155 3435 215221 3436
rect 216443 3500 216509 3501
rect 216443 3436 216444 3500
rect 216508 3436 216509 3500
rect 216443 3435 216509 3436
rect 217794 3454 218414 38898
rect 218654 3637 218714 243475
rect 218838 158541 218898 308755
rect 219022 158677 219082 308891
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 219203 262852 219269 262853
rect 219203 262788 219204 262852
rect 219268 262788 219269 262852
rect 219203 262787 219269 262788
rect 219019 158676 219085 158677
rect 219019 158612 219020 158676
rect 219084 158612 219085 158676
rect 219019 158611 219085 158612
rect 218835 158540 218901 158541
rect 218835 158476 218836 158540
rect 218900 158476 218901 158540
rect 218835 158475 218901 158476
rect 218651 3636 218717 3637
rect 218651 3572 218652 3636
rect 218716 3572 218717 3636
rect 218651 3571 218717 3572
rect 219206 3501 219266 262787
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 235950 476237 236010 479710
rect 237238 476237 237298 479710
rect 238158 479710 238292 479770
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 238158 476373 238218 479710
rect 238155 476372 238221 476373
rect 238155 476308 238156 476372
rect 238220 476308 238221 476372
rect 238155 476307 238221 476308
rect 239630 476237 239690 479710
rect 240550 476237 240610 479710
rect 241838 476237 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 243126 476373 243186 479710
rect 244230 476509 244290 479710
rect 245334 479710 245500 479770
rect 246438 479710 246588 479770
rect 247542 479710 247676 479770
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 250064 479710 250178 479770
rect 244227 476508 244293 476509
rect 244227 476444 244228 476508
rect 244292 476444 244293 476508
rect 244227 476443 244293 476444
rect 245334 476373 245394 479710
rect 243123 476372 243189 476373
rect 243123 476308 243124 476372
rect 243188 476308 243189 476372
rect 243123 476307 243189 476308
rect 245331 476372 245397 476373
rect 245331 476308 245332 476372
rect 245396 476308 245397 476372
rect 245331 476307 245397 476308
rect 246438 476237 246498 479710
rect 247542 476237 247602 479710
rect 248278 476645 248338 479710
rect 248275 476644 248341 476645
rect 248275 476580 248276 476644
rect 248340 476580 248341 476644
rect 248275 476579 248341 476580
rect 248646 476237 248706 479710
rect 250118 476237 250178 479710
rect 250670 479710 250804 479770
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 251288 479710 251466 479770
rect 250670 476645 250730 479710
rect 250667 476644 250733 476645
rect 250667 476580 250668 476644
rect 250732 476580 250733 476644
rect 250667 476579 250733 476580
rect 251406 476373 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 251403 476372 251469 476373
rect 251403 476308 251404 476372
rect 251468 476308 251469 476372
rect 251403 476307 251469 476308
rect 252326 476237 252386 479710
rect 253430 476917 253490 479710
rect 253427 476916 253493 476917
rect 253427 476852 253428 476916
rect 253492 476852 253493 476916
rect 253427 476851 253493 476852
rect 253614 476645 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 258496 479770 258556 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 253611 476644 253677 476645
rect 253611 476580 253612 476644
rect 253676 476580 253677 476644
rect 253611 476579 253677 476580
rect 254534 476237 254594 479710
rect 255822 476917 255882 479710
rect 255819 476916 255885 476917
rect 255819 476852 255820 476916
rect 255884 476852 255885 476916
rect 255819 476851 255885 476852
rect 256190 476781 256250 479710
rect 256187 476780 256253 476781
rect 256187 476716 256188 476780
rect 256252 476716 256253 476780
rect 256187 476715 256253 476716
rect 257110 476373 257170 479710
rect 257846 479710 258148 479770
rect 258398 479710 258556 479770
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 259448 479710 259562 479770
rect 257107 476372 257173 476373
rect 257107 476308 257108 476372
rect 257172 476308 257173 476372
rect 257846 476370 257906 479710
rect 258398 476373 258458 479710
rect 258395 476372 258461 476373
rect 257846 476310 258090 476370
rect 257107 476307 257173 476308
rect 258030 476237 258090 476310
rect 258395 476308 258396 476372
rect 258460 476308 258461 476372
rect 258395 476307 258461 476308
rect 259502 476237 259562 479710
rect 260606 479710 260732 479770
rect 260974 479710 261140 479770
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 260606 476509 260666 479710
rect 260603 476508 260669 476509
rect 260603 476444 260604 476508
rect 260668 476444 260669 476508
rect 260603 476443 260669 476444
rect 260974 476373 261034 479710
rect 260971 476372 261037 476373
rect 260971 476308 260972 476372
rect 261036 476308 261037 476372
rect 260971 476307 261037 476308
rect 261710 476237 261770 479710
rect 262814 476237 262874 479710
rect 263550 476645 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476644 263613 476645
rect 263547 476580 263548 476644
rect 263612 476580 263613 476644
rect 263547 476579 263613 476580
rect 263918 476237 263978 479710
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 476645 266002 479710
rect 265939 476644 266005 476645
rect 265939 476580 265940 476644
rect 266004 476580 266005 476644
rect 265939 476579 266005 476580
rect 266494 476373 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 266491 476372 266557 476373
rect 266491 476308 266492 476372
rect 266556 476308 266557 476372
rect 266491 476307 266557 476308
rect 267598 476237 267658 479710
rect 268334 476509 268394 479710
rect 268331 476508 268397 476509
rect 268331 476444 268332 476508
rect 268396 476444 268397 476508
rect 268331 476443 268397 476444
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 271144 479710 271338 479770
rect 270910 476917 270970 479710
rect 270907 476916 270973 476917
rect 270907 476852 270908 476916
rect 270972 476852 270973 476916
rect 270907 476851 270973 476852
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273486 479710 273652 479770
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 272198 476645 272258 479710
rect 272195 476644 272261 476645
rect 272195 476580 272196 476644
rect 272260 476580 272261 476644
rect 272195 476579 272261 476580
rect 273302 476373 273362 479710
rect 273486 476509 273546 479710
rect 273483 476508 273549 476509
rect 273483 476444 273484 476508
rect 273548 476444 273549 476508
rect 273483 476443 273549 476444
rect 273299 476372 273365 476373
rect 273299 476308 273300 476372
rect 273364 476308 273365 476372
rect 273299 476307 273365 476308
rect 274406 476237 274466 479710
rect 275878 476237 275938 479710
rect 276062 476373 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476372 276125 476373
rect 276059 476308 276060 476372
rect 276124 476308 276125 476372
rect 276059 476307 276125 476308
rect 276982 476237 277042 479710
rect 278086 476237 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 279168 479710 279250 479770
rect 278454 477053 278514 479710
rect 278451 477052 278517 477053
rect 278451 476988 278452 477052
rect 278516 476988 278517 477052
rect 278451 476987 278517 476988
rect 279190 476237 279250 479710
rect 280846 479710 280996 479770
rect 283422 479710 283580 479770
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 293448 479770 293508 480080
rect 285968 479710 286058 479770
rect 280846 476373 280906 479710
rect 280843 476372 280909 476373
rect 280843 476308 280844 476372
rect 280908 476308 280909 476372
rect 280843 476307 280909 476308
rect 283422 476237 283482 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293358 479710 293508 479770
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293358 476237 293418 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305870 479710 306020 479770
rect 308446 479710 308604 479770
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 318472 479770 318532 480080
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476781 303538 479710
rect 305870 477053 305930 479710
rect 308446 477053 308506 479710
rect 305867 477052 305933 477053
rect 305867 476988 305868 477052
rect 305932 476988 305933 477052
rect 305867 476987 305933 476988
rect 308443 477052 308509 477053
rect 308443 476988 308444 477052
rect 308508 476988 308509 477052
rect 308443 476987 308509 476988
rect 311022 476917 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318382 479710 318532 479770
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 320920 479710 321018 479770
rect 311019 476916 311085 476917
rect 311019 476852 311020 476916
rect 311084 476852 311085 476916
rect 311019 476851 311085 476852
rect 303475 476780 303541 476781
rect 303475 476716 303476 476780
rect 303540 476716 303541 476780
rect 303475 476715 303541 476716
rect 313414 476509 313474 479710
rect 315806 476509 315866 479710
rect 313411 476508 313477 476509
rect 313411 476444 313412 476508
rect 313476 476444 313477 476508
rect 313411 476443 313477 476444
rect 315803 476508 315869 476509
rect 315803 476444 315804 476508
rect 315868 476444 315869 476508
rect 315803 476443 315869 476444
rect 318382 476373 318442 479710
rect 320958 476373 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 476917 323410 479710
rect 323347 476916 323413 476917
rect 323347 476852 323348 476916
rect 323412 476852 323413 476916
rect 323347 476851 323413 476852
rect 318379 476372 318445 476373
rect 318379 476308 318380 476372
rect 318444 476308 318445 476372
rect 318379 476307 318445 476308
rect 320955 476372 321021 476373
rect 320955 476308 320956 476372
rect 321020 476308 321021 476372
rect 320955 476307 321021 476308
rect 325926 476237 325986 479710
rect 235947 476236 236013 476237
rect 235947 476172 235948 476236
rect 236012 476172 236013 476236
rect 235947 476171 236013 476172
rect 237235 476236 237301 476237
rect 237235 476172 237236 476236
rect 237300 476172 237301 476236
rect 237235 476171 237301 476172
rect 239627 476236 239693 476237
rect 239627 476172 239628 476236
rect 239692 476172 239693 476236
rect 239627 476171 239693 476172
rect 240547 476236 240613 476237
rect 240547 476172 240548 476236
rect 240612 476172 240613 476236
rect 240547 476171 240613 476172
rect 241835 476236 241901 476237
rect 241835 476172 241836 476236
rect 241900 476172 241901 476236
rect 241835 476171 241901 476172
rect 246435 476236 246501 476237
rect 246435 476172 246436 476236
rect 246500 476172 246501 476236
rect 246435 476171 246501 476172
rect 247539 476236 247605 476237
rect 247539 476172 247540 476236
rect 247604 476172 247605 476236
rect 247539 476171 247605 476172
rect 248643 476236 248709 476237
rect 248643 476172 248644 476236
rect 248708 476172 248709 476236
rect 248643 476171 248709 476172
rect 250115 476236 250181 476237
rect 250115 476172 250116 476236
rect 250180 476172 250181 476236
rect 250115 476171 250181 476172
rect 252323 476236 252389 476237
rect 252323 476172 252324 476236
rect 252388 476172 252389 476236
rect 252323 476171 252389 476172
rect 254531 476236 254597 476237
rect 254531 476172 254532 476236
rect 254596 476172 254597 476236
rect 254531 476171 254597 476172
rect 258027 476236 258093 476237
rect 258027 476172 258028 476236
rect 258092 476172 258093 476236
rect 258027 476171 258093 476172
rect 259499 476236 259565 476237
rect 259499 476172 259500 476236
rect 259564 476172 259565 476236
rect 259499 476171 259565 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 262811 476236 262877 476237
rect 262811 476172 262812 476236
rect 262876 476172 262877 476236
rect 262811 476171 262877 476172
rect 263915 476236 263981 476237
rect 263915 476172 263916 476236
rect 263980 476172 263981 476236
rect 263915 476171 263981 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 267595 476236 267661 476237
rect 267595 476172 267596 476236
rect 267660 476172 267661 476236
rect 267595 476171 267661 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 274403 476236 274469 476237
rect 274403 476172 274404 476236
rect 274468 476172 274469 476236
rect 274403 476171 274469 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278083 476236 278149 476237
rect 278083 476172 278084 476236
rect 278148 476172 278149 476236
rect 278083 476171 278149 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 283419 476236 283485 476237
rect 283419 476172 283420 476236
rect 283484 476172 283485 476236
rect 283419 476171 283485 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293355 476236 293421 476237
rect 293355 476172 293356 476236
rect 293420 476172 293421 476236
rect 293355 476171 293421 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 325923 476236 325989 476237
rect 325923 476172 325924 476236
rect 325988 476172 325989 476236
rect 325923 476171 325989 476172
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 444835 362414 470898
rect 366294 706108 366914 711900
rect 366294 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 366914 706108
rect 366294 705788 366914 705872
rect 366294 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 366914 705788
rect 366294 691954 366914 705552
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 363459 443324 363525 443325
rect 363459 443260 363460 443324
rect 363524 443260 363525 443324
rect 363459 443259 363525 443260
rect 360331 442236 360397 442237
rect 360331 442172 360332 442236
rect 360396 442172 360397 442236
rect 360331 442171 360397 442172
rect 361619 442236 361685 442237
rect 361619 442172 361620 442236
rect 361684 442172 361685 442236
rect 361619 442171 361685 442172
rect 251968 439954 252288 439986
rect 251968 439718 252010 439954
rect 252246 439718 252288 439954
rect 251968 439634 252288 439718
rect 251968 439398 252010 439634
rect 252246 439398 252288 439634
rect 251968 439366 252288 439398
rect 282688 439954 283008 439986
rect 282688 439718 282730 439954
rect 282966 439718 283008 439954
rect 282688 439634 283008 439718
rect 282688 439398 282730 439634
rect 282966 439398 283008 439634
rect 282688 439366 283008 439398
rect 313408 439954 313728 439986
rect 313408 439718 313450 439954
rect 313686 439718 313728 439954
rect 313408 439634 313728 439718
rect 313408 439398 313450 439634
rect 313686 439398 313728 439634
rect 313408 439366 313728 439398
rect 344128 439954 344448 439986
rect 344128 439718 344170 439954
rect 344406 439718 344448 439954
rect 344128 439634 344448 439718
rect 344128 439398 344170 439634
rect 344406 439398 344448 439634
rect 344128 439366 344448 439398
rect 236608 435454 236928 435486
rect 236608 435218 236650 435454
rect 236886 435218 236928 435454
rect 236608 435134 236928 435218
rect 236608 434898 236650 435134
rect 236886 434898 236928 435134
rect 236608 434866 236928 434898
rect 267328 435454 267648 435486
rect 267328 435218 267370 435454
rect 267606 435218 267648 435454
rect 267328 435134 267648 435218
rect 267328 434898 267370 435134
rect 267606 434898 267648 435134
rect 267328 434866 267648 434898
rect 298048 435454 298368 435486
rect 298048 435218 298090 435454
rect 298326 435218 298368 435454
rect 298048 435134 298368 435218
rect 298048 434898 298090 435134
rect 298326 434898 298368 435134
rect 298048 434866 298368 434898
rect 328768 435454 329088 435486
rect 328768 435218 328810 435454
rect 329046 435218 329088 435454
rect 328768 435134 329088 435218
rect 328768 434898 328810 435134
rect 329046 434898 329088 435134
rect 328768 434866 329088 434898
rect 359488 435454 359808 435486
rect 359488 435218 359530 435454
rect 359766 435218 359808 435454
rect 359488 435134 359808 435218
rect 359488 434898 359530 435134
rect 359766 434898 359808 435134
rect 359488 434866 359808 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 251968 403954 252288 403986
rect 251968 403718 252010 403954
rect 252246 403718 252288 403954
rect 251968 403634 252288 403718
rect 251968 403398 252010 403634
rect 252246 403398 252288 403634
rect 251968 403366 252288 403398
rect 282688 403954 283008 403986
rect 282688 403718 282730 403954
rect 282966 403718 283008 403954
rect 282688 403634 283008 403718
rect 282688 403398 282730 403634
rect 282966 403398 283008 403634
rect 282688 403366 283008 403398
rect 313408 403954 313728 403986
rect 313408 403718 313450 403954
rect 313686 403718 313728 403954
rect 313408 403634 313728 403718
rect 313408 403398 313450 403634
rect 313686 403398 313728 403634
rect 313408 403366 313728 403398
rect 344128 403954 344448 403986
rect 344128 403718 344170 403954
rect 344406 403718 344448 403954
rect 344128 403634 344448 403718
rect 344128 403398 344170 403634
rect 344406 403398 344448 403634
rect 344128 403366 344448 403398
rect 236608 399454 236928 399486
rect 236608 399218 236650 399454
rect 236886 399218 236928 399454
rect 236608 399134 236928 399218
rect 236608 398898 236650 399134
rect 236886 398898 236928 399134
rect 236608 398866 236928 398898
rect 267328 399454 267648 399486
rect 267328 399218 267370 399454
rect 267606 399218 267648 399454
rect 267328 399134 267648 399218
rect 267328 398898 267370 399134
rect 267606 398898 267648 399134
rect 267328 398866 267648 398898
rect 298048 399454 298368 399486
rect 298048 399218 298090 399454
rect 298326 399218 298368 399454
rect 298048 399134 298368 399218
rect 298048 398898 298090 399134
rect 298326 398898 298368 399134
rect 298048 398866 298368 398898
rect 328768 399454 329088 399486
rect 328768 399218 328810 399454
rect 329046 399218 329088 399454
rect 328768 399134 329088 399218
rect 328768 398898 328810 399134
rect 329046 398898 329088 399134
rect 328768 398866 329088 398898
rect 359488 399454 359808 399486
rect 359488 399218 359530 399454
rect 359766 399218 359808 399454
rect 359488 399134 359808 399218
rect 359488 398898 359530 399134
rect 359766 398898 359808 399134
rect 359488 398866 359808 398898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 251968 367954 252288 367986
rect 251968 367718 252010 367954
rect 252246 367718 252288 367954
rect 251968 367634 252288 367718
rect 251968 367398 252010 367634
rect 252246 367398 252288 367634
rect 251968 367366 252288 367398
rect 282688 367954 283008 367986
rect 282688 367718 282730 367954
rect 282966 367718 283008 367954
rect 282688 367634 283008 367718
rect 282688 367398 282730 367634
rect 282966 367398 283008 367634
rect 282688 367366 283008 367398
rect 313408 367954 313728 367986
rect 313408 367718 313450 367954
rect 313686 367718 313728 367954
rect 313408 367634 313728 367718
rect 313408 367398 313450 367634
rect 313686 367398 313728 367634
rect 313408 367366 313728 367398
rect 344128 367954 344448 367986
rect 344128 367718 344170 367954
rect 344406 367718 344448 367954
rect 344128 367634 344448 367718
rect 344128 367398 344170 367634
rect 344406 367398 344448 367634
rect 344128 367366 344448 367398
rect 236608 363454 236928 363486
rect 236608 363218 236650 363454
rect 236886 363218 236928 363454
rect 236608 363134 236928 363218
rect 236608 362898 236650 363134
rect 236886 362898 236928 363134
rect 236608 362866 236928 362898
rect 267328 363454 267648 363486
rect 267328 363218 267370 363454
rect 267606 363218 267648 363454
rect 267328 363134 267648 363218
rect 267328 362898 267370 363134
rect 267606 362898 267648 363134
rect 267328 362866 267648 362898
rect 298048 363454 298368 363486
rect 298048 363218 298090 363454
rect 298326 363218 298368 363454
rect 298048 363134 298368 363218
rect 298048 362898 298090 363134
rect 298326 362898 298368 363134
rect 298048 362866 298368 362898
rect 328768 363454 329088 363486
rect 328768 363218 328810 363454
rect 329046 363218 329088 363454
rect 328768 363134 329088 363218
rect 328768 362898 328810 363134
rect 329046 362898 329088 363134
rect 328768 362866 329088 362898
rect 359488 363454 359808 363486
rect 359488 363218 359530 363454
rect 359766 363218 359808 363454
rect 359488 363134 359808 363218
rect 359488 362898 359530 363134
rect 359766 362898 359808 363134
rect 359488 362866 359808 362898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 251968 331954 252288 331986
rect 251968 331718 252010 331954
rect 252246 331718 252288 331954
rect 251968 331634 252288 331718
rect 251968 331398 252010 331634
rect 252246 331398 252288 331634
rect 251968 331366 252288 331398
rect 282688 331954 283008 331986
rect 282688 331718 282730 331954
rect 282966 331718 283008 331954
rect 282688 331634 283008 331718
rect 282688 331398 282730 331634
rect 282966 331398 283008 331634
rect 282688 331366 283008 331398
rect 313408 331954 313728 331986
rect 313408 331718 313450 331954
rect 313686 331718 313728 331954
rect 313408 331634 313728 331718
rect 313408 331398 313450 331634
rect 313686 331398 313728 331634
rect 313408 331366 313728 331398
rect 344128 331954 344448 331986
rect 344128 331718 344170 331954
rect 344406 331718 344448 331954
rect 344128 331634 344448 331718
rect 344128 331398 344170 331634
rect 344406 331398 344448 331634
rect 344128 331366 344448 331398
rect 236608 327454 236928 327486
rect 236608 327218 236650 327454
rect 236886 327218 236928 327454
rect 236608 327134 236928 327218
rect 236608 326898 236650 327134
rect 236886 326898 236928 327134
rect 236608 326866 236928 326898
rect 267328 327454 267648 327486
rect 267328 327218 267370 327454
rect 267606 327218 267648 327454
rect 267328 327134 267648 327218
rect 267328 326898 267370 327134
rect 267606 326898 267648 327134
rect 267328 326866 267648 326898
rect 298048 327454 298368 327486
rect 298048 327218 298090 327454
rect 298326 327218 298368 327454
rect 298048 327134 298368 327218
rect 298048 326898 298090 327134
rect 298326 326898 298368 327134
rect 298048 326866 298368 326898
rect 328768 327454 329088 327486
rect 328768 327218 328810 327454
rect 329046 327218 329088 327454
rect 328768 327134 329088 327218
rect 328768 326898 328810 327134
rect 329046 326898 329088 327134
rect 328768 326866 329088 326898
rect 359488 327454 359808 327486
rect 359488 327218 359530 327454
rect 359766 327218 359808 327454
rect 359488 327134 359808 327218
rect 359488 326898 359530 327134
rect 359766 326898 359808 327134
rect 359488 326866 359808 326898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 245308 245414 245898
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 245308 249914 250398
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 245308 254414 254898
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 245308 258914 259398
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 245308 263414 263898
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 245308 267914 268398
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 245308 281414 245898
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 245308 285914 250398
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 245308 290414 254898
rect 294294 295954 294914 308400
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 245308 294914 259398
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 358859 264212 358925 264213
rect 358859 264148 358860 264212
rect 358924 264148 358925 264212
rect 358859 264147 358925 264148
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 358123 245580 358189 245581
rect 358123 245516 358124 245580
rect 358188 245516 358189 245580
rect 358123 245515 358189 245516
rect 357571 244764 357637 244765
rect 357571 244700 357572 244764
rect 357636 244700 357637 244764
rect 357571 244699 357637 244700
rect 220272 223954 220620 223986
rect 220272 223718 220328 223954
rect 220564 223718 220620 223954
rect 220272 223634 220620 223718
rect 220272 223398 220328 223634
rect 220564 223398 220620 223634
rect 220272 223366 220620 223398
rect 356000 223954 356348 223986
rect 356000 223718 356056 223954
rect 356292 223718 356348 223954
rect 356000 223634 356348 223718
rect 356000 223398 356056 223634
rect 356292 223398 356348 223634
rect 356000 223366 356348 223398
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 187954 220620 187986
rect 220272 187718 220328 187954
rect 220564 187718 220620 187954
rect 220272 187634 220620 187718
rect 220272 187398 220328 187634
rect 220564 187398 220620 187634
rect 220272 187366 220620 187398
rect 356000 187954 356348 187986
rect 356000 187718 356056 187954
rect 356292 187718 356348 187954
rect 356000 187634 356348 187718
rect 356000 187398 356056 187634
rect 356292 187398 356348 187634
rect 356000 187366 356348 187398
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 159490 236116 160106
rect 237144 159490 237204 160106
rect 238232 159490 238292 160106
rect 236056 159430 236562 159490
rect 237144 159430 237298 159490
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 214419 3364 214485 3365
rect 214419 3300 214420 3364
rect 214484 3300 214485 3364
rect 214419 3299 214485 3300
rect 213294 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 213914 -7376
rect 213294 -7696 213914 -7612
rect 213294 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 213914 -7696
rect 213294 -7964 213914 -7932
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 219203 3500 219269 3501
rect 219203 3436 219204 3500
rect 219268 3436 219269 3500
rect 219203 3435 219269 3436
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -656 218414 2898
rect 217794 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 218414 -656
rect 217794 -976 218414 -892
rect 217794 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 218414 -976
rect 217794 -7964 218414 -1212
rect 222294 -1616 222914 7398
rect 222294 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 222914 -1616
rect 222294 -1936 222914 -1852
rect 222294 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 222914 -1936
rect 222294 -7964 222914 -2172
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2576 227414 11898
rect 226794 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 227414 -2576
rect 226794 -2896 227414 -2812
rect 226794 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 227414 -2896
rect 226794 -7964 227414 -3132
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3536 231914 16398
rect 231294 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 231914 -3536
rect 231294 -3856 231914 -3772
rect 231294 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 231914 -3856
rect 231294 -7964 231914 -4092
rect 235794 129454 236414 158000
rect 236502 157453 236562 159430
rect 237238 158541 237298 159430
rect 238158 159430 238292 159490
rect 239592 159490 239652 160106
rect 240544 159490 240604 160106
rect 241768 159490 241828 160106
rect 243128 159490 243188 160106
rect 239592 159430 239690 159490
rect 240544 159430 240610 159490
rect 241768 159430 241898 159490
rect 238158 158677 238218 159430
rect 239630 158677 239690 159430
rect 238155 158676 238221 158677
rect 238155 158612 238156 158676
rect 238220 158612 238221 158676
rect 238155 158611 238221 158612
rect 239627 158676 239693 158677
rect 239627 158612 239628 158676
rect 239692 158612 239693 158676
rect 239627 158611 239693 158612
rect 237235 158540 237301 158541
rect 237235 158476 237236 158540
rect 237300 158476 237301 158540
rect 237235 158475 237301 158476
rect 240550 158405 240610 159430
rect 241838 158677 241898 159430
rect 243126 159430 243188 159490
rect 244216 159490 244276 160106
rect 245440 159490 245500 160106
rect 246528 159490 246588 160106
rect 247616 159490 247676 160106
rect 248296 159490 248356 160106
rect 248704 159490 248764 160106
rect 244216 159430 244290 159490
rect 245440 159430 245578 159490
rect 246528 159430 246682 159490
rect 247616 159430 247786 159490
rect 243126 158813 243186 159430
rect 243123 158812 243189 158813
rect 243123 158748 243124 158812
rect 243188 158748 243189 158812
rect 243123 158747 243189 158748
rect 244230 158677 244290 159430
rect 241835 158676 241901 158677
rect 241835 158612 241836 158676
rect 241900 158612 241901 158676
rect 241835 158611 241901 158612
rect 244227 158676 244293 158677
rect 244227 158612 244228 158676
rect 244292 158612 244293 158676
rect 244227 158611 244293 158612
rect 240547 158404 240613 158405
rect 240547 158340 240548 158404
rect 240612 158340 240613 158404
rect 240547 158339 240613 158340
rect 236499 157452 236565 157453
rect 236499 157388 236500 157452
rect 236564 157388 236565 157452
rect 236499 157387 236565 157388
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4496 236414 20898
rect 235794 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 236414 -4496
rect 235794 -4816 236414 -4732
rect 235794 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 236414 -4816
rect 235794 -7964 236414 -5052
rect 240294 133954 240914 158000
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5456 240914 25398
rect 240294 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 240914 -5456
rect 240294 -5776 240914 -5692
rect 240294 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 240914 -5776
rect 240294 -7964 240914 -6012
rect 244794 138454 245414 158000
rect 245518 157861 245578 159430
rect 246622 158133 246682 159430
rect 246619 158132 246685 158133
rect 246619 158068 246620 158132
rect 246684 158068 246685 158132
rect 246619 158067 246685 158068
rect 247726 157861 247786 159430
rect 248278 159430 248356 159490
rect 248646 159430 248764 159490
rect 250064 159490 250124 160106
rect 250744 159490 250804 160106
rect 251288 159490 251348 160106
rect 252376 159490 252436 160106
rect 253464 159490 253524 160106
rect 250064 159430 250178 159490
rect 250744 159430 250914 159490
rect 251288 159430 251466 159490
rect 248278 158677 248338 159430
rect 248275 158676 248341 158677
rect 248275 158612 248276 158676
rect 248340 158612 248341 158676
rect 248275 158611 248341 158612
rect 248646 157861 248706 159430
rect 245515 157860 245581 157861
rect 245515 157796 245516 157860
rect 245580 157796 245581 157860
rect 245515 157795 245581 157796
rect 247723 157860 247789 157861
rect 247723 157796 247724 157860
rect 247788 157796 247789 157860
rect 247723 157795 247789 157796
rect 248643 157860 248709 157861
rect 248643 157796 248644 157860
rect 248708 157796 248709 157860
rect 248643 157795 248709 157796
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6416 245414 29898
rect 244794 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 245414 -6416
rect 244794 -6736 245414 -6652
rect 244794 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 245414 -6736
rect 244794 -7964 245414 -6972
rect 249294 142954 249914 158000
rect 250118 157861 250178 159430
rect 250854 158677 250914 159430
rect 251406 158677 251466 159430
rect 252326 159430 252436 159490
rect 253430 159430 253524 159490
rect 253600 159490 253660 160106
rect 254552 159490 254612 160106
rect 253600 159430 253674 159490
rect 250851 158676 250917 158677
rect 250851 158612 250852 158676
rect 250916 158612 250917 158676
rect 250851 158611 250917 158612
rect 251403 158676 251469 158677
rect 251403 158612 251404 158676
rect 251468 158612 251469 158676
rect 251403 158611 251469 158612
rect 252326 158405 252386 159430
rect 252323 158404 252389 158405
rect 252323 158340 252324 158404
rect 252388 158340 252389 158404
rect 252323 158339 252389 158340
rect 253430 157861 253490 159430
rect 253614 158949 253674 159430
rect 254534 159430 254612 159490
rect 255912 159490 255972 160106
rect 256048 159629 256108 160106
rect 256045 159628 256111 159629
rect 256045 159564 256046 159628
rect 256110 159564 256111 159628
rect 256045 159563 256111 159564
rect 257000 159490 257060 160106
rect 258088 159490 258148 160106
rect 258496 159490 258556 160106
rect 259448 159490 259508 160106
rect 260672 159490 260732 160106
rect 261080 159490 261140 160106
rect 261760 159490 261820 160106
rect 262848 159490 262908 160106
rect 255912 159430 256066 159490
rect 257000 159430 257170 159490
rect 258088 159430 258274 159490
rect 258496 159430 258642 159490
rect 259448 159430 259562 159490
rect 260672 159430 260850 159490
rect 261080 159430 261218 159490
rect 253611 158948 253677 158949
rect 253611 158884 253612 158948
rect 253676 158884 253677 158948
rect 253611 158883 253677 158884
rect 254534 158133 254594 159430
rect 256006 159085 256066 159430
rect 256003 159084 256069 159085
rect 256003 159020 256004 159084
rect 256068 159020 256069 159084
rect 256003 159019 256069 159020
rect 257110 158677 257170 159430
rect 258214 159221 258274 159430
rect 258211 159220 258277 159221
rect 258211 159156 258212 159220
rect 258276 159156 258277 159220
rect 258211 159155 258277 159156
rect 257107 158676 257173 158677
rect 257107 158612 257108 158676
rect 257172 158612 257173 158676
rect 257107 158611 257173 158612
rect 258582 158269 258642 159430
rect 259502 158677 259562 159430
rect 259499 158676 259565 158677
rect 259499 158612 259500 158676
rect 259564 158612 259565 158676
rect 259499 158611 259565 158612
rect 258579 158268 258645 158269
rect 258579 158204 258580 158268
rect 258644 158204 258645 158268
rect 258579 158203 258645 158204
rect 254531 158132 254597 158133
rect 254531 158068 254532 158132
rect 254596 158068 254597 158132
rect 254531 158067 254597 158068
rect 250115 157860 250181 157861
rect 250115 157796 250116 157860
rect 250180 157796 250181 157860
rect 250115 157795 250181 157796
rect 253427 157860 253493 157861
rect 253427 157796 253428 157860
rect 253492 157796 253493 157860
rect 253427 157795 253493 157796
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7376 249914 34398
rect 249294 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 249914 -7376
rect 249294 -7696 249914 -7612
rect 249294 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 249914 -7696
rect 249294 -7964 249914 -7932
rect 253794 147454 254414 158000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -656 254414 2898
rect 253794 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 254414 -656
rect 253794 -976 254414 -892
rect 253794 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 254414 -976
rect 253794 -7964 254414 -1212
rect 258294 151954 258914 158000
rect 260790 157997 260850 159430
rect 260787 157996 260853 157997
rect 260787 157932 260788 157996
rect 260852 157932 260853 157996
rect 260787 157931 260853 157932
rect 261158 157589 261218 159430
rect 261710 159430 261820 159490
rect 262814 159430 262908 159490
rect 263528 159490 263588 160106
rect 263936 159490 263996 160106
rect 263528 159430 263610 159490
rect 261710 158677 261770 159430
rect 262814 159357 262874 159430
rect 262811 159356 262877 159357
rect 262811 159292 262812 159356
rect 262876 159292 262877 159356
rect 262811 159291 262877 159292
rect 261707 158676 261773 158677
rect 261707 158612 261708 158676
rect 261772 158612 261773 158676
rect 261707 158611 261773 158612
rect 261155 157588 261221 157589
rect 261155 157524 261156 157588
rect 261220 157524 261221 157588
rect 261155 157523 261221 157524
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1616 258914 7398
rect 258294 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 258914 -1616
rect 258294 -1936 258914 -1852
rect 258294 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 258914 -1936
rect 258294 -7964 258914 -2172
rect 262794 156454 263414 158000
rect 263550 157589 263610 159430
rect 263918 159430 263996 159490
rect 265296 159490 265356 160106
rect 265976 159490 266036 160106
rect 265296 159430 265450 159490
rect 263918 158677 263978 159430
rect 265390 158677 265450 159430
rect 265942 159430 266036 159490
rect 266384 159490 266444 160106
rect 267608 159490 267668 160106
rect 266384 159430 266554 159490
rect 263915 158676 263981 158677
rect 263915 158612 263916 158676
rect 263980 158612 263981 158676
rect 263915 158611 263981 158612
rect 265387 158676 265453 158677
rect 265387 158612 265388 158676
rect 265452 158612 265453 158676
rect 265387 158611 265453 158612
rect 265942 157589 266002 159430
rect 266494 157725 266554 159430
rect 267046 159430 267668 159490
rect 268288 159490 268348 160106
rect 268696 159490 268756 160106
rect 269784 159490 269844 160106
rect 271008 159629 271068 160106
rect 271005 159628 271071 159629
rect 271005 159564 271006 159628
rect 271070 159564 271071 159628
rect 271005 159563 271071 159564
rect 271144 159490 271204 160106
rect 272232 159490 272292 160106
rect 273320 159490 273380 160106
rect 268288 159430 268394 159490
rect 268696 159430 268762 159490
rect 269784 159430 269866 159490
rect 267046 157861 267106 159430
rect 268334 158677 268394 159430
rect 268702 158677 268762 159430
rect 269806 158677 269866 159430
rect 271094 159430 271204 159490
rect 272198 159430 272292 159490
rect 273302 159430 273380 159490
rect 273592 159490 273652 160106
rect 274408 159490 274468 160106
rect 275768 159629 275828 160106
rect 275765 159628 275831 159629
rect 275765 159564 275766 159628
rect 275830 159564 275831 159628
rect 275765 159563 275831 159564
rect 273592 159430 273730 159490
rect 271094 158677 271154 159430
rect 272198 158677 272258 159430
rect 273302 158677 273362 159430
rect 268331 158676 268397 158677
rect 268331 158612 268332 158676
rect 268396 158612 268397 158676
rect 268331 158611 268397 158612
rect 268699 158676 268765 158677
rect 268699 158612 268700 158676
rect 268764 158612 268765 158676
rect 268699 158611 268765 158612
rect 269803 158676 269869 158677
rect 269803 158612 269804 158676
rect 269868 158612 269869 158676
rect 269803 158611 269869 158612
rect 271091 158676 271157 158677
rect 271091 158612 271092 158676
rect 271156 158612 271157 158676
rect 271091 158611 271157 158612
rect 272195 158676 272261 158677
rect 272195 158612 272196 158676
rect 272260 158612 272261 158676
rect 272195 158611 272261 158612
rect 273299 158676 273365 158677
rect 273299 158612 273300 158676
rect 273364 158612 273365 158676
rect 273299 158611 273365 158612
rect 267043 157860 267109 157861
rect 267043 157796 267044 157860
rect 267108 157796 267109 157860
rect 267043 157795 267109 157796
rect 266491 157724 266557 157725
rect 266491 157660 266492 157724
rect 266556 157660 266557 157724
rect 266491 157659 266557 157660
rect 263547 157588 263613 157589
rect 263547 157524 263548 157588
rect 263612 157524 263613 157588
rect 263547 157523 263613 157524
rect 265939 157588 266005 157589
rect 265939 157524 265940 157588
rect 266004 157524 266005 157588
rect 265939 157523 266005 157524
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2576 263414 11898
rect 262794 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 263414 -2576
rect 262794 -2896 263414 -2812
rect 262794 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 263414 -2896
rect 262794 -7964 263414 -3132
rect 267294 124954 267914 158000
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3536 267914 16398
rect 267294 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 267914 -3536
rect 267294 -3856 267914 -3772
rect 267294 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 267914 -3856
rect 267294 -7964 267914 -4092
rect 271794 129454 272414 158000
rect 273670 157725 273730 159430
rect 274406 159430 274468 159490
rect 276040 159490 276100 160106
rect 276992 159901 277052 160106
rect 278080 159901 278140 160106
rect 276989 159900 277055 159901
rect 276989 159836 276990 159900
rect 277054 159836 277055 159900
rect 276989 159835 277055 159836
rect 278077 159900 278143 159901
rect 278077 159836 278078 159900
rect 278142 159836 278143 159900
rect 278488 159898 278548 160106
rect 279168 159901 279228 160106
rect 278077 159835 278143 159836
rect 278454 159838 278548 159898
rect 279165 159900 279231 159901
rect 276040 159430 276122 159490
rect 274406 158677 274466 159430
rect 276062 158677 276122 159430
rect 274403 158676 274469 158677
rect 274403 158612 274404 158676
rect 274468 158612 274469 158676
rect 274403 158611 274469 158612
rect 276059 158676 276125 158677
rect 276059 158612 276060 158676
rect 276124 158612 276125 158676
rect 276059 158611 276125 158612
rect 273667 157724 273733 157725
rect 273667 157660 273668 157724
rect 273732 157660 273733 157724
rect 273667 157659 273733 157660
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4496 272414 20898
rect 271794 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 272414 -4496
rect 271794 -4816 272414 -4732
rect 271794 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 272414 -4816
rect 271794 -7964 272414 -5052
rect 276294 133954 276914 158000
rect 278454 157725 278514 159838
rect 279165 159836 279166 159900
rect 279230 159836 279231 159900
rect 279165 159835 279231 159836
rect 280936 159490 280996 160106
rect 283520 159898 283580 160106
rect 285968 159901 286028 160106
rect 285965 159900 286031 159901
rect 283520 159838 283666 159898
rect 280936 159430 281090 159490
rect 281030 158677 281090 159430
rect 283606 158677 283666 159838
rect 285965 159836 285966 159900
rect 286030 159836 286031 159900
rect 285965 159835 286031 159836
rect 288280 159490 288340 160106
rect 291000 159629 291060 160106
rect 290997 159628 291063 159629
rect 290997 159564 290998 159628
rect 291062 159564 291063 159628
rect 290997 159563 291063 159564
rect 288206 159430 288340 159490
rect 293448 159490 293508 160106
rect 295896 159490 295956 160106
rect 298480 159490 298540 160106
rect 300928 159490 300988 160106
rect 303512 159490 303572 160106
rect 293448 159430 293602 159490
rect 295896 159430 295994 159490
rect 298480 159430 298570 159490
rect 281027 158676 281093 158677
rect 281027 158612 281028 158676
rect 281092 158612 281093 158676
rect 281027 158611 281093 158612
rect 283603 158676 283669 158677
rect 283603 158612 283604 158676
rect 283668 158612 283669 158676
rect 283603 158611 283669 158612
rect 278451 157724 278517 157725
rect 278451 157660 278452 157724
rect 278516 157660 278517 157724
rect 278451 157659 278517 157660
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5456 276914 25398
rect 276294 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 276914 -5456
rect 276294 -5776 276914 -5692
rect 276294 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 276914 -5776
rect 276294 -7964 276914 -6012
rect 280794 138454 281414 158000
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6416 281414 29898
rect 280794 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 281414 -6416
rect 280794 -6736 281414 -6652
rect 280794 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 281414 -6736
rect 280794 -7964 281414 -6972
rect 285294 142954 285914 158000
rect 288206 157589 288266 159430
rect 293542 158677 293602 159430
rect 295934 158677 295994 159430
rect 298510 158677 298570 159430
rect 300902 159430 300988 159490
rect 303478 159430 303572 159490
rect 305960 159490 306020 160106
rect 308544 159490 308604 160106
rect 310992 159490 311052 160106
rect 313440 159490 313500 160106
rect 315888 159490 315948 160106
rect 305960 159430 306114 159490
rect 308544 159430 308690 159490
rect 310992 159430 311082 159490
rect 300902 158677 300962 159430
rect 303478 158677 303538 159430
rect 306054 158677 306114 159430
rect 308630 158677 308690 159430
rect 311022 158677 311082 159430
rect 313414 159430 313500 159490
rect 315806 159430 315948 159490
rect 318472 159490 318532 160106
rect 320920 159490 320980 160106
rect 323368 159490 323428 160106
rect 325952 159490 326012 160106
rect 318472 159430 318626 159490
rect 320920 159430 321018 159490
rect 313414 158677 313474 159430
rect 315806 158677 315866 159430
rect 318566 158677 318626 159430
rect 320958 158677 321018 159430
rect 323350 159430 323428 159490
rect 325926 159430 326012 159490
rect 323350 158677 323410 159430
rect 325926 158677 325986 159430
rect 357574 158813 357634 244699
rect 357571 158812 357637 158813
rect 357571 158748 357572 158812
rect 357636 158748 357637 158812
rect 357571 158747 357637 158748
rect 293539 158676 293605 158677
rect 293539 158612 293540 158676
rect 293604 158612 293605 158676
rect 293539 158611 293605 158612
rect 295931 158676 295997 158677
rect 295931 158612 295932 158676
rect 295996 158612 295997 158676
rect 295931 158611 295997 158612
rect 298507 158676 298573 158677
rect 298507 158612 298508 158676
rect 298572 158612 298573 158676
rect 298507 158611 298573 158612
rect 300899 158676 300965 158677
rect 300899 158612 300900 158676
rect 300964 158612 300965 158676
rect 300899 158611 300965 158612
rect 303475 158676 303541 158677
rect 303475 158612 303476 158676
rect 303540 158612 303541 158676
rect 303475 158611 303541 158612
rect 306051 158676 306117 158677
rect 306051 158612 306052 158676
rect 306116 158612 306117 158676
rect 306051 158611 306117 158612
rect 308627 158676 308693 158677
rect 308627 158612 308628 158676
rect 308692 158612 308693 158676
rect 308627 158611 308693 158612
rect 311019 158676 311085 158677
rect 311019 158612 311020 158676
rect 311084 158612 311085 158676
rect 311019 158611 311085 158612
rect 313411 158676 313477 158677
rect 313411 158612 313412 158676
rect 313476 158612 313477 158676
rect 313411 158611 313477 158612
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 318563 158676 318629 158677
rect 318563 158612 318564 158676
rect 318628 158612 318629 158676
rect 318563 158611 318629 158612
rect 320955 158676 321021 158677
rect 320955 158612 320956 158676
rect 321020 158612 321021 158676
rect 320955 158611 321021 158612
rect 323347 158676 323413 158677
rect 323347 158612 323348 158676
rect 323412 158612 323413 158676
rect 323347 158611 323413 158612
rect 325923 158676 325989 158677
rect 325923 158612 325924 158676
rect 325988 158612 325989 158676
rect 325923 158611 325989 158612
rect 288203 157588 288269 157589
rect 288203 157524 288204 157588
rect 288268 157524 288269 157588
rect 288203 157523 288269 157524
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7376 285914 34398
rect 285294 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 285914 -7376
rect 285294 -7696 285914 -7612
rect 285294 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 285914 -7696
rect 285294 -7964 285914 -7932
rect 289794 147454 290414 158000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -656 290414 2898
rect 289794 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 290414 -656
rect 289794 -976 290414 -892
rect 289794 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 290414 -976
rect 289794 -7964 290414 -1212
rect 294294 151954 294914 158000
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1616 294914 7398
rect 294294 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 294914 -1616
rect 294294 -1936 294914 -1852
rect 294294 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 294914 -1936
rect 294294 -7964 294914 -2172
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2576 299414 11898
rect 298794 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 299414 -2576
rect 298794 -2896 299414 -2812
rect 298794 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 299414 -2896
rect 298794 -7964 299414 -3132
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3536 303914 16398
rect 303294 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 303914 -3536
rect 303294 -3856 303914 -3772
rect 303294 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 303914 -3856
rect 303294 -7964 303914 -4092
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4496 308414 20898
rect 307794 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 308414 -4496
rect 307794 -4816 308414 -4732
rect 307794 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 308414 -4816
rect 307794 -7964 308414 -5052
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5456 312914 25398
rect 312294 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 312914 -5456
rect 312294 -5776 312914 -5692
rect 312294 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 312914 -5776
rect 312294 -7964 312914 -6012
rect 316794 138454 317414 158000
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6416 317414 29898
rect 316794 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 317414 -6416
rect 316794 -6736 317414 -6652
rect 316794 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 317414 -6736
rect 316794 -7964 317414 -6972
rect 321294 142954 321914 158000
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7376 321914 34398
rect 321294 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 321914 -7376
rect 321294 -7696 321914 -7612
rect 321294 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 321914 -7696
rect 321294 -7964 321914 -7932
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -656 326414 2898
rect 325794 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 326414 -656
rect 325794 -976 326414 -892
rect 325794 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 326414 -976
rect 325794 -7964 326414 -1212
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1616 330914 7398
rect 330294 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 330914 -1616
rect 330294 -1936 330914 -1852
rect 330294 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 330914 -1936
rect 330294 -7964 330914 -2172
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2576 335414 11898
rect 334794 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 335414 -2576
rect 334794 -2896 335414 -2812
rect 334794 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 335414 -2896
rect 334794 -7964 335414 -3132
rect 339294 124954 339914 158000
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3536 339914 16398
rect 339294 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 339914 -3536
rect 339294 -3856 339914 -3772
rect 339294 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 339914 -3856
rect 339294 -7964 339914 -4092
rect 343794 129454 344414 158000
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4496 344414 20898
rect 343794 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 344414 -4496
rect 343794 -4816 344414 -4732
rect 343794 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 344414 -4816
rect 343794 -7964 344414 -5052
rect 348294 133954 348914 158000
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5456 348914 25398
rect 348294 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 348914 -5456
rect 348294 -5776 348914 -5692
rect 348294 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 348914 -5776
rect 348294 -7964 348914 -6012
rect 352794 138454 353414 158000
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6416 353414 29898
rect 352794 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 353414 -6416
rect 352794 -6736 353414 -6652
rect 352794 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 353414 -6736
rect 352794 -7964 353414 -6972
rect 357294 142954 357914 158000
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7376 357914 34398
rect 358126 3637 358186 245515
rect 358307 245444 358373 245445
rect 358307 245380 358308 245444
rect 358372 245380 358373 245444
rect 358307 245379 358373 245380
rect 358123 3636 358189 3637
rect 358123 3572 358124 3636
rect 358188 3572 358189 3636
rect 358123 3571 358189 3572
rect 358310 3501 358370 245379
rect 358491 245308 358557 245309
rect 358491 245244 358492 245308
rect 358556 245244 358557 245308
rect 358491 245243 358557 245244
rect 358494 3773 358554 245243
rect 358491 3772 358557 3773
rect 358491 3708 358492 3772
rect 358556 3708 358557 3772
rect 358491 3707 358557 3708
rect 358862 3501 358922 264147
rect 360147 246260 360213 246261
rect 360147 246196 360148 246260
rect 360212 246196 360213 246260
rect 360147 246195 360213 246196
rect 359043 245172 359109 245173
rect 359043 245108 359044 245172
rect 359108 245108 359109 245172
rect 359043 245107 359109 245108
rect 358307 3500 358373 3501
rect 358307 3436 358308 3500
rect 358372 3436 358373 3500
rect 358307 3435 358373 3436
rect 358859 3500 358925 3501
rect 358859 3436 358860 3500
rect 358924 3436 358925 3500
rect 358859 3435 358925 3436
rect 359046 2957 359106 245107
rect 359227 245036 359293 245037
rect 359227 244972 359228 245036
rect 359292 244972 359293 245036
rect 359227 244971 359293 244972
rect 359230 3093 359290 244971
rect 359411 244900 359477 244901
rect 359411 244836 359412 244900
rect 359476 244836 359477 244900
rect 359411 244835 359477 244836
rect 359414 3365 359474 244835
rect 360150 3501 360210 246195
rect 360334 44301 360394 442171
rect 360515 244628 360581 244629
rect 360515 244564 360516 244628
rect 360580 244564 360581 244628
rect 360515 244563 360581 244564
rect 360331 44300 360397 44301
rect 360331 44236 360332 44300
rect 360396 44236 360397 44300
rect 360331 44235 360397 44236
rect 360518 4045 360578 244563
rect 360699 244492 360765 244493
rect 360699 244428 360700 244492
rect 360764 244428 360765 244492
rect 360699 244427 360765 244428
rect 360515 4044 360581 4045
rect 360515 3980 360516 4044
rect 360580 3980 360581 4044
rect 360515 3979 360581 3980
rect 360147 3500 360213 3501
rect 360147 3436 360148 3500
rect 360212 3436 360213 3500
rect 360147 3435 360213 3436
rect 359411 3364 359477 3365
rect 359411 3300 359412 3364
rect 359476 3300 359477 3364
rect 359411 3299 359477 3300
rect 360702 3229 360762 244427
rect 361622 5677 361682 442171
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 362907 265572 362973 265573
rect 362907 265508 362908 265572
rect 362972 265508 362973 265572
rect 362907 265507 362973 265508
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 362539 254692 362605 254693
rect 362539 254628 362540 254692
rect 362604 254628 362605 254692
rect 362539 254627 362605 254628
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361619 5676 361685 5677
rect 361619 5612 361620 5676
rect 361684 5612 361685 5676
rect 361619 5611 361685 5612
rect 361794 3454 362414 38898
rect 362542 3501 362602 254627
rect 362910 3501 362970 265507
rect 363462 71909 363522 443259
rect 363827 441692 363893 441693
rect 363827 441628 363828 441692
rect 363892 441628 363893 441692
rect 363827 441627 363893 441628
rect 363643 303244 363709 303245
rect 363643 303180 363644 303244
rect 363708 303180 363709 303244
rect 363643 303179 363709 303180
rect 363459 71908 363525 71909
rect 363459 71844 363460 71908
rect 363524 71844 363525 71908
rect 363459 71843 363525 71844
rect 363646 3501 363706 303179
rect 363830 191861 363890 441627
rect 366294 439954 366914 475398
rect 370794 707068 371414 711900
rect 370794 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 371414 707068
rect 370794 706748 371414 706832
rect 370794 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 371414 706748
rect 370794 696454 371414 706512
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 368979 444548 369045 444549
rect 368979 444484 368980 444548
rect 369044 444484 369045 444548
rect 368979 444483 369045 444484
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 364931 301476 364997 301477
rect 364931 301412 364932 301476
rect 364996 301412 364997 301476
rect 364931 301411 364997 301412
rect 364379 282164 364445 282165
rect 364379 282100 364380 282164
rect 364444 282100 364445 282164
rect 364379 282099 364445 282100
rect 363827 191860 363893 191861
rect 363827 191796 363828 191860
rect 363892 191796 363893 191860
rect 363827 191795 363893 191796
rect 364382 3637 364442 282099
rect 364563 248164 364629 248165
rect 364563 248100 364564 248164
rect 364628 248100 364629 248164
rect 364563 248099 364629 248100
rect 364566 159629 364626 248099
rect 364563 159628 364629 159629
rect 364563 159564 364564 159628
rect 364628 159564 364629 159628
rect 364563 159563 364629 159564
rect 364934 3909 364994 301411
rect 366294 295954 366914 331398
rect 367691 303108 367757 303109
rect 367691 303044 367692 303108
rect 367756 303044 367757 303108
rect 367691 303043 367757 303044
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 367139 283524 367205 283525
rect 367139 283460 367140 283524
rect 367204 283460 367205 283524
rect 367139 283459 367205 283460
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 365667 254556 365733 254557
rect 365667 254492 365668 254556
rect 365732 254492 365733 254556
rect 365667 254491 365733 254492
rect 364931 3908 364997 3909
rect 364931 3844 364932 3908
rect 364996 3844 364997 3908
rect 364931 3843 364997 3844
rect 365670 3637 365730 254491
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 364379 3636 364445 3637
rect 364379 3572 364380 3636
rect 364444 3572 364445 3636
rect 364379 3571 364445 3572
rect 365667 3636 365733 3637
rect 365667 3572 365668 3636
rect 365732 3572 365733 3636
rect 365667 3571 365733 3572
rect 360699 3228 360765 3229
rect 360699 3164 360700 3228
rect 360764 3164 360765 3228
rect 360699 3163 360765 3164
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 362539 3500 362605 3501
rect 362539 3436 362540 3500
rect 362604 3436 362605 3500
rect 362539 3435 362605 3436
rect 362907 3500 362973 3501
rect 362907 3436 362908 3500
rect 362972 3436 362973 3500
rect 362907 3435 362973 3436
rect 363643 3500 363709 3501
rect 363643 3436 363644 3500
rect 363708 3436 363709 3500
rect 363643 3435 363709 3436
rect 361794 3134 362414 3218
rect 359227 3092 359293 3093
rect 359227 3028 359228 3092
rect 359292 3028 359293 3092
rect 359227 3027 359293 3028
rect 359043 2956 359109 2957
rect 359043 2892 359044 2956
rect 359108 2892 359109 2956
rect 359043 2891 359109 2892
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 357294 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 357914 -7376
rect 357294 -7696 357914 -7612
rect 357294 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 357914 -7696
rect 357294 -7964 357914 -7932
rect 361794 -656 362414 2898
rect 361794 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 362414 -656
rect 361794 -976 362414 -892
rect 361794 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 362414 -976
rect 361794 -7964 362414 -1212
rect 366294 -1616 366914 7398
rect 367142 3637 367202 283459
rect 367323 250884 367389 250885
rect 367323 250820 367324 250884
rect 367388 250820 367389 250884
rect 367323 250819 367389 250820
rect 367326 4045 367386 250819
rect 367323 4044 367389 4045
rect 367323 3980 367324 4044
rect 367388 3980 367389 4044
rect 367323 3979 367389 3980
rect 367694 3773 367754 303043
rect 368427 297396 368493 297397
rect 368427 297332 368428 297396
rect 368492 297332 368493 297396
rect 368427 297331 368493 297332
rect 367691 3772 367757 3773
rect 367691 3708 367692 3772
rect 367756 3708 367757 3772
rect 367691 3707 367757 3708
rect 368430 3637 368490 297331
rect 368982 4861 369042 444483
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 369163 304196 369229 304197
rect 369163 304132 369164 304196
rect 369228 304132 369229 304196
rect 369163 304131 369229 304132
rect 368979 4860 369045 4861
rect 368979 4796 368980 4860
rect 369044 4796 369045 4860
rect 368979 4795 369045 4796
rect 367139 3636 367205 3637
rect 367139 3572 367140 3636
rect 367204 3572 367205 3636
rect 367139 3571 367205 3572
rect 368427 3636 368493 3637
rect 368427 3572 368428 3636
rect 368492 3572 368493 3636
rect 368427 3571 368493 3572
rect 369166 3365 369226 304131
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 369899 269788 369965 269789
rect 369899 269724 369900 269788
rect 369964 269724 369965 269788
rect 369899 269723 369965 269724
rect 369902 3637 369962 269723
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 369899 3636 369965 3637
rect 369899 3572 369900 3636
rect 369964 3572 369965 3636
rect 369899 3571 369965 3572
rect 369163 3364 369229 3365
rect 369163 3300 369164 3364
rect 369228 3300 369229 3364
rect 369163 3299 369229 3300
rect 366294 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 366914 -1616
rect 366294 -1936 366914 -1852
rect 366294 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 366914 -1936
rect 366294 -7964 366914 -2172
rect 370794 -2576 371414 11898
rect 370794 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 371414 -2576
rect 370794 -2896 371414 -2812
rect 370794 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 371414 -2896
rect 370794 -7964 371414 -3132
rect 375294 708028 375914 711900
rect 375294 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 375914 708028
rect 375294 707708 375914 707792
rect 375294 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 375914 707708
rect 375294 700954 375914 707472
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3536 375914 16398
rect 375294 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 375914 -3536
rect 375294 -3856 375914 -3772
rect 375294 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 375914 -3856
rect 375294 -7964 375914 -4092
rect 379794 708988 380414 711900
rect 379794 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 380414 708988
rect 379794 708668 380414 708752
rect 379794 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 380414 708668
rect 379794 669454 380414 708432
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4496 380414 20898
rect 379794 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 380414 -4496
rect 379794 -4816 380414 -4732
rect 379794 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 380414 -4816
rect 379794 -7964 380414 -5052
rect 384294 709948 384914 711900
rect 384294 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 384914 709948
rect 384294 709628 384914 709712
rect 384294 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 384914 709628
rect 384294 673954 384914 709392
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5456 384914 25398
rect 384294 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 384914 -5456
rect 384294 -5776 384914 -5692
rect 384294 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 384914 -5776
rect 384294 -7964 384914 -6012
rect 388794 710908 389414 711900
rect 388794 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 389414 710908
rect 388794 710588 389414 710672
rect 388794 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 389414 710588
rect 388794 678454 389414 710352
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6416 389414 29898
rect 388794 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 389414 -6416
rect 388794 -6736 389414 -6652
rect 388794 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 389414 -6736
rect 388794 -7964 389414 -6972
rect 393294 711868 393914 711900
rect 393294 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 393914 711868
rect 393294 711548 393914 711632
rect 393294 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 393914 711548
rect 393294 682954 393914 711312
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7376 393914 34398
rect 393294 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 393914 -7376
rect 393294 -7696 393914 -7612
rect 393294 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 393914 -7696
rect 393294 -7964 393914 -7932
rect 397794 705148 398414 711900
rect 397794 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 398414 705148
rect 397794 704828 398414 704912
rect 397794 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 398414 704828
rect 397794 687454 398414 704592
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -656 398414 2898
rect 397794 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 398414 -656
rect 397794 -976 398414 -892
rect 397794 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 398414 -976
rect 397794 -7964 398414 -1212
rect 402294 706108 402914 711900
rect 402294 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 402914 706108
rect 402294 705788 402914 705872
rect 402294 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 402914 705788
rect 402294 691954 402914 705552
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1616 402914 7398
rect 402294 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 402914 -1616
rect 402294 -1936 402914 -1852
rect 402294 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 402914 -1936
rect 402294 -7964 402914 -2172
rect 406794 707068 407414 711900
rect 406794 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 407414 707068
rect 406794 706748 407414 706832
rect 406794 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 407414 706748
rect 406794 696454 407414 706512
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2576 407414 11898
rect 406794 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 407414 -2576
rect 406794 -2896 407414 -2812
rect 406794 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 407414 -2896
rect 406794 -7964 407414 -3132
rect 411294 708028 411914 711900
rect 411294 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 411914 708028
rect 411294 707708 411914 707792
rect 411294 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 411914 707708
rect 411294 700954 411914 707472
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3536 411914 16398
rect 411294 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 411914 -3536
rect 411294 -3856 411914 -3772
rect 411294 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 411914 -3856
rect 411294 -7964 411914 -4092
rect 415794 708988 416414 711900
rect 415794 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 416414 708988
rect 415794 708668 416414 708752
rect 415794 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 416414 708668
rect 415794 669454 416414 708432
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4496 416414 20898
rect 415794 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 416414 -4496
rect 415794 -4816 416414 -4732
rect 415794 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 416414 -4816
rect 415794 -7964 416414 -5052
rect 420294 709948 420914 711900
rect 420294 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 420914 709948
rect 420294 709628 420914 709712
rect 420294 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 420914 709628
rect 420294 673954 420914 709392
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5456 420914 25398
rect 420294 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 420914 -5456
rect 420294 -5776 420914 -5692
rect 420294 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 420914 -5776
rect 420294 -7964 420914 -6012
rect 424794 710908 425414 711900
rect 424794 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 425414 710908
rect 424794 710588 425414 710672
rect 424794 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 425414 710588
rect 424794 678454 425414 710352
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6416 425414 29898
rect 424794 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 425414 -6416
rect 424794 -6736 425414 -6652
rect 424794 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 425414 -6736
rect 424794 -7964 425414 -6972
rect 429294 711868 429914 711900
rect 429294 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 429914 711868
rect 429294 711548 429914 711632
rect 429294 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 429914 711548
rect 429294 682954 429914 711312
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7376 429914 34398
rect 429294 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 429914 -7376
rect 429294 -7696 429914 -7612
rect 429294 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 429914 -7696
rect 429294 -7964 429914 -7932
rect 433794 705148 434414 711900
rect 433794 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 434414 705148
rect 433794 704828 434414 704912
rect 433794 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 434414 704828
rect 433794 687454 434414 704592
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -656 434414 2898
rect 433794 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 434414 -656
rect 433794 -976 434414 -892
rect 433794 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 434414 -976
rect 433794 -7964 434414 -1212
rect 438294 706108 438914 711900
rect 438294 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 438914 706108
rect 438294 705788 438914 705872
rect 438294 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 438914 705788
rect 438294 691954 438914 705552
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1616 438914 7398
rect 438294 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 438914 -1616
rect 438294 -1936 438914 -1852
rect 438294 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 438914 -1936
rect 438294 -7964 438914 -2172
rect 442794 707068 443414 711900
rect 442794 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 443414 707068
rect 442794 706748 443414 706832
rect 442794 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 443414 706748
rect 442794 696454 443414 706512
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2576 443414 11898
rect 442794 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 443414 -2576
rect 442794 -2896 443414 -2812
rect 442794 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 443414 -2896
rect 442794 -7964 443414 -3132
rect 447294 708028 447914 711900
rect 447294 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 447914 708028
rect 447294 707708 447914 707792
rect 447294 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 447914 707708
rect 447294 700954 447914 707472
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3536 447914 16398
rect 447294 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 447914 -3536
rect 447294 -3856 447914 -3772
rect 447294 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 447914 -3856
rect 447294 -7964 447914 -4092
rect 451794 708988 452414 711900
rect 451794 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 452414 708988
rect 451794 708668 452414 708752
rect 451794 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 452414 708668
rect 451794 669454 452414 708432
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4496 452414 20898
rect 451794 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 452414 -4496
rect 451794 -4816 452414 -4732
rect 451794 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 452414 -4816
rect 451794 -7964 452414 -5052
rect 456294 709948 456914 711900
rect 456294 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 456914 709948
rect 456294 709628 456914 709712
rect 456294 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 456914 709628
rect 456294 673954 456914 709392
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5456 456914 25398
rect 456294 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 456914 -5456
rect 456294 -5776 456914 -5692
rect 456294 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 456914 -5776
rect 456294 -7964 456914 -6012
rect 460794 710908 461414 711900
rect 460794 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 461414 710908
rect 460794 710588 461414 710672
rect 460794 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 461414 710588
rect 460794 678454 461414 710352
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6416 461414 29898
rect 460794 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 461414 -6416
rect 460794 -6736 461414 -6652
rect 460794 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 461414 -6736
rect 460794 -7964 461414 -6972
rect 465294 711868 465914 711900
rect 465294 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 465914 711868
rect 465294 711548 465914 711632
rect 465294 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 465914 711548
rect 465294 682954 465914 711312
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7376 465914 34398
rect 465294 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 465914 -7376
rect 465294 -7696 465914 -7612
rect 465294 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 465914 -7696
rect 465294 -7964 465914 -7932
rect 469794 705148 470414 711900
rect 469794 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 470414 705148
rect 469794 704828 470414 704912
rect 469794 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 470414 704828
rect 469794 687454 470414 704592
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -656 470414 2898
rect 469794 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 470414 -656
rect 469794 -976 470414 -892
rect 469794 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 470414 -976
rect 469794 -7964 470414 -1212
rect 474294 706108 474914 711900
rect 474294 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 474914 706108
rect 474294 705788 474914 705872
rect 474294 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 474914 705788
rect 474294 691954 474914 705552
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1616 474914 7398
rect 474294 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 474914 -1616
rect 474294 -1936 474914 -1852
rect 474294 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 474914 -1936
rect 474294 -7964 474914 -2172
rect 478794 707068 479414 711900
rect 478794 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 479414 707068
rect 478794 706748 479414 706832
rect 478794 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 479414 706748
rect 478794 696454 479414 706512
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2576 479414 11898
rect 478794 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 479414 -2576
rect 478794 -2896 479414 -2812
rect 478794 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 479414 -2896
rect 478794 -7964 479414 -3132
rect 483294 708028 483914 711900
rect 483294 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 483914 708028
rect 483294 707708 483914 707792
rect 483294 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 483914 707708
rect 483294 700954 483914 707472
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3536 483914 16398
rect 483294 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 483914 -3536
rect 483294 -3856 483914 -3772
rect 483294 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 483914 -3856
rect 483294 -7964 483914 -4092
rect 487794 708988 488414 711900
rect 487794 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 488414 708988
rect 487794 708668 488414 708752
rect 487794 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 488414 708668
rect 487794 669454 488414 708432
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4496 488414 20898
rect 487794 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 488414 -4496
rect 487794 -4816 488414 -4732
rect 487794 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 488414 -4816
rect 487794 -7964 488414 -5052
rect 492294 709948 492914 711900
rect 492294 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 492914 709948
rect 492294 709628 492914 709712
rect 492294 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 492914 709628
rect 492294 673954 492914 709392
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5456 492914 25398
rect 492294 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 492914 -5456
rect 492294 -5776 492914 -5692
rect 492294 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 492914 -5776
rect 492294 -7964 492914 -6012
rect 496794 710908 497414 711900
rect 496794 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 497414 710908
rect 496794 710588 497414 710672
rect 496794 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 497414 710588
rect 496794 678454 497414 710352
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6416 497414 29898
rect 496794 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 497414 -6416
rect 496794 -6736 497414 -6652
rect 496794 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 497414 -6736
rect 496794 -7964 497414 -6972
rect 501294 711868 501914 711900
rect 501294 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 501914 711868
rect 501294 711548 501914 711632
rect 501294 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 501914 711548
rect 501294 682954 501914 711312
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7376 501914 34398
rect 501294 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 501914 -7376
rect 501294 -7696 501914 -7612
rect 501294 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 501914 -7696
rect 501294 -7964 501914 -7932
rect 505794 705148 506414 711900
rect 505794 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 506414 705148
rect 505794 704828 506414 704912
rect 505794 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 506414 704828
rect 505794 687454 506414 704592
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -656 506414 2898
rect 505794 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 506414 -656
rect 505794 -976 506414 -892
rect 505794 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 506414 -976
rect 505794 -7964 506414 -1212
rect 510294 706108 510914 711900
rect 510294 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 510914 706108
rect 510294 705788 510914 705872
rect 510294 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 510914 705788
rect 510294 691954 510914 705552
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1616 510914 7398
rect 510294 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 510914 -1616
rect 510294 -1936 510914 -1852
rect 510294 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 510914 -1936
rect 510294 -7964 510914 -2172
rect 514794 707068 515414 711900
rect 514794 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 515414 707068
rect 514794 706748 515414 706832
rect 514794 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 515414 706748
rect 514794 696454 515414 706512
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2576 515414 11898
rect 514794 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 515414 -2576
rect 514794 -2896 515414 -2812
rect 514794 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 515414 -2896
rect 514794 -7964 515414 -3132
rect 519294 708028 519914 711900
rect 519294 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 519914 708028
rect 519294 707708 519914 707792
rect 519294 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 519914 707708
rect 519294 700954 519914 707472
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3536 519914 16398
rect 519294 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 519914 -3536
rect 519294 -3856 519914 -3772
rect 519294 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 519914 -3856
rect 519294 -7964 519914 -4092
rect 523794 708988 524414 711900
rect 523794 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 524414 708988
rect 523794 708668 524414 708752
rect 523794 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 524414 708668
rect 523794 669454 524414 708432
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4496 524414 20898
rect 523794 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 524414 -4496
rect 523794 -4816 524414 -4732
rect 523794 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 524414 -4816
rect 523794 -7964 524414 -5052
rect 528294 709948 528914 711900
rect 528294 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 528914 709948
rect 528294 709628 528914 709712
rect 528294 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 528914 709628
rect 528294 673954 528914 709392
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5456 528914 25398
rect 528294 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 528914 -5456
rect 528294 -5776 528914 -5692
rect 528294 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 528914 -5776
rect 528294 -7964 528914 -6012
rect 532794 710908 533414 711900
rect 532794 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 533414 710908
rect 532794 710588 533414 710672
rect 532794 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 533414 710588
rect 532794 678454 533414 710352
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6416 533414 29898
rect 532794 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 533414 -6416
rect 532794 -6736 533414 -6652
rect 532794 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 533414 -6736
rect 532794 -7964 533414 -6972
rect 537294 711868 537914 711900
rect 537294 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 537914 711868
rect 537294 711548 537914 711632
rect 537294 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 537914 711548
rect 537294 682954 537914 711312
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7376 537914 34398
rect 537294 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 537914 -7376
rect 537294 -7696 537914 -7612
rect 537294 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 537914 -7696
rect 537294 -7964 537914 -7932
rect 541794 705148 542414 711900
rect 541794 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 542414 705148
rect 541794 704828 542414 704912
rect 541794 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 542414 704828
rect 541794 687454 542414 704592
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -656 542414 2898
rect 541794 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 542414 -656
rect 541794 -976 542414 -892
rect 541794 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 542414 -976
rect 541794 -7964 542414 -1212
rect 546294 706108 546914 711900
rect 546294 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 546914 706108
rect 546294 705788 546914 705872
rect 546294 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 546914 705788
rect 546294 691954 546914 705552
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1616 546914 7398
rect 546294 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 546914 -1616
rect 546294 -1936 546914 -1852
rect 546294 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 546914 -1936
rect 546294 -7964 546914 -2172
rect 550794 707068 551414 711900
rect 550794 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 551414 707068
rect 550794 706748 551414 706832
rect 550794 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 551414 706748
rect 550794 696454 551414 706512
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2576 551414 11898
rect 550794 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 551414 -2576
rect 550794 -2896 551414 -2812
rect 550794 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 551414 -2896
rect 550794 -7964 551414 -3132
rect 555294 708028 555914 711900
rect 555294 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 555914 708028
rect 555294 707708 555914 707792
rect 555294 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 555914 707708
rect 555294 700954 555914 707472
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3536 555914 16398
rect 555294 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 555914 -3536
rect 555294 -3856 555914 -3772
rect 555294 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 555914 -3856
rect 555294 -7964 555914 -4092
rect 559794 708988 560414 711900
rect 559794 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 560414 708988
rect 559794 708668 560414 708752
rect 559794 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 560414 708668
rect 559794 669454 560414 708432
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4496 560414 20898
rect 559794 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 560414 -4496
rect 559794 -4816 560414 -4732
rect 559794 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 560414 -4816
rect 559794 -7964 560414 -5052
rect 564294 709948 564914 711900
rect 564294 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 564914 709948
rect 564294 709628 564914 709712
rect 564294 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 564914 709628
rect 564294 673954 564914 709392
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5456 564914 25398
rect 564294 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 564914 -5456
rect 564294 -5776 564914 -5692
rect 564294 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 564914 -5776
rect 564294 -7964 564914 -6012
rect 568794 710908 569414 711900
rect 568794 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 569414 710908
rect 568794 710588 569414 710672
rect 568794 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 569414 710588
rect 568794 678454 569414 710352
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6416 569414 29898
rect 568794 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 569414 -6416
rect 568794 -6736 569414 -6652
rect 568794 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 569414 -6736
rect 568794 -7964 569414 -6972
rect 573294 711868 573914 711900
rect 573294 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 573914 711868
rect 573294 711548 573914 711632
rect 573294 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 573914 711548
rect 573294 682954 573914 711312
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7376 573914 34398
rect 573294 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 573914 -7376
rect 573294 -7696 573914 -7612
rect 573294 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 573914 -7696
rect 573294 -7964 573914 -7932
rect 577794 705148 578414 711900
rect 577794 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 578414 705148
rect 577794 704828 578414 704912
rect 577794 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 578414 704828
rect 577794 687454 578414 704592
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -656 578414 2898
rect 577794 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 578414 -656
rect 577794 -976 578414 -892
rect 577794 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 578414 -976
rect 577794 -7964 578414 -1212
rect 582294 706108 582914 711900
rect 592340 711868 592960 711900
rect 592340 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect 592340 711548 592960 711632
rect 592340 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect 591380 710908 592000 710940
rect 591380 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect 591380 710588 592000 710672
rect 591380 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect 590420 709948 591040 709980
rect 590420 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect 590420 709628 591040 709712
rect 590420 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect 589460 708988 590080 709020
rect 589460 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect 589460 708668 590080 708752
rect 589460 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect 588500 708028 589120 708060
rect 588500 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect 588500 707708 589120 707792
rect 588500 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect 587540 707068 588160 707100
rect 587540 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect 587540 706748 588160 706832
rect 587540 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect 582294 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 582914 706108
rect 582294 705788 582914 705872
rect 582294 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 582914 705788
rect 582294 691954 582914 705552
rect 586580 706108 587200 706140
rect 586580 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect 586580 705788 587200 705872
rect 586580 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1616 582914 7398
rect 585620 705148 586240 705180
rect 585620 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect 585620 704828 586240 704912
rect 585620 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect 585620 687454 586240 704592
rect 585620 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 586240 687454
rect 585620 687134 586240 687218
rect 585620 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 586240 687134
rect 585620 651454 586240 686898
rect 585620 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 586240 651454
rect 585620 651134 586240 651218
rect 585620 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 586240 651134
rect 585620 615454 586240 650898
rect 585620 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 586240 615454
rect 585620 615134 586240 615218
rect 585620 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 586240 615134
rect 585620 579454 586240 614898
rect 585620 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 586240 579454
rect 585620 579134 586240 579218
rect 585620 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 586240 579134
rect 585620 543454 586240 578898
rect 585620 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 586240 543454
rect 585620 543134 586240 543218
rect 585620 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 586240 543134
rect 585620 507454 586240 542898
rect 585620 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 586240 507454
rect 585620 507134 586240 507218
rect 585620 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 586240 507134
rect 585620 471454 586240 506898
rect 585620 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 586240 471454
rect 585620 471134 586240 471218
rect 585620 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 586240 471134
rect 585620 435454 586240 470898
rect 585620 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 586240 435454
rect 585620 435134 586240 435218
rect 585620 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 586240 435134
rect 585620 399454 586240 434898
rect 585620 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 586240 399454
rect 585620 399134 586240 399218
rect 585620 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 586240 399134
rect 585620 363454 586240 398898
rect 585620 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 586240 363454
rect 585620 363134 586240 363218
rect 585620 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 586240 363134
rect 585620 327454 586240 362898
rect 585620 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 586240 327454
rect 585620 327134 586240 327218
rect 585620 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 586240 327134
rect 585620 291454 586240 326898
rect 585620 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 586240 291454
rect 585620 291134 586240 291218
rect 585620 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 586240 291134
rect 585620 255454 586240 290898
rect 585620 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 586240 255454
rect 585620 255134 586240 255218
rect 585620 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 586240 255134
rect 585620 219454 586240 254898
rect 585620 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 586240 219454
rect 585620 219134 586240 219218
rect 585620 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 586240 219134
rect 585620 183454 586240 218898
rect 585620 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 586240 183454
rect 585620 183134 586240 183218
rect 585620 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 586240 183134
rect 585620 147454 586240 182898
rect 585620 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 586240 147454
rect 585620 147134 586240 147218
rect 585620 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 586240 147134
rect 585620 111454 586240 146898
rect 585620 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 586240 111454
rect 585620 111134 586240 111218
rect 585620 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 586240 111134
rect 585620 75454 586240 110898
rect 585620 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 586240 75454
rect 585620 75134 586240 75218
rect 585620 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 586240 75134
rect 585620 39454 586240 74898
rect 585620 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 586240 39454
rect 585620 39134 586240 39218
rect 585620 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 586240 39134
rect 585620 3454 586240 38898
rect 585620 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 586240 3454
rect 585620 3134 586240 3218
rect 585620 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 586240 3134
rect 585620 -656 586240 2898
rect 585620 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect 585620 -976 586240 -892
rect 585620 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect 585620 -1244 586240 -1212
rect 586580 691954 587200 705552
rect 586580 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 587200 691954
rect 586580 691634 587200 691718
rect 586580 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 587200 691634
rect 586580 655954 587200 691398
rect 586580 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 587200 655954
rect 586580 655634 587200 655718
rect 586580 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 587200 655634
rect 586580 619954 587200 655398
rect 586580 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 587200 619954
rect 586580 619634 587200 619718
rect 586580 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 587200 619634
rect 586580 583954 587200 619398
rect 586580 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 587200 583954
rect 586580 583634 587200 583718
rect 586580 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 587200 583634
rect 586580 547954 587200 583398
rect 586580 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 587200 547954
rect 586580 547634 587200 547718
rect 586580 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 587200 547634
rect 586580 511954 587200 547398
rect 586580 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 587200 511954
rect 586580 511634 587200 511718
rect 586580 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 587200 511634
rect 586580 475954 587200 511398
rect 586580 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 587200 475954
rect 586580 475634 587200 475718
rect 586580 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 587200 475634
rect 586580 439954 587200 475398
rect 586580 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 587200 439954
rect 586580 439634 587200 439718
rect 586580 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 587200 439634
rect 586580 403954 587200 439398
rect 586580 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 587200 403954
rect 586580 403634 587200 403718
rect 586580 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 587200 403634
rect 586580 367954 587200 403398
rect 586580 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 587200 367954
rect 586580 367634 587200 367718
rect 586580 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 587200 367634
rect 586580 331954 587200 367398
rect 586580 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 587200 331954
rect 586580 331634 587200 331718
rect 586580 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 587200 331634
rect 586580 295954 587200 331398
rect 586580 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 587200 295954
rect 586580 295634 587200 295718
rect 586580 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 587200 295634
rect 586580 259954 587200 295398
rect 586580 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 587200 259954
rect 586580 259634 587200 259718
rect 586580 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 587200 259634
rect 586580 223954 587200 259398
rect 586580 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 587200 223954
rect 586580 223634 587200 223718
rect 586580 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 587200 223634
rect 586580 187954 587200 223398
rect 586580 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 587200 187954
rect 586580 187634 587200 187718
rect 586580 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 587200 187634
rect 586580 151954 587200 187398
rect 586580 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 587200 151954
rect 586580 151634 587200 151718
rect 586580 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 587200 151634
rect 586580 115954 587200 151398
rect 586580 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 587200 115954
rect 586580 115634 587200 115718
rect 586580 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 587200 115634
rect 586580 79954 587200 115398
rect 586580 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 587200 79954
rect 586580 79634 587200 79718
rect 586580 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 587200 79634
rect 586580 43954 587200 79398
rect 586580 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 587200 43954
rect 586580 43634 587200 43718
rect 586580 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 587200 43634
rect 586580 7954 587200 43398
rect 586580 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 587200 7954
rect 586580 7634 587200 7718
rect 586580 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 587200 7634
rect 582294 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 582914 -1616
rect 582294 -1936 582914 -1852
rect 582294 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 582914 -1936
rect 582294 -7964 582914 -2172
rect 586580 -1616 587200 7398
rect 586580 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect 586580 -1936 587200 -1852
rect 586580 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect 586580 -2204 587200 -2172
rect 587540 696454 588160 706512
rect 587540 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 588160 696454
rect 587540 696134 588160 696218
rect 587540 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 588160 696134
rect 587540 660454 588160 695898
rect 587540 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 588160 660454
rect 587540 660134 588160 660218
rect 587540 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 588160 660134
rect 587540 624454 588160 659898
rect 587540 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 588160 624454
rect 587540 624134 588160 624218
rect 587540 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 588160 624134
rect 587540 588454 588160 623898
rect 587540 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 588160 588454
rect 587540 588134 588160 588218
rect 587540 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 588160 588134
rect 587540 552454 588160 587898
rect 587540 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 588160 552454
rect 587540 552134 588160 552218
rect 587540 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 588160 552134
rect 587540 516454 588160 551898
rect 587540 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 588160 516454
rect 587540 516134 588160 516218
rect 587540 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 588160 516134
rect 587540 480454 588160 515898
rect 587540 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 588160 480454
rect 587540 480134 588160 480218
rect 587540 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 588160 480134
rect 587540 444454 588160 479898
rect 587540 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 588160 444454
rect 587540 444134 588160 444218
rect 587540 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 588160 444134
rect 587540 408454 588160 443898
rect 587540 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 588160 408454
rect 587540 408134 588160 408218
rect 587540 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 588160 408134
rect 587540 372454 588160 407898
rect 587540 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 588160 372454
rect 587540 372134 588160 372218
rect 587540 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 588160 372134
rect 587540 336454 588160 371898
rect 587540 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 588160 336454
rect 587540 336134 588160 336218
rect 587540 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 588160 336134
rect 587540 300454 588160 335898
rect 587540 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 588160 300454
rect 587540 300134 588160 300218
rect 587540 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 588160 300134
rect 587540 264454 588160 299898
rect 587540 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 588160 264454
rect 587540 264134 588160 264218
rect 587540 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 588160 264134
rect 587540 228454 588160 263898
rect 587540 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 588160 228454
rect 587540 228134 588160 228218
rect 587540 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 588160 228134
rect 587540 192454 588160 227898
rect 587540 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 588160 192454
rect 587540 192134 588160 192218
rect 587540 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 588160 192134
rect 587540 156454 588160 191898
rect 587540 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 588160 156454
rect 587540 156134 588160 156218
rect 587540 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 588160 156134
rect 587540 120454 588160 155898
rect 587540 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 588160 120454
rect 587540 120134 588160 120218
rect 587540 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 588160 120134
rect 587540 84454 588160 119898
rect 587540 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 588160 84454
rect 587540 84134 588160 84218
rect 587540 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 588160 84134
rect 587540 48454 588160 83898
rect 587540 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 588160 48454
rect 587540 48134 588160 48218
rect 587540 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 588160 48134
rect 587540 12454 588160 47898
rect 587540 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 588160 12454
rect 587540 12134 588160 12218
rect 587540 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 588160 12134
rect 587540 -2576 588160 11898
rect 587540 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect 587540 -2896 588160 -2812
rect 587540 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect 587540 -3164 588160 -3132
rect 588500 700954 589120 707472
rect 588500 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 589120 700954
rect 588500 700634 589120 700718
rect 588500 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 589120 700634
rect 588500 664954 589120 700398
rect 588500 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 589120 664954
rect 588500 664634 589120 664718
rect 588500 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 589120 664634
rect 588500 628954 589120 664398
rect 588500 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 589120 628954
rect 588500 628634 589120 628718
rect 588500 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 589120 628634
rect 588500 592954 589120 628398
rect 588500 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 589120 592954
rect 588500 592634 589120 592718
rect 588500 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 589120 592634
rect 588500 556954 589120 592398
rect 588500 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 589120 556954
rect 588500 556634 589120 556718
rect 588500 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 589120 556634
rect 588500 520954 589120 556398
rect 588500 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 589120 520954
rect 588500 520634 589120 520718
rect 588500 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 589120 520634
rect 588500 484954 589120 520398
rect 588500 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 589120 484954
rect 588500 484634 589120 484718
rect 588500 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 589120 484634
rect 588500 448954 589120 484398
rect 588500 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 589120 448954
rect 588500 448634 589120 448718
rect 588500 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 589120 448634
rect 588500 412954 589120 448398
rect 588500 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 589120 412954
rect 588500 412634 589120 412718
rect 588500 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 589120 412634
rect 588500 376954 589120 412398
rect 588500 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 589120 376954
rect 588500 376634 589120 376718
rect 588500 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 589120 376634
rect 588500 340954 589120 376398
rect 588500 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 589120 340954
rect 588500 340634 589120 340718
rect 588500 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 589120 340634
rect 588500 304954 589120 340398
rect 588500 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 589120 304954
rect 588500 304634 589120 304718
rect 588500 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 589120 304634
rect 588500 268954 589120 304398
rect 588500 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 589120 268954
rect 588500 268634 589120 268718
rect 588500 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 589120 268634
rect 588500 232954 589120 268398
rect 588500 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 589120 232954
rect 588500 232634 589120 232718
rect 588500 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 589120 232634
rect 588500 196954 589120 232398
rect 588500 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 589120 196954
rect 588500 196634 589120 196718
rect 588500 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 589120 196634
rect 588500 160954 589120 196398
rect 588500 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 589120 160954
rect 588500 160634 589120 160718
rect 588500 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 589120 160634
rect 588500 124954 589120 160398
rect 588500 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 589120 124954
rect 588500 124634 589120 124718
rect 588500 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 589120 124634
rect 588500 88954 589120 124398
rect 588500 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 589120 88954
rect 588500 88634 589120 88718
rect 588500 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 589120 88634
rect 588500 52954 589120 88398
rect 588500 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 589120 52954
rect 588500 52634 589120 52718
rect 588500 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 589120 52634
rect 588500 16954 589120 52398
rect 588500 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 589120 16954
rect 588500 16634 589120 16718
rect 588500 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 589120 16634
rect 588500 -3536 589120 16398
rect 588500 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect 588500 -3856 589120 -3772
rect 588500 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect 588500 -4124 589120 -4092
rect 589460 669454 590080 708432
rect 589460 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 590080 669454
rect 589460 669134 590080 669218
rect 589460 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 590080 669134
rect 589460 633454 590080 668898
rect 589460 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 590080 633454
rect 589460 633134 590080 633218
rect 589460 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 590080 633134
rect 589460 597454 590080 632898
rect 589460 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 590080 597454
rect 589460 597134 590080 597218
rect 589460 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 590080 597134
rect 589460 561454 590080 596898
rect 589460 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 590080 561454
rect 589460 561134 590080 561218
rect 589460 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 590080 561134
rect 589460 525454 590080 560898
rect 589460 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 590080 525454
rect 589460 525134 590080 525218
rect 589460 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 590080 525134
rect 589460 489454 590080 524898
rect 589460 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 590080 489454
rect 589460 489134 590080 489218
rect 589460 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 590080 489134
rect 589460 453454 590080 488898
rect 589460 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 590080 453454
rect 589460 453134 590080 453218
rect 589460 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 590080 453134
rect 589460 417454 590080 452898
rect 589460 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 590080 417454
rect 589460 417134 590080 417218
rect 589460 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 590080 417134
rect 589460 381454 590080 416898
rect 589460 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 590080 381454
rect 589460 381134 590080 381218
rect 589460 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 590080 381134
rect 589460 345454 590080 380898
rect 589460 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 590080 345454
rect 589460 345134 590080 345218
rect 589460 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 590080 345134
rect 589460 309454 590080 344898
rect 589460 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 590080 309454
rect 589460 309134 590080 309218
rect 589460 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 590080 309134
rect 589460 273454 590080 308898
rect 589460 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 590080 273454
rect 589460 273134 590080 273218
rect 589460 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 590080 273134
rect 589460 237454 590080 272898
rect 589460 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 590080 237454
rect 589460 237134 590080 237218
rect 589460 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 590080 237134
rect 589460 201454 590080 236898
rect 589460 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 590080 201454
rect 589460 201134 590080 201218
rect 589460 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 590080 201134
rect 589460 165454 590080 200898
rect 589460 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 590080 165454
rect 589460 165134 590080 165218
rect 589460 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 590080 165134
rect 589460 129454 590080 164898
rect 589460 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 590080 129454
rect 589460 129134 590080 129218
rect 589460 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 590080 129134
rect 589460 93454 590080 128898
rect 589460 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 590080 93454
rect 589460 93134 590080 93218
rect 589460 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 590080 93134
rect 589460 57454 590080 92898
rect 589460 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 590080 57454
rect 589460 57134 590080 57218
rect 589460 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 590080 57134
rect 589460 21454 590080 56898
rect 589460 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 590080 21454
rect 589460 21134 590080 21218
rect 589460 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 590080 21134
rect 589460 -4496 590080 20898
rect 589460 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect 589460 -4816 590080 -4732
rect 589460 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect 589460 -5084 590080 -5052
rect 590420 673954 591040 709392
rect 590420 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 591040 673954
rect 590420 673634 591040 673718
rect 590420 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 591040 673634
rect 590420 637954 591040 673398
rect 590420 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 591040 637954
rect 590420 637634 591040 637718
rect 590420 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 591040 637634
rect 590420 601954 591040 637398
rect 590420 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 591040 601954
rect 590420 601634 591040 601718
rect 590420 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 591040 601634
rect 590420 565954 591040 601398
rect 590420 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 591040 565954
rect 590420 565634 591040 565718
rect 590420 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 591040 565634
rect 590420 529954 591040 565398
rect 590420 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 591040 529954
rect 590420 529634 591040 529718
rect 590420 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 591040 529634
rect 590420 493954 591040 529398
rect 590420 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 591040 493954
rect 590420 493634 591040 493718
rect 590420 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 591040 493634
rect 590420 457954 591040 493398
rect 590420 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 591040 457954
rect 590420 457634 591040 457718
rect 590420 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 591040 457634
rect 590420 421954 591040 457398
rect 590420 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 591040 421954
rect 590420 421634 591040 421718
rect 590420 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 591040 421634
rect 590420 385954 591040 421398
rect 590420 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 591040 385954
rect 590420 385634 591040 385718
rect 590420 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 591040 385634
rect 590420 349954 591040 385398
rect 590420 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 591040 349954
rect 590420 349634 591040 349718
rect 590420 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 591040 349634
rect 590420 313954 591040 349398
rect 590420 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 591040 313954
rect 590420 313634 591040 313718
rect 590420 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 591040 313634
rect 590420 277954 591040 313398
rect 590420 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 591040 277954
rect 590420 277634 591040 277718
rect 590420 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 591040 277634
rect 590420 241954 591040 277398
rect 590420 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 591040 241954
rect 590420 241634 591040 241718
rect 590420 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 591040 241634
rect 590420 205954 591040 241398
rect 590420 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 591040 205954
rect 590420 205634 591040 205718
rect 590420 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 591040 205634
rect 590420 169954 591040 205398
rect 590420 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 591040 169954
rect 590420 169634 591040 169718
rect 590420 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 591040 169634
rect 590420 133954 591040 169398
rect 590420 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 591040 133954
rect 590420 133634 591040 133718
rect 590420 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 591040 133634
rect 590420 97954 591040 133398
rect 590420 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 591040 97954
rect 590420 97634 591040 97718
rect 590420 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 591040 97634
rect 590420 61954 591040 97398
rect 590420 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 591040 61954
rect 590420 61634 591040 61718
rect 590420 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 591040 61634
rect 590420 25954 591040 61398
rect 590420 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 591040 25954
rect 590420 25634 591040 25718
rect 590420 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 591040 25634
rect 590420 -5456 591040 25398
rect 590420 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect 590420 -5776 591040 -5692
rect 590420 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect 590420 -6044 591040 -6012
rect 591380 678454 592000 710352
rect 591380 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592000 678454
rect 591380 678134 592000 678218
rect 591380 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592000 678134
rect 591380 642454 592000 677898
rect 591380 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592000 642454
rect 591380 642134 592000 642218
rect 591380 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592000 642134
rect 591380 606454 592000 641898
rect 591380 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592000 606454
rect 591380 606134 592000 606218
rect 591380 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592000 606134
rect 591380 570454 592000 605898
rect 591380 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592000 570454
rect 591380 570134 592000 570218
rect 591380 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592000 570134
rect 591380 534454 592000 569898
rect 591380 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592000 534454
rect 591380 534134 592000 534218
rect 591380 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592000 534134
rect 591380 498454 592000 533898
rect 591380 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592000 498454
rect 591380 498134 592000 498218
rect 591380 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592000 498134
rect 591380 462454 592000 497898
rect 591380 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592000 462454
rect 591380 462134 592000 462218
rect 591380 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592000 462134
rect 591380 426454 592000 461898
rect 591380 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592000 426454
rect 591380 426134 592000 426218
rect 591380 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592000 426134
rect 591380 390454 592000 425898
rect 591380 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592000 390454
rect 591380 390134 592000 390218
rect 591380 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592000 390134
rect 591380 354454 592000 389898
rect 591380 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592000 354454
rect 591380 354134 592000 354218
rect 591380 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592000 354134
rect 591380 318454 592000 353898
rect 591380 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592000 318454
rect 591380 318134 592000 318218
rect 591380 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592000 318134
rect 591380 282454 592000 317898
rect 591380 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592000 282454
rect 591380 282134 592000 282218
rect 591380 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592000 282134
rect 591380 246454 592000 281898
rect 591380 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592000 246454
rect 591380 246134 592000 246218
rect 591380 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592000 246134
rect 591380 210454 592000 245898
rect 591380 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592000 210454
rect 591380 210134 592000 210218
rect 591380 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592000 210134
rect 591380 174454 592000 209898
rect 591380 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592000 174454
rect 591380 174134 592000 174218
rect 591380 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592000 174134
rect 591380 138454 592000 173898
rect 591380 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592000 138454
rect 591380 138134 592000 138218
rect 591380 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592000 138134
rect 591380 102454 592000 137898
rect 591380 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592000 102454
rect 591380 102134 592000 102218
rect 591380 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592000 102134
rect 591380 66454 592000 101898
rect 591380 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592000 66454
rect 591380 66134 592000 66218
rect 591380 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592000 66134
rect 591380 30454 592000 65898
rect 591380 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592000 30454
rect 591380 30134 592000 30218
rect 591380 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592000 30134
rect 591380 -6416 592000 29898
rect 591380 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect 591380 -6736 592000 -6652
rect 591380 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect 591380 -7004 592000 -6972
rect 592340 682954 592960 711312
rect 592340 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect 592340 682634 592960 682718
rect 592340 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect 592340 646954 592960 682398
rect 592340 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect 592340 646634 592960 646718
rect 592340 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect 592340 610954 592960 646398
rect 592340 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect 592340 610634 592960 610718
rect 592340 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect 592340 574954 592960 610398
rect 592340 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect 592340 574634 592960 574718
rect 592340 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect 592340 538954 592960 574398
rect 592340 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect 592340 538634 592960 538718
rect 592340 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect 592340 502954 592960 538398
rect 592340 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect 592340 502634 592960 502718
rect 592340 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect 592340 466954 592960 502398
rect 592340 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect 592340 466634 592960 466718
rect 592340 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect 592340 430954 592960 466398
rect 592340 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect 592340 430634 592960 430718
rect 592340 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect 592340 394954 592960 430398
rect 592340 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect 592340 394634 592960 394718
rect 592340 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect 592340 358954 592960 394398
rect 592340 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect 592340 358634 592960 358718
rect 592340 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect 592340 322954 592960 358398
rect 592340 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect 592340 322634 592960 322718
rect 592340 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect 592340 286954 592960 322398
rect 592340 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect 592340 286634 592960 286718
rect 592340 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect 592340 250954 592960 286398
rect 592340 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect 592340 250634 592960 250718
rect 592340 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect 592340 214954 592960 250398
rect 592340 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect 592340 214634 592960 214718
rect 592340 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect 592340 178954 592960 214398
rect 592340 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect 592340 178634 592960 178718
rect 592340 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect 592340 142954 592960 178398
rect 592340 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect 592340 142634 592960 142718
rect 592340 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect 592340 106954 592960 142398
rect 592340 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect 592340 106634 592960 106718
rect 592340 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect 592340 70954 592960 106398
rect 592340 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect 592340 70634 592960 70718
rect 592340 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect 592340 34954 592960 70398
rect 592340 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect 592340 34634 592960 34718
rect 592340 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect 592340 -7376 592960 34398
rect 592340 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect 592340 -7696 592960 -7612
rect 592340 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect 592340 -7964 592960 -7932
<< via4 >>
rect -9004 711632 -8768 711868
rect -8684 711632 -8448 711868
rect -9004 711312 -8768 711548
rect -8684 711312 -8448 711548
rect -9004 682718 -8768 682954
rect -8684 682718 -8448 682954
rect -9004 682398 -8768 682634
rect -8684 682398 -8448 682634
rect -9004 646718 -8768 646954
rect -8684 646718 -8448 646954
rect -9004 646398 -8768 646634
rect -8684 646398 -8448 646634
rect -9004 610718 -8768 610954
rect -8684 610718 -8448 610954
rect -9004 610398 -8768 610634
rect -8684 610398 -8448 610634
rect -9004 574718 -8768 574954
rect -8684 574718 -8448 574954
rect -9004 574398 -8768 574634
rect -8684 574398 -8448 574634
rect -9004 538718 -8768 538954
rect -8684 538718 -8448 538954
rect -9004 538398 -8768 538634
rect -8684 538398 -8448 538634
rect -9004 502718 -8768 502954
rect -8684 502718 -8448 502954
rect -9004 502398 -8768 502634
rect -8684 502398 -8448 502634
rect -9004 466718 -8768 466954
rect -8684 466718 -8448 466954
rect -9004 466398 -8768 466634
rect -8684 466398 -8448 466634
rect -9004 430718 -8768 430954
rect -8684 430718 -8448 430954
rect -9004 430398 -8768 430634
rect -8684 430398 -8448 430634
rect -9004 394718 -8768 394954
rect -8684 394718 -8448 394954
rect -9004 394398 -8768 394634
rect -8684 394398 -8448 394634
rect -9004 358718 -8768 358954
rect -8684 358718 -8448 358954
rect -9004 358398 -8768 358634
rect -8684 358398 -8448 358634
rect -9004 322718 -8768 322954
rect -8684 322718 -8448 322954
rect -9004 322398 -8768 322634
rect -8684 322398 -8448 322634
rect -9004 286718 -8768 286954
rect -8684 286718 -8448 286954
rect -9004 286398 -8768 286634
rect -8684 286398 -8448 286634
rect -9004 250718 -8768 250954
rect -8684 250718 -8448 250954
rect -9004 250398 -8768 250634
rect -8684 250398 -8448 250634
rect -9004 214718 -8768 214954
rect -8684 214718 -8448 214954
rect -9004 214398 -8768 214634
rect -8684 214398 -8448 214634
rect -9004 178718 -8768 178954
rect -8684 178718 -8448 178954
rect -9004 178398 -8768 178634
rect -8684 178398 -8448 178634
rect -9004 142718 -8768 142954
rect -8684 142718 -8448 142954
rect -9004 142398 -8768 142634
rect -8684 142398 -8448 142634
rect -9004 106718 -8768 106954
rect -8684 106718 -8448 106954
rect -9004 106398 -8768 106634
rect -8684 106398 -8448 106634
rect -9004 70718 -8768 70954
rect -8684 70718 -8448 70954
rect -9004 70398 -8768 70634
rect -8684 70398 -8448 70634
rect -9004 34718 -8768 34954
rect -8684 34718 -8448 34954
rect -9004 34398 -8768 34634
rect -8684 34398 -8448 34634
rect -8044 710672 -7808 710908
rect -7724 710672 -7488 710908
rect -8044 710352 -7808 710588
rect -7724 710352 -7488 710588
rect -8044 678218 -7808 678454
rect -7724 678218 -7488 678454
rect -8044 677898 -7808 678134
rect -7724 677898 -7488 678134
rect -8044 642218 -7808 642454
rect -7724 642218 -7488 642454
rect -8044 641898 -7808 642134
rect -7724 641898 -7488 642134
rect -8044 606218 -7808 606454
rect -7724 606218 -7488 606454
rect -8044 605898 -7808 606134
rect -7724 605898 -7488 606134
rect -8044 570218 -7808 570454
rect -7724 570218 -7488 570454
rect -8044 569898 -7808 570134
rect -7724 569898 -7488 570134
rect -8044 534218 -7808 534454
rect -7724 534218 -7488 534454
rect -8044 533898 -7808 534134
rect -7724 533898 -7488 534134
rect -8044 498218 -7808 498454
rect -7724 498218 -7488 498454
rect -8044 497898 -7808 498134
rect -7724 497898 -7488 498134
rect -8044 462218 -7808 462454
rect -7724 462218 -7488 462454
rect -8044 461898 -7808 462134
rect -7724 461898 -7488 462134
rect -8044 426218 -7808 426454
rect -7724 426218 -7488 426454
rect -8044 425898 -7808 426134
rect -7724 425898 -7488 426134
rect -8044 390218 -7808 390454
rect -7724 390218 -7488 390454
rect -8044 389898 -7808 390134
rect -7724 389898 -7488 390134
rect -8044 354218 -7808 354454
rect -7724 354218 -7488 354454
rect -8044 353898 -7808 354134
rect -7724 353898 -7488 354134
rect -8044 318218 -7808 318454
rect -7724 318218 -7488 318454
rect -8044 317898 -7808 318134
rect -7724 317898 -7488 318134
rect -8044 282218 -7808 282454
rect -7724 282218 -7488 282454
rect -8044 281898 -7808 282134
rect -7724 281898 -7488 282134
rect -8044 246218 -7808 246454
rect -7724 246218 -7488 246454
rect -8044 245898 -7808 246134
rect -7724 245898 -7488 246134
rect -8044 210218 -7808 210454
rect -7724 210218 -7488 210454
rect -8044 209898 -7808 210134
rect -7724 209898 -7488 210134
rect -8044 174218 -7808 174454
rect -7724 174218 -7488 174454
rect -8044 173898 -7808 174134
rect -7724 173898 -7488 174134
rect -8044 138218 -7808 138454
rect -7724 138218 -7488 138454
rect -8044 137898 -7808 138134
rect -7724 137898 -7488 138134
rect -8044 102218 -7808 102454
rect -7724 102218 -7488 102454
rect -8044 101898 -7808 102134
rect -7724 101898 -7488 102134
rect -8044 66218 -7808 66454
rect -7724 66218 -7488 66454
rect -8044 65898 -7808 66134
rect -7724 65898 -7488 66134
rect -8044 30218 -7808 30454
rect -7724 30218 -7488 30454
rect -8044 29898 -7808 30134
rect -7724 29898 -7488 30134
rect -7084 709712 -6848 709948
rect -6764 709712 -6528 709948
rect -7084 709392 -6848 709628
rect -6764 709392 -6528 709628
rect -7084 673718 -6848 673954
rect -6764 673718 -6528 673954
rect -7084 673398 -6848 673634
rect -6764 673398 -6528 673634
rect -7084 637718 -6848 637954
rect -6764 637718 -6528 637954
rect -7084 637398 -6848 637634
rect -6764 637398 -6528 637634
rect -7084 601718 -6848 601954
rect -6764 601718 -6528 601954
rect -7084 601398 -6848 601634
rect -6764 601398 -6528 601634
rect -7084 565718 -6848 565954
rect -6764 565718 -6528 565954
rect -7084 565398 -6848 565634
rect -6764 565398 -6528 565634
rect -7084 529718 -6848 529954
rect -6764 529718 -6528 529954
rect -7084 529398 -6848 529634
rect -6764 529398 -6528 529634
rect -7084 493718 -6848 493954
rect -6764 493718 -6528 493954
rect -7084 493398 -6848 493634
rect -6764 493398 -6528 493634
rect -7084 457718 -6848 457954
rect -6764 457718 -6528 457954
rect -7084 457398 -6848 457634
rect -6764 457398 -6528 457634
rect -7084 421718 -6848 421954
rect -6764 421718 -6528 421954
rect -7084 421398 -6848 421634
rect -6764 421398 -6528 421634
rect -7084 385718 -6848 385954
rect -6764 385718 -6528 385954
rect -7084 385398 -6848 385634
rect -6764 385398 -6528 385634
rect -7084 349718 -6848 349954
rect -6764 349718 -6528 349954
rect -7084 349398 -6848 349634
rect -6764 349398 -6528 349634
rect -7084 313718 -6848 313954
rect -6764 313718 -6528 313954
rect -7084 313398 -6848 313634
rect -6764 313398 -6528 313634
rect -7084 277718 -6848 277954
rect -6764 277718 -6528 277954
rect -7084 277398 -6848 277634
rect -6764 277398 -6528 277634
rect -7084 241718 -6848 241954
rect -6764 241718 -6528 241954
rect -7084 241398 -6848 241634
rect -6764 241398 -6528 241634
rect -7084 205718 -6848 205954
rect -6764 205718 -6528 205954
rect -7084 205398 -6848 205634
rect -6764 205398 -6528 205634
rect -7084 169718 -6848 169954
rect -6764 169718 -6528 169954
rect -7084 169398 -6848 169634
rect -6764 169398 -6528 169634
rect -7084 133718 -6848 133954
rect -6764 133718 -6528 133954
rect -7084 133398 -6848 133634
rect -6764 133398 -6528 133634
rect -7084 97718 -6848 97954
rect -6764 97718 -6528 97954
rect -7084 97398 -6848 97634
rect -6764 97398 -6528 97634
rect -7084 61718 -6848 61954
rect -6764 61718 -6528 61954
rect -7084 61398 -6848 61634
rect -6764 61398 -6528 61634
rect -7084 25718 -6848 25954
rect -6764 25718 -6528 25954
rect -7084 25398 -6848 25634
rect -6764 25398 -6528 25634
rect -6124 708752 -5888 708988
rect -5804 708752 -5568 708988
rect -6124 708432 -5888 708668
rect -5804 708432 -5568 708668
rect -6124 669218 -5888 669454
rect -5804 669218 -5568 669454
rect -6124 668898 -5888 669134
rect -5804 668898 -5568 669134
rect -6124 633218 -5888 633454
rect -5804 633218 -5568 633454
rect -6124 632898 -5888 633134
rect -5804 632898 -5568 633134
rect -6124 597218 -5888 597454
rect -5804 597218 -5568 597454
rect -6124 596898 -5888 597134
rect -5804 596898 -5568 597134
rect -6124 561218 -5888 561454
rect -5804 561218 -5568 561454
rect -6124 560898 -5888 561134
rect -5804 560898 -5568 561134
rect -6124 525218 -5888 525454
rect -5804 525218 -5568 525454
rect -6124 524898 -5888 525134
rect -5804 524898 -5568 525134
rect -6124 489218 -5888 489454
rect -5804 489218 -5568 489454
rect -6124 488898 -5888 489134
rect -5804 488898 -5568 489134
rect -6124 453218 -5888 453454
rect -5804 453218 -5568 453454
rect -6124 452898 -5888 453134
rect -5804 452898 -5568 453134
rect -6124 417218 -5888 417454
rect -5804 417218 -5568 417454
rect -6124 416898 -5888 417134
rect -5804 416898 -5568 417134
rect -6124 381218 -5888 381454
rect -5804 381218 -5568 381454
rect -6124 380898 -5888 381134
rect -5804 380898 -5568 381134
rect -6124 345218 -5888 345454
rect -5804 345218 -5568 345454
rect -6124 344898 -5888 345134
rect -5804 344898 -5568 345134
rect -6124 309218 -5888 309454
rect -5804 309218 -5568 309454
rect -6124 308898 -5888 309134
rect -5804 308898 -5568 309134
rect -6124 273218 -5888 273454
rect -5804 273218 -5568 273454
rect -6124 272898 -5888 273134
rect -5804 272898 -5568 273134
rect -6124 237218 -5888 237454
rect -5804 237218 -5568 237454
rect -6124 236898 -5888 237134
rect -5804 236898 -5568 237134
rect -6124 201218 -5888 201454
rect -5804 201218 -5568 201454
rect -6124 200898 -5888 201134
rect -5804 200898 -5568 201134
rect -6124 165218 -5888 165454
rect -5804 165218 -5568 165454
rect -6124 164898 -5888 165134
rect -5804 164898 -5568 165134
rect -6124 129218 -5888 129454
rect -5804 129218 -5568 129454
rect -6124 128898 -5888 129134
rect -5804 128898 -5568 129134
rect -6124 93218 -5888 93454
rect -5804 93218 -5568 93454
rect -6124 92898 -5888 93134
rect -5804 92898 -5568 93134
rect -6124 57218 -5888 57454
rect -5804 57218 -5568 57454
rect -6124 56898 -5888 57134
rect -5804 56898 -5568 57134
rect -6124 21218 -5888 21454
rect -5804 21218 -5568 21454
rect -6124 20898 -5888 21134
rect -5804 20898 -5568 21134
rect -5164 707792 -4928 708028
rect -4844 707792 -4608 708028
rect -5164 707472 -4928 707708
rect -4844 707472 -4608 707708
rect -5164 700718 -4928 700954
rect -4844 700718 -4608 700954
rect -5164 700398 -4928 700634
rect -4844 700398 -4608 700634
rect -5164 664718 -4928 664954
rect -4844 664718 -4608 664954
rect -5164 664398 -4928 664634
rect -4844 664398 -4608 664634
rect -5164 628718 -4928 628954
rect -4844 628718 -4608 628954
rect -5164 628398 -4928 628634
rect -4844 628398 -4608 628634
rect -5164 592718 -4928 592954
rect -4844 592718 -4608 592954
rect -5164 592398 -4928 592634
rect -4844 592398 -4608 592634
rect -5164 556718 -4928 556954
rect -4844 556718 -4608 556954
rect -5164 556398 -4928 556634
rect -4844 556398 -4608 556634
rect -5164 520718 -4928 520954
rect -4844 520718 -4608 520954
rect -5164 520398 -4928 520634
rect -4844 520398 -4608 520634
rect -5164 484718 -4928 484954
rect -4844 484718 -4608 484954
rect -5164 484398 -4928 484634
rect -4844 484398 -4608 484634
rect -5164 448718 -4928 448954
rect -4844 448718 -4608 448954
rect -5164 448398 -4928 448634
rect -4844 448398 -4608 448634
rect -5164 412718 -4928 412954
rect -4844 412718 -4608 412954
rect -5164 412398 -4928 412634
rect -4844 412398 -4608 412634
rect -5164 376718 -4928 376954
rect -4844 376718 -4608 376954
rect -5164 376398 -4928 376634
rect -4844 376398 -4608 376634
rect -5164 340718 -4928 340954
rect -4844 340718 -4608 340954
rect -5164 340398 -4928 340634
rect -4844 340398 -4608 340634
rect -5164 304718 -4928 304954
rect -4844 304718 -4608 304954
rect -5164 304398 -4928 304634
rect -4844 304398 -4608 304634
rect -5164 268718 -4928 268954
rect -4844 268718 -4608 268954
rect -5164 268398 -4928 268634
rect -4844 268398 -4608 268634
rect -5164 232718 -4928 232954
rect -4844 232718 -4608 232954
rect -5164 232398 -4928 232634
rect -4844 232398 -4608 232634
rect -5164 196718 -4928 196954
rect -4844 196718 -4608 196954
rect -5164 196398 -4928 196634
rect -4844 196398 -4608 196634
rect -5164 160718 -4928 160954
rect -4844 160718 -4608 160954
rect -5164 160398 -4928 160634
rect -4844 160398 -4608 160634
rect -5164 124718 -4928 124954
rect -4844 124718 -4608 124954
rect -5164 124398 -4928 124634
rect -4844 124398 -4608 124634
rect -5164 88718 -4928 88954
rect -4844 88718 -4608 88954
rect -5164 88398 -4928 88634
rect -4844 88398 -4608 88634
rect -5164 52718 -4928 52954
rect -4844 52718 -4608 52954
rect -5164 52398 -4928 52634
rect -4844 52398 -4608 52634
rect -5164 16718 -4928 16954
rect -4844 16718 -4608 16954
rect -5164 16398 -4928 16634
rect -4844 16398 -4608 16634
rect -4204 706832 -3968 707068
rect -3884 706832 -3648 707068
rect -4204 706512 -3968 706748
rect -3884 706512 -3648 706748
rect -4204 696218 -3968 696454
rect -3884 696218 -3648 696454
rect -4204 695898 -3968 696134
rect -3884 695898 -3648 696134
rect -4204 660218 -3968 660454
rect -3884 660218 -3648 660454
rect -4204 659898 -3968 660134
rect -3884 659898 -3648 660134
rect -4204 624218 -3968 624454
rect -3884 624218 -3648 624454
rect -4204 623898 -3968 624134
rect -3884 623898 -3648 624134
rect -4204 588218 -3968 588454
rect -3884 588218 -3648 588454
rect -4204 587898 -3968 588134
rect -3884 587898 -3648 588134
rect -4204 552218 -3968 552454
rect -3884 552218 -3648 552454
rect -4204 551898 -3968 552134
rect -3884 551898 -3648 552134
rect -4204 516218 -3968 516454
rect -3884 516218 -3648 516454
rect -4204 515898 -3968 516134
rect -3884 515898 -3648 516134
rect -4204 480218 -3968 480454
rect -3884 480218 -3648 480454
rect -4204 479898 -3968 480134
rect -3884 479898 -3648 480134
rect -4204 444218 -3968 444454
rect -3884 444218 -3648 444454
rect -4204 443898 -3968 444134
rect -3884 443898 -3648 444134
rect -4204 408218 -3968 408454
rect -3884 408218 -3648 408454
rect -4204 407898 -3968 408134
rect -3884 407898 -3648 408134
rect -4204 372218 -3968 372454
rect -3884 372218 -3648 372454
rect -4204 371898 -3968 372134
rect -3884 371898 -3648 372134
rect -4204 336218 -3968 336454
rect -3884 336218 -3648 336454
rect -4204 335898 -3968 336134
rect -3884 335898 -3648 336134
rect -4204 300218 -3968 300454
rect -3884 300218 -3648 300454
rect -4204 299898 -3968 300134
rect -3884 299898 -3648 300134
rect -4204 264218 -3968 264454
rect -3884 264218 -3648 264454
rect -4204 263898 -3968 264134
rect -3884 263898 -3648 264134
rect -4204 228218 -3968 228454
rect -3884 228218 -3648 228454
rect -4204 227898 -3968 228134
rect -3884 227898 -3648 228134
rect -4204 192218 -3968 192454
rect -3884 192218 -3648 192454
rect -4204 191898 -3968 192134
rect -3884 191898 -3648 192134
rect -4204 156218 -3968 156454
rect -3884 156218 -3648 156454
rect -4204 155898 -3968 156134
rect -3884 155898 -3648 156134
rect -4204 120218 -3968 120454
rect -3884 120218 -3648 120454
rect -4204 119898 -3968 120134
rect -3884 119898 -3648 120134
rect -4204 84218 -3968 84454
rect -3884 84218 -3648 84454
rect -4204 83898 -3968 84134
rect -3884 83898 -3648 84134
rect -4204 48218 -3968 48454
rect -3884 48218 -3648 48454
rect -4204 47898 -3968 48134
rect -3884 47898 -3648 48134
rect -4204 12218 -3968 12454
rect -3884 12218 -3648 12454
rect -4204 11898 -3968 12134
rect -3884 11898 -3648 12134
rect -3244 705872 -3008 706108
rect -2924 705872 -2688 706108
rect -3244 705552 -3008 705788
rect -2924 705552 -2688 705788
rect -3244 691718 -3008 691954
rect -2924 691718 -2688 691954
rect -3244 691398 -3008 691634
rect -2924 691398 -2688 691634
rect -3244 655718 -3008 655954
rect -2924 655718 -2688 655954
rect -3244 655398 -3008 655634
rect -2924 655398 -2688 655634
rect -3244 619718 -3008 619954
rect -2924 619718 -2688 619954
rect -3244 619398 -3008 619634
rect -2924 619398 -2688 619634
rect -3244 583718 -3008 583954
rect -2924 583718 -2688 583954
rect -3244 583398 -3008 583634
rect -2924 583398 -2688 583634
rect -3244 547718 -3008 547954
rect -2924 547718 -2688 547954
rect -3244 547398 -3008 547634
rect -2924 547398 -2688 547634
rect -3244 511718 -3008 511954
rect -2924 511718 -2688 511954
rect -3244 511398 -3008 511634
rect -2924 511398 -2688 511634
rect -3244 475718 -3008 475954
rect -2924 475718 -2688 475954
rect -3244 475398 -3008 475634
rect -2924 475398 -2688 475634
rect -3244 439718 -3008 439954
rect -2924 439718 -2688 439954
rect -3244 439398 -3008 439634
rect -2924 439398 -2688 439634
rect -3244 403718 -3008 403954
rect -2924 403718 -2688 403954
rect -3244 403398 -3008 403634
rect -2924 403398 -2688 403634
rect -3244 367718 -3008 367954
rect -2924 367718 -2688 367954
rect -3244 367398 -3008 367634
rect -2924 367398 -2688 367634
rect -3244 331718 -3008 331954
rect -2924 331718 -2688 331954
rect -3244 331398 -3008 331634
rect -2924 331398 -2688 331634
rect -3244 295718 -3008 295954
rect -2924 295718 -2688 295954
rect -3244 295398 -3008 295634
rect -2924 295398 -2688 295634
rect -3244 259718 -3008 259954
rect -2924 259718 -2688 259954
rect -3244 259398 -3008 259634
rect -2924 259398 -2688 259634
rect -3244 223718 -3008 223954
rect -2924 223718 -2688 223954
rect -3244 223398 -3008 223634
rect -2924 223398 -2688 223634
rect -3244 187718 -3008 187954
rect -2924 187718 -2688 187954
rect -3244 187398 -3008 187634
rect -2924 187398 -2688 187634
rect -3244 151718 -3008 151954
rect -2924 151718 -2688 151954
rect -3244 151398 -3008 151634
rect -2924 151398 -2688 151634
rect -3244 115718 -3008 115954
rect -2924 115718 -2688 115954
rect -3244 115398 -3008 115634
rect -2924 115398 -2688 115634
rect -3244 79718 -3008 79954
rect -2924 79718 -2688 79954
rect -3244 79398 -3008 79634
rect -2924 79398 -2688 79634
rect -3244 43718 -3008 43954
rect -2924 43718 -2688 43954
rect -3244 43398 -3008 43634
rect -2924 43398 -2688 43634
rect -3244 7718 -3008 7954
rect -2924 7718 -2688 7954
rect -3244 7398 -3008 7634
rect -2924 7398 -2688 7634
rect -2284 704912 -2048 705148
rect -1964 704912 -1728 705148
rect -2284 704592 -2048 704828
rect -1964 704592 -1728 704828
rect -2284 687218 -2048 687454
rect -1964 687218 -1728 687454
rect -2284 686898 -2048 687134
rect -1964 686898 -1728 687134
rect -2284 651218 -2048 651454
rect -1964 651218 -1728 651454
rect -2284 650898 -2048 651134
rect -1964 650898 -1728 651134
rect -2284 615218 -2048 615454
rect -1964 615218 -1728 615454
rect -2284 614898 -2048 615134
rect -1964 614898 -1728 615134
rect -2284 579218 -2048 579454
rect -1964 579218 -1728 579454
rect -2284 578898 -2048 579134
rect -1964 578898 -1728 579134
rect -2284 543218 -2048 543454
rect -1964 543218 -1728 543454
rect -2284 542898 -2048 543134
rect -1964 542898 -1728 543134
rect -2284 507218 -2048 507454
rect -1964 507218 -1728 507454
rect -2284 506898 -2048 507134
rect -1964 506898 -1728 507134
rect -2284 471218 -2048 471454
rect -1964 471218 -1728 471454
rect -2284 470898 -2048 471134
rect -1964 470898 -1728 471134
rect -2284 435218 -2048 435454
rect -1964 435218 -1728 435454
rect -2284 434898 -2048 435134
rect -1964 434898 -1728 435134
rect -2284 399218 -2048 399454
rect -1964 399218 -1728 399454
rect -2284 398898 -2048 399134
rect -1964 398898 -1728 399134
rect -2284 363218 -2048 363454
rect -1964 363218 -1728 363454
rect -2284 362898 -2048 363134
rect -1964 362898 -1728 363134
rect -2284 327218 -2048 327454
rect -1964 327218 -1728 327454
rect -2284 326898 -2048 327134
rect -1964 326898 -1728 327134
rect -2284 291218 -2048 291454
rect -1964 291218 -1728 291454
rect -2284 290898 -2048 291134
rect -1964 290898 -1728 291134
rect -2284 255218 -2048 255454
rect -1964 255218 -1728 255454
rect -2284 254898 -2048 255134
rect -1964 254898 -1728 255134
rect -2284 219218 -2048 219454
rect -1964 219218 -1728 219454
rect -2284 218898 -2048 219134
rect -1964 218898 -1728 219134
rect -2284 183218 -2048 183454
rect -1964 183218 -1728 183454
rect -2284 182898 -2048 183134
rect -1964 182898 -1728 183134
rect -2284 147218 -2048 147454
rect -1964 147218 -1728 147454
rect -2284 146898 -2048 147134
rect -1964 146898 -1728 147134
rect -2284 111218 -2048 111454
rect -1964 111218 -1728 111454
rect -2284 110898 -2048 111134
rect -1964 110898 -1728 111134
rect -2284 75218 -2048 75454
rect -1964 75218 -1728 75454
rect -2284 74898 -2048 75134
rect -1964 74898 -1728 75134
rect -2284 39218 -2048 39454
rect -1964 39218 -1728 39454
rect -2284 38898 -2048 39134
rect -1964 38898 -1728 39134
rect -2284 3218 -2048 3454
rect -1964 3218 -1728 3454
rect -2284 2898 -2048 3134
rect -1964 2898 -1728 3134
rect -2284 -892 -2048 -656
rect -1964 -892 -1728 -656
rect -2284 -1212 -2048 -976
rect -1964 -1212 -1728 -976
rect 1826 704912 2062 705148
rect 2146 704912 2382 705148
rect 1826 704592 2062 704828
rect 2146 704592 2382 704828
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -892 2062 -656
rect 2146 -892 2382 -656
rect 1826 -1212 2062 -976
rect 2146 -1212 2382 -976
rect -3244 -1852 -3008 -1616
rect -2924 -1852 -2688 -1616
rect -3244 -2172 -3008 -1936
rect -2924 -2172 -2688 -1936
rect -4204 -2812 -3968 -2576
rect -3884 -2812 -3648 -2576
rect -4204 -3132 -3968 -2896
rect -3884 -3132 -3648 -2896
rect -5164 -3772 -4928 -3536
rect -4844 -3772 -4608 -3536
rect -5164 -4092 -4928 -3856
rect -4844 -4092 -4608 -3856
rect -6124 -4732 -5888 -4496
rect -5804 -4732 -5568 -4496
rect -6124 -5052 -5888 -4816
rect -5804 -5052 -5568 -4816
rect -7084 -5692 -6848 -5456
rect -6764 -5692 -6528 -5456
rect -7084 -6012 -6848 -5776
rect -6764 -6012 -6528 -5776
rect -8044 -6652 -7808 -6416
rect -7724 -6652 -7488 -6416
rect -8044 -6972 -7808 -6736
rect -7724 -6972 -7488 -6736
rect -9004 -7612 -8768 -7376
rect -8684 -7612 -8448 -7376
rect -9004 -7932 -8768 -7696
rect -8684 -7932 -8448 -7696
rect 6326 705872 6562 706108
rect 6646 705872 6882 706108
rect 6326 705552 6562 705788
rect 6646 705552 6882 705788
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1852 6562 -1616
rect 6646 -1852 6882 -1616
rect 6326 -2172 6562 -1936
rect 6646 -2172 6882 -1936
rect 10826 706832 11062 707068
rect 11146 706832 11382 707068
rect 10826 706512 11062 706748
rect 11146 706512 11382 706748
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2812 11062 -2576
rect 11146 -2812 11382 -2576
rect 10826 -3132 11062 -2896
rect 11146 -3132 11382 -2896
rect 15326 707792 15562 708028
rect 15646 707792 15882 708028
rect 15326 707472 15562 707708
rect 15646 707472 15882 707708
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3772 15562 -3536
rect 15646 -3772 15882 -3536
rect 15326 -4092 15562 -3856
rect 15646 -4092 15882 -3856
rect 19826 708752 20062 708988
rect 20146 708752 20382 708988
rect 19826 708432 20062 708668
rect 20146 708432 20382 708668
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4732 20062 -4496
rect 20146 -4732 20382 -4496
rect 19826 -5052 20062 -4816
rect 20146 -5052 20382 -4816
rect 24326 709712 24562 709948
rect 24646 709712 24882 709948
rect 24326 709392 24562 709628
rect 24646 709392 24882 709628
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5692 24562 -5456
rect 24646 -5692 24882 -5456
rect 24326 -6012 24562 -5776
rect 24646 -6012 24882 -5776
rect 28826 710672 29062 710908
rect 29146 710672 29382 710908
rect 28826 710352 29062 710588
rect 29146 710352 29382 710588
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6652 29062 -6416
rect 29146 -6652 29382 -6416
rect 28826 -6972 29062 -6736
rect 29146 -6972 29382 -6736
rect 33326 711632 33562 711868
rect 33646 711632 33882 711868
rect 33326 711312 33562 711548
rect 33646 711312 33882 711548
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7612 33562 -7376
rect 33646 -7612 33882 -7376
rect 33326 -7932 33562 -7696
rect 33646 -7932 33882 -7696
rect 37826 704912 38062 705148
rect 38146 704912 38382 705148
rect 37826 704592 38062 704828
rect 38146 704592 38382 704828
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -892 38062 -656
rect 38146 -892 38382 -656
rect 37826 -1212 38062 -976
rect 38146 -1212 38382 -976
rect 42326 705872 42562 706108
rect 42646 705872 42882 706108
rect 42326 705552 42562 705788
rect 42646 705552 42882 705788
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1852 42562 -1616
rect 42646 -1852 42882 -1616
rect 42326 -2172 42562 -1936
rect 42646 -2172 42882 -1936
rect 46826 706832 47062 707068
rect 47146 706832 47382 707068
rect 46826 706512 47062 706748
rect 47146 706512 47382 706748
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2812 47062 -2576
rect 47146 -2812 47382 -2576
rect 46826 -3132 47062 -2896
rect 47146 -3132 47382 -2896
rect 51326 707792 51562 708028
rect 51646 707792 51882 708028
rect 51326 707472 51562 707708
rect 51646 707472 51882 707708
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3772 51562 -3536
rect 51646 -3772 51882 -3536
rect 51326 -4092 51562 -3856
rect 51646 -4092 51882 -3856
rect 55826 708752 56062 708988
rect 56146 708752 56382 708988
rect 55826 708432 56062 708668
rect 56146 708432 56382 708668
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4732 56062 -4496
rect 56146 -4732 56382 -4496
rect 55826 -5052 56062 -4816
rect 56146 -5052 56382 -4816
rect 60326 709712 60562 709948
rect 60646 709712 60882 709948
rect 60326 709392 60562 709628
rect 60646 709392 60882 709628
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5692 60562 -5456
rect 60646 -5692 60882 -5456
rect 60326 -6012 60562 -5776
rect 60646 -6012 60882 -5776
rect 64826 710672 65062 710908
rect 65146 710672 65382 710908
rect 64826 710352 65062 710588
rect 65146 710352 65382 710588
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6652 65062 -6416
rect 65146 -6652 65382 -6416
rect 64826 -6972 65062 -6736
rect 65146 -6972 65382 -6736
rect 69326 711632 69562 711868
rect 69646 711632 69882 711868
rect 69326 711312 69562 711548
rect 69646 711312 69882 711548
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7612 69562 -7376
rect 69646 -7612 69882 -7376
rect 69326 -7932 69562 -7696
rect 69646 -7932 69882 -7696
rect 73826 704912 74062 705148
rect 74146 704912 74382 705148
rect 73826 704592 74062 704828
rect 74146 704592 74382 704828
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -892 74062 -656
rect 74146 -892 74382 -656
rect 73826 -1212 74062 -976
rect 74146 -1212 74382 -976
rect 78326 705872 78562 706108
rect 78646 705872 78882 706108
rect 78326 705552 78562 705788
rect 78646 705552 78882 705788
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1852 78562 -1616
rect 78646 -1852 78882 -1616
rect 78326 -2172 78562 -1936
rect 78646 -2172 78882 -1936
rect 82826 706832 83062 707068
rect 83146 706832 83382 707068
rect 82826 706512 83062 706748
rect 83146 706512 83382 706748
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2812 83062 -2576
rect 83146 -2812 83382 -2576
rect 82826 -3132 83062 -2896
rect 83146 -3132 83382 -2896
rect 87326 707792 87562 708028
rect 87646 707792 87882 708028
rect 87326 707472 87562 707708
rect 87646 707472 87882 707708
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3772 87562 -3536
rect 87646 -3772 87882 -3536
rect 87326 -4092 87562 -3856
rect 87646 -4092 87882 -3856
rect 91826 708752 92062 708988
rect 92146 708752 92382 708988
rect 91826 708432 92062 708668
rect 92146 708432 92382 708668
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4732 92062 -4496
rect 92146 -4732 92382 -4496
rect 91826 -5052 92062 -4816
rect 92146 -5052 92382 -4816
rect 96326 709712 96562 709948
rect 96646 709712 96882 709948
rect 96326 709392 96562 709628
rect 96646 709392 96882 709628
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5692 96562 -5456
rect 96646 -5692 96882 -5456
rect 96326 -6012 96562 -5776
rect 96646 -6012 96882 -5776
rect 100826 710672 101062 710908
rect 101146 710672 101382 710908
rect 100826 710352 101062 710588
rect 101146 710352 101382 710588
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6652 101062 -6416
rect 101146 -6652 101382 -6416
rect 100826 -6972 101062 -6736
rect 101146 -6972 101382 -6736
rect 105326 711632 105562 711868
rect 105646 711632 105882 711868
rect 105326 711312 105562 711548
rect 105646 711312 105882 711548
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7612 105562 -7376
rect 105646 -7612 105882 -7376
rect 105326 -7932 105562 -7696
rect 105646 -7932 105882 -7696
rect 109826 704912 110062 705148
rect 110146 704912 110382 705148
rect 109826 704592 110062 704828
rect 110146 704592 110382 704828
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -892 110062 -656
rect 110146 -892 110382 -656
rect 109826 -1212 110062 -976
rect 110146 -1212 110382 -976
rect 114326 705872 114562 706108
rect 114646 705872 114882 706108
rect 114326 705552 114562 705788
rect 114646 705552 114882 705788
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1852 114562 -1616
rect 114646 -1852 114882 -1616
rect 114326 -2172 114562 -1936
rect 114646 -2172 114882 -1936
rect 118826 706832 119062 707068
rect 119146 706832 119382 707068
rect 118826 706512 119062 706748
rect 119146 706512 119382 706748
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2812 119062 -2576
rect 119146 -2812 119382 -2576
rect 118826 -3132 119062 -2896
rect 119146 -3132 119382 -2896
rect 123326 707792 123562 708028
rect 123646 707792 123882 708028
rect 123326 707472 123562 707708
rect 123646 707472 123882 707708
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3772 123562 -3536
rect 123646 -3772 123882 -3536
rect 123326 -4092 123562 -3856
rect 123646 -4092 123882 -3856
rect 127826 708752 128062 708988
rect 128146 708752 128382 708988
rect 127826 708432 128062 708668
rect 128146 708432 128382 708668
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4732 128062 -4496
rect 128146 -4732 128382 -4496
rect 127826 -5052 128062 -4816
rect 128146 -5052 128382 -4816
rect 132326 709712 132562 709948
rect 132646 709712 132882 709948
rect 132326 709392 132562 709628
rect 132646 709392 132882 709628
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5692 132562 -5456
rect 132646 -5692 132882 -5456
rect 132326 -6012 132562 -5776
rect 132646 -6012 132882 -5776
rect 136826 710672 137062 710908
rect 137146 710672 137382 710908
rect 136826 710352 137062 710588
rect 137146 710352 137382 710588
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6652 137062 -6416
rect 137146 -6652 137382 -6416
rect 136826 -6972 137062 -6736
rect 137146 -6972 137382 -6736
rect 141326 711632 141562 711868
rect 141646 711632 141882 711868
rect 141326 711312 141562 711548
rect 141646 711312 141882 711548
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7612 141562 -7376
rect 141646 -7612 141882 -7376
rect 141326 -7932 141562 -7696
rect 141646 -7932 141882 -7696
rect 145826 704912 146062 705148
rect 146146 704912 146382 705148
rect 145826 704592 146062 704828
rect 146146 704592 146382 704828
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -892 146062 -656
rect 146146 -892 146382 -656
rect 145826 -1212 146062 -976
rect 146146 -1212 146382 -976
rect 150326 705872 150562 706108
rect 150646 705872 150882 706108
rect 150326 705552 150562 705788
rect 150646 705552 150882 705788
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1852 150562 -1616
rect 150646 -1852 150882 -1616
rect 150326 -2172 150562 -1936
rect 150646 -2172 150882 -1936
rect 154826 706832 155062 707068
rect 155146 706832 155382 707068
rect 154826 706512 155062 706748
rect 155146 706512 155382 706748
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2812 155062 -2576
rect 155146 -2812 155382 -2576
rect 154826 -3132 155062 -2896
rect 155146 -3132 155382 -2896
rect 159326 707792 159562 708028
rect 159646 707792 159882 708028
rect 159326 707472 159562 707708
rect 159646 707472 159882 707708
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3772 159562 -3536
rect 159646 -3772 159882 -3536
rect 159326 -4092 159562 -3856
rect 159646 -4092 159882 -3856
rect 163826 708752 164062 708988
rect 164146 708752 164382 708988
rect 163826 708432 164062 708668
rect 164146 708432 164382 708668
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4732 164062 -4496
rect 164146 -4732 164382 -4496
rect 163826 -5052 164062 -4816
rect 164146 -5052 164382 -4816
rect 168326 709712 168562 709948
rect 168646 709712 168882 709948
rect 168326 709392 168562 709628
rect 168646 709392 168882 709628
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5692 168562 -5456
rect 168646 -5692 168882 -5456
rect 168326 -6012 168562 -5776
rect 168646 -6012 168882 -5776
rect 172826 710672 173062 710908
rect 173146 710672 173382 710908
rect 172826 710352 173062 710588
rect 173146 710352 173382 710588
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6652 173062 -6416
rect 173146 -6652 173382 -6416
rect 172826 -6972 173062 -6736
rect 173146 -6972 173382 -6736
rect 177326 711632 177562 711868
rect 177646 711632 177882 711868
rect 177326 711312 177562 711548
rect 177646 711312 177882 711548
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7612 177562 -7376
rect 177646 -7612 177882 -7376
rect 177326 -7932 177562 -7696
rect 177646 -7932 177882 -7696
rect 181826 704912 182062 705148
rect 182146 704912 182382 705148
rect 181826 704592 182062 704828
rect 182146 704592 182382 704828
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -892 182062 -656
rect 182146 -892 182382 -656
rect 181826 -1212 182062 -976
rect 182146 -1212 182382 -976
rect 186326 705872 186562 706108
rect 186646 705872 186882 706108
rect 186326 705552 186562 705788
rect 186646 705552 186882 705788
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1852 186562 -1616
rect 186646 -1852 186882 -1616
rect 186326 -2172 186562 -1936
rect 186646 -2172 186882 -1936
rect 190826 706832 191062 707068
rect 191146 706832 191382 707068
rect 190826 706512 191062 706748
rect 191146 706512 191382 706748
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2812 191062 -2576
rect 191146 -2812 191382 -2576
rect 190826 -3132 191062 -2896
rect 191146 -3132 191382 -2896
rect 195326 707792 195562 708028
rect 195646 707792 195882 708028
rect 195326 707472 195562 707708
rect 195646 707472 195882 707708
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3772 195562 -3536
rect 195646 -3772 195882 -3536
rect 195326 -4092 195562 -3856
rect 195646 -4092 195882 -3856
rect 199826 708752 200062 708988
rect 200146 708752 200382 708988
rect 199826 708432 200062 708668
rect 200146 708432 200382 708668
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4732 200062 -4496
rect 200146 -4732 200382 -4496
rect 199826 -5052 200062 -4816
rect 200146 -5052 200382 -4816
rect 204326 709712 204562 709948
rect 204646 709712 204882 709948
rect 204326 709392 204562 709628
rect 204646 709392 204882 709628
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5692 204562 -5456
rect 204646 -5692 204882 -5456
rect 204326 -6012 204562 -5776
rect 204646 -6012 204882 -5776
rect 208826 710672 209062 710908
rect 209146 710672 209382 710908
rect 208826 710352 209062 710588
rect 209146 710352 209382 710588
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 213326 711632 213562 711868
rect 213646 711632 213882 711868
rect 213326 711312 213562 711548
rect 213646 711312 213882 711548
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704912 218062 705148
rect 218146 704912 218382 705148
rect 217826 704592 218062 704828
rect 218146 704592 218382 704828
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705872 222562 706108
rect 222646 705872 222882 706108
rect 222326 705552 222562 705788
rect 222646 705552 222882 705788
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706832 227062 707068
rect 227146 706832 227382 707068
rect 226826 706512 227062 706748
rect 227146 706512 227382 706748
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707792 231562 708028
rect 231646 707792 231882 708028
rect 231326 707472 231562 707708
rect 231646 707472 231882 707708
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708752 236062 708988
rect 236146 708752 236382 708988
rect 235826 708432 236062 708668
rect 236146 708432 236382 708668
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709712 240562 709948
rect 240646 709712 240882 709948
rect 240326 709392 240562 709628
rect 240646 709392 240882 709628
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710672 245062 710908
rect 245146 710672 245382 710908
rect 244826 710352 245062 710588
rect 245146 710352 245382 710588
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711632 249562 711868
rect 249646 711632 249882 711868
rect 249326 711312 249562 711548
rect 249646 711312 249882 711548
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704912 254062 705148
rect 254146 704912 254382 705148
rect 253826 704592 254062 704828
rect 254146 704592 254382 704828
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705872 258562 706108
rect 258646 705872 258882 706108
rect 258326 705552 258562 705788
rect 258646 705552 258882 705788
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706832 263062 707068
rect 263146 706832 263382 707068
rect 262826 706512 263062 706748
rect 263146 706512 263382 706748
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707792 267562 708028
rect 267646 707792 267882 708028
rect 267326 707472 267562 707708
rect 267646 707472 267882 707708
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708752 272062 708988
rect 272146 708752 272382 708988
rect 271826 708432 272062 708668
rect 272146 708432 272382 708668
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709712 276562 709948
rect 276646 709712 276882 709948
rect 276326 709392 276562 709628
rect 276646 709392 276882 709628
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710672 281062 710908
rect 281146 710672 281382 710908
rect 280826 710352 281062 710588
rect 281146 710352 281382 710588
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711632 285562 711868
rect 285646 711632 285882 711868
rect 285326 711312 285562 711548
rect 285646 711312 285882 711548
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704912 290062 705148
rect 290146 704912 290382 705148
rect 289826 704592 290062 704828
rect 290146 704592 290382 704828
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705872 294562 706108
rect 294646 705872 294882 706108
rect 294326 705552 294562 705788
rect 294646 705552 294882 705788
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706832 299062 707068
rect 299146 706832 299382 707068
rect 298826 706512 299062 706748
rect 299146 706512 299382 706748
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707792 303562 708028
rect 303646 707792 303882 708028
rect 303326 707472 303562 707708
rect 303646 707472 303882 707708
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708752 308062 708988
rect 308146 708752 308382 708988
rect 307826 708432 308062 708668
rect 308146 708432 308382 708668
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709712 312562 709948
rect 312646 709712 312882 709948
rect 312326 709392 312562 709628
rect 312646 709392 312882 709628
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710672 317062 710908
rect 317146 710672 317382 710908
rect 316826 710352 317062 710588
rect 317146 710352 317382 710588
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711632 321562 711868
rect 321646 711632 321882 711868
rect 321326 711312 321562 711548
rect 321646 711312 321882 711548
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704912 326062 705148
rect 326146 704912 326382 705148
rect 325826 704592 326062 704828
rect 326146 704592 326382 704828
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705872 330562 706108
rect 330646 705872 330882 706108
rect 330326 705552 330562 705788
rect 330646 705552 330882 705788
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706832 335062 707068
rect 335146 706832 335382 707068
rect 334826 706512 335062 706748
rect 335146 706512 335382 706748
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707792 339562 708028
rect 339646 707792 339882 708028
rect 339326 707472 339562 707708
rect 339646 707472 339882 707708
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708752 344062 708988
rect 344146 708752 344382 708988
rect 343826 708432 344062 708668
rect 344146 708432 344382 708668
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709712 348562 709948
rect 348646 709712 348882 709948
rect 348326 709392 348562 709628
rect 348646 709392 348882 709628
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710672 353062 710908
rect 353146 710672 353382 710908
rect 352826 710352 353062 710588
rect 353146 710352 353382 710588
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711632 357562 711868
rect 357646 711632 357882 711868
rect 357326 711312 357562 711548
rect 357646 711312 357882 711548
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704912 362062 705148
rect 362146 704912 362382 705148
rect 361826 704592 362062 704828
rect 362146 704592 362382 704828
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 208826 -6652 209062 -6416
rect 209146 -6652 209382 -6416
rect 208826 -6972 209062 -6736
rect 209146 -6972 209382 -6736
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705872 366562 706108
rect 366646 705872 366882 706108
rect 366326 705552 366562 705788
rect 366646 705552 366882 705788
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 252010 439718 252246 439954
rect 252010 439398 252246 439634
rect 282730 439718 282966 439954
rect 282730 439398 282966 439634
rect 313450 439718 313686 439954
rect 313450 439398 313686 439634
rect 344170 439718 344406 439954
rect 344170 439398 344406 439634
rect 236650 435218 236886 435454
rect 236650 434898 236886 435134
rect 267370 435218 267606 435454
rect 267370 434898 267606 435134
rect 298090 435218 298326 435454
rect 298090 434898 298326 435134
rect 328810 435218 329046 435454
rect 328810 434898 329046 435134
rect 359530 435218 359766 435454
rect 359530 434898 359766 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 252010 403718 252246 403954
rect 252010 403398 252246 403634
rect 282730 403718 282966 403954
rect 282730 403398 282966 403634
rect 313450 403718 313686 403954
rect 313450 403398 313686 403634
rect 344170 403718 344406 403954
rect 344170 403398 344406 403634
rect 236650 399218 236886 399454
rect 236650 398898 236886 399134
rect 267370 399218 267606 399454
rect 267370 398898 267606 399134
rect 298090 399218 298326 399454
rect 298090 398898 298326 399134
rect 328810 399218 329046 399454
rect 328810 398898 329046 399134
rect 359530 399218 359766 399454
rect 359530 398898 359766 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 252010 367718 252246 367954
rect 252010 367398 252246 367634
rect 282730 367718 282966 367954
rect 282730 367398 282966 367634
rect 313450 367718 313686 367954
rect 313450 367398 313686 367634
rect 344170 367718 344406 367954
rect 344170 367398 344406 367634
rect 236650 363218 236886 363454
rect 236650 362898 236886 363134
rect 267370 363218 267606 363454
rect 267370 362898 267606 363134
rect 298090 363218 298326 363454
rect 298090 362898 298326 363134
rect 328810 363218 329046 363454
rect 328810 362898 329046 363134
rect 359530 363218 359766 363454
rect 359530 362898 359766 363134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 252010 331718 252246 331954
rect 252010 331398 252246 331634
rect 282730 331718 282966 331954
rect 282730 331398 282966 331634
rect 313450 331718 313686 331954
rect 313450 331398 313686 331634
rect 344170 331718 344406 331954
rect 344170 331398 344406 331634
rect 236650 327218 236886 327454
rect 236650 326898 236886 327134
rect 267370 327218 267606 327454
rect 267370 326898 267606 327134
rect 298090 327218 298326 327454
rect 298090 326898 298326 327134
rect 328810 327218 329046 327454
rect 328810 326898 329046 327134
rect 359530 327218 359766 327454
rect 359530 326898 359766 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 220328 223718 220564 223954
rect 220328 223398 220564 223634
rect 356056 223718 356292 223954
rect 356056 223398 356292 223634
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 187718 220564 187954
rect 220328 187398 220564 187634
rect 356056 187718 356292 187954
rect 356056 187398 356292 187634
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 213326 -7612 213562 -7376
rect 213646 -7612 213882 -7376
rect 213326 -7932 213562 -7696
rect 213646 -7932 213882 -7696
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -892 218062 -656
rect 218146 -892 218382 -656
rect 217826 -1212 218062 -976
rect 218146 -1212 218382 -976
rect 222326 -1852 222562 -1616
rect 222646 -1852 222882 -1616
rect 222326 -2172 222562 -1936
rect 222646 -2172 222882 -1936
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2812 227062 -2576
rect 227146 -2812 227382 -2576
rect 226826 -3132 227062 -2896
rect 227146 -3132 227382 -2896
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3772 231562 -3536
rect 231646 -3772 231882 -3536
rect 231326 -4092 231562 -3856
rect 231646 -4092 231882 -3856
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4732 236062 -4496
rect 236146 -4732 236382 -4496
rect 235826 -5052 236062 -4816
rect 236146 -5052 236382 -4816
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5692 240562 -5456
rect 240646 -5692 240882 -5456
rect 240326 -6012 240562 -5776
rect 240646 -6012 240882 -5776
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6652 245062 -6416
rect 245146 -6652 245382 -6416
rect 244826 -6972 245062 -6736
rect 245146 -6972 245382 -6736
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7612 249562 -7376
rect 249646 -7612 249882 -7376
rect 249326 -7932 249562 -7696
rect 249646 -7932 249882 -7696
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -892 254062 -656
rect 254146 -892 254382 -656
rect 253826 -1212 254062 -976
rect 254146 -1212 254382 -976
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1852 258562 -1616
rect 258646 -1852 258882 -1616
rect 258326 -2172 258562 -1936
rect 258646 -2172 258882 -1936
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2812 263062 -2576
rect 263146 -2812 263382 -2576
rect 262826 -3132 263062 -2896
rect 263146 -3132 263382 -2896
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3772 267562 -3536
rect 267646 -3772 267882 -3536
rect 267326 -4092 267562 -3856
rect 267646 -4092 267882 -3856
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4732 272062 -4496
rect 272146 -4732 272382 -4496
rect 271826 -5052 272062 -4816
rect 272146 -5052 272382 -4816
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5692 276562 -5456
rect 276646 -5692 276882 -5456
rect 276326 -6012 276562 -5776
rect 276646 -6012 276882 -5776
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6652 281062 -6416
rect 281146 -6652 281382 -6416
rect 280826 -6972 281062 -6736
rect 281146 -6972 281382 -6736
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7612 285562 -7376
rect 285646 -7612 285882 -7376
rect 285326 -7932 285562 -7696
rect 285646 -7932 285882 -7696
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -892 290062 -656
rect 290146 -892 290382 -656
rect 289826 -1212 290062 -976
rect 290146 -1212 290382 -976
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1852 294562 -1616
rect 294646 -1852 294882 -1616
rect 294326 -2172 294562 -1936
rect 294646 -2172 294882 -1936
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2812 299062 -2576
rect 299146 -2812 299382 -2576
rect 298826 -3132 299062 -2896
rect 299146 -3132 299382 -2896
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3772 303562 -3536
rect 303646 -3772 303882 -3536
rect 303326 -4092 303562 -3856
rect 303646 -4092 303882 -3856
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4732 308062 -4496
rect 308146 -4732 308382 -4496
rect 307826 -5052 308062 -4816
rect 308146 -5052 308382 -4816
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5692 312562 -5456
rect 312646 -5692 312882 -5456
rect 312326 -6012 312562 -5776
rect 312646 -6012 312882 -5776
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6652 317062 -6416
rect 317146 -6652 317382 -6416
rect 316826 -6972 317062 -6736
rect 317146 -6972 317382 -6736
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7612 321562 -7376
rect 321646 -7612 321882 -7376
rect 321326 -7932 321562 -7696
rect 321646 -7932 321882 -7696
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -892 326062 -656
rect 326146 -892 326382 -656
rect 325826 -1212 326062 -976
rect 326146 -1212 326382 -976
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1852 330562 -1616
rect 330646 -1852 330882 -1616
rect 330326 -2172 330562 -1936
rect 330646 -2172 330882 -1936
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2812 335062 -2576
rect 335146 -2812 335382 -2576
rect 334826 -3132 335062 -2896
rect 335146 -3132 335382 -2896
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3772 339562 -3536
rect 339646 -3772 339882 -3536
rect 339326 -4092 339562 -3856
rect 339646 -4092 339882 -3856
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4732 344062 -4496
rect 344146 -4732 344382 -4496
rect 343826 -5052 344062 -4816
rect 344146 -5052 344382 -4816
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5692 348562 -5456
rect 348646 -5692 348882 -5456
rect 348326 -6012 348562 -5776
rect 348646 -6012 348882 -5776
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6652 353062 -6416
rect 353146 -6652 353382 -6416
rect 352826 -6972 353062 -6736
rect 353146 -6972 353382 -6736
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 370826 706832 371062 707068
rect 371146 706832 371382 707068
rect 370826 706512 371062 706748
rect 371146 706512 371382 706748
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 357326 -7612 357562 -7376
rect 357646 -7612 357882 -7376
rect 357326 -7932 357562 -7696
rect 357646 -7932 357882 -7696
rect 361826 -892 362062 -656
rect 362146 -892 362382 -656
rect 361826 -1212 362062 -976
rect 362146 -1212 362382 -976
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 366326 -1852 366562 -1616
rect 366646 -1852 366882 -1616
rect 366326 -2172 366562 -1936
rect 366646 -2172 366882 -1936
rect 370826 -2812 371062 -2576
rect 371146 -2812 371382 -2576
rect 370826 -3132 371062 -2896
rect 371146 -3132 371382 -2896
rect 375326 707792 375562 708028
rect 375646 707792 375882 708028
rect 375326 707472 375562 707708
rect 375646 707472 375882 707708
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3772 375562 -3536
rect 375646 -3772 375882 -3536
rect 375326 -4092 375562 -3856
rect 375646 -4092 375882 -3856
rect 379826 708752 380062 708988
rect 380146 708752 380382 708988
rect 379826 708432 380062 708668
rect 380146 708432 380382 708668
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4732 380062 -4496
rect 380146 -4732 380382 -4496
rect 379826 -5052 380062 -4816
rect 380146 -5052 380382 -4816
rect 384326 709712 384562 709948
rect 384646 709712 384882 709948
rect 384326 709392 384562 709628
rect 384646 709392 384882 709628
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5692 384562 -5456
rect 384646 -5692 384882 -5456
rect 384326 -6012 384562 -5776
rect 384646 -6012 384882 -5776
rect 388826 710672 389062 710908
rect 389146 710672 389382 710908
rect 388826 710352 389062 710588
rect 389146 710352 389382 710588
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6652 389062 -6416
rect 389146 -6652 389382 -6416
rect 388826 -6972 389062 -6736
rect 389146 -6972 389382 -6736
rect 393326 711632 393562 711868
rect 393646 711632 393882 711868
rect 393326 711312 393562 711548
rect 393646 711312 393882 711548
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7612 393562 -7376
rect 393646 -7612 393882 -7376
rect 393326 -7932 393562 -7696
rect 393646 -7932 393882 -7696
rect 397826 704912 398062 705148
rect 398146 704912 398382 705148
rect 397826 704592 398062 704828
rect 398146 704592 398382 704828
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -892 398062 -656
rect 398146 -892 398382 -656
rect 397826 -1212 398062 -976
rect 398146 -1212 398382 -976
rect 402326 705872 402562 706108
rect 402646 705872 402882 706108
rect 402326 705552 402562 705788
rect 402646 705552 402882 705788
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1852 402562 -1616
rect 402646 -1852 402882 -1616
rect 402326 -2172 402562 -1936
rect 402646 -2172 402882 -1936
rect 406826 706832 407062 707068
rect 407146 706832 407382 707068
rect 406826 706512 407062 706748
rect 407146 706512 407382 706748
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2812 407062 -2576
rect 407146 -2812 407382 -2576
rect 406826 -3132 407062 -2896
rect 407146 -3132 407382 -2896
rect 411326 707792 411562 708028
rect 411646 707792 411882 708028
rect 411326 707472 411562 707708
rect 411646 707472 411882 707708
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3772 411562 -3536
rect 411646 -3772 411882 -3536
rect 411326 -4092 411562 -3856
rect 411646 -4092 411882 -3856
rect 415826 708752 416062 708988
rect 416146 708752 416382 708988
rect 415826 708432 416062 708668
rect 416146 708432 416382 708668
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4732 416062 -4496
rect 416146 -4732 416382 -4496
rect 415826 -5052 416062 -4816
rect 416146 -5052 416382 -4816
rect 420326 709712 420562 709948
rect 420646 709712 420882 709948
rect 420326 709392 420562 709628
rect 420646 709392 420882 709628
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5692 420562 -5456
rect 420646 -5692 420882 -5456
rect 420326 -6012 420562 -5776
rect 420646 -6012 420882 -5776
rect 424826 710672 425062 710908
rect 425146 710672 425382 710908
rect 424826 710352 425062 710588
rect 425146 710352 425382 710588
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6652 425062 -6416
rect 425146 -6652 425382 -6416
rect 424826 -6972 425062 -6736
rect 425146 -6972 425382 -6736
rect 429326 711632 429562 711868
rect 429646 711632 429882 711868
rect 429326 711312 429562 711548
rect 429646 711312 429882 711548
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7612 429562 -7376
rect 429646 -7612 429882 -7376
rect 429326 -7932 429562 -7696
rect 429646 -7932 429882 -7696
rect 433826 704912 434062 705148
rect 434146 704912 434382 705148
rect 433826 704592 434062 704828
rect 434146 704592 434382 704828
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -892 434062 -656
rect 434146 -892 434382 -656
rect 433826 -1212 434062 -976
rect 434146 -1212 434382 -976
rect 438326 705872 438562 706108
rect 438646 705872 438882 706108
rect 438326 705552 438562 705788
rect 438646 705552 438882 705788
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1852 438562 -1616
rect 438646 -1852 438882 -1616
rect 438326 -2172 438562 -1936
rect 438646 -2172 438882 -1936
rect 442826 706832 443062 707068
rect 443146 706832 443382 707068
rect 442826 706512 443062 706748
rect 443146 706512 443382 706748
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2812 443062 -2576
rect 443146 -2812 443382 -2576
rect 442826 -3132 443062 -2896
rect 443146 -3132 443382 -2896
rect 447326 707792 447562 708028
rect 447646 707792 447882 708028
rect 447326 707472 447562 707708
rect 447646 707472 447882 707708
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3772 447562 -3536
rect 447646 -3772 447882 -3536
rect 447326 -4092 447562 -3856
rect 447646 -4092 447882 -3856
rect 451826 708752 452062 708988
rect 452146 708752 452382 708988
rect 451826 708432 452062 708668
rect 452146 708432 452382 708668
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4732 452062 -4496
rect 452146 -4732 452382 -4496
rect 451826 -5052 452062 -4816
rect 452146 -5052 452382 -4816
rect 456326 709712 456562 709948
rect 456646 709712 456882 709948
rect 456326 709392 456562 709628
rect 456646 709392 456882 709628
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5692 456562 -5456
rect 456646 -5692 456882 -5456
rect 456326 -6012 456562 -5776
rect 456646 -6012 456882 -5776
rect 460826 710672 461062 710908
rect 461146 710672 461382 710908
rect 460826 710352 461062 710588
rect 461146 710352 461382 710588
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6652 461062 -6416
rect 461146 -6652 461382 -6416
rect 460826 -6972 461062 -6736
rect 461146 -6972 461382 -6736
rect 465326 711632 465562 711868
rect 465646 711632 465882 711868
rect 465326 711312 465562 711548
rect 465646 711312 465882 711548
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7612 465562 -7376
rect 465646 -7612 465882 -7376
rect 465326 -7932 465562 -7696
rect 465646 -7932 465882 -7696
rect 469826 704912 470062 705148
rect 470146 704912 470382 705148
rect 469826 704592 470062 704828
rect 470146 704592 470382 704828
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -892 470062 -656
rect 470146 -892 470382 -656
rect 469826 -1212 470062 -976
rect 470146 -1212 470382 -976
rect 474326 705872 474562 706108
rect 474646 705872 474882 706108
rect 474326 705552 474562 705788
rect 474646 705552 474882 705788
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1852 474562 -1616
rect 474646 -1852 474882 -1616
rect 474326 -2172 474562 -1936
rect 474646 -2172 474882 -1936
rect 478826 706832 479062 707068
rect 479146 706832 479382 707068
rect 478826 706512 479062 706748
rect 479146 706512 479382 706748
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2812 479062 -2576
rect 479146 -2812 479382 -2576
rect 478826 -3132 479062 -2896
rect 479146 -3132 479382 -2896
rect 483326 707792 483562 708028
rect 483646 707792 483882 708028
rect 483326 707472 483562 707708
rect 483646 707472 483882 707708
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3772 483562 -3536
rect 483646 -3772 483882 -3536
rect 483326 -4092 483562 -3856
rect 483646 -4092 483882 -3856
rect 487826 708752 488062 708988
rect 488146 708752 488382 708988
rect 487826 708432 488062 708668
rect 488146 708432 488382 708668
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4732 488062 -4496
rect 488146 -4732 488382 -4496
rect 487826 -5052 488062 -4816
rect 488146 -5052 488382 -4816
rect 492326 709712 492562 709948
rect 492646 709712 492882 709948
rect 492326 709392 492562 709628
rect 492646 709392 492882 709628
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5692 492562 -5456
rect 492646 -5692 492882 -5456
rect 492326 -6012 492562 -5776
rect 492646 -6012 492882 -5776
rect 496826 710672 497062 710908
rect 497146 710672 497382 710908
rect 496826 710352 497062 710588
rect 497146 710352 497382 710588
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6652 497062 -6416
rect 497146 -6652 497382 -6416
rect 496826 -6972 497062 -6736
rect 497146 -6972 497382 -6736
rect 501326 711632 501562 711868
rect 501646 711632 501882 711868
rect 501326 711312 501562 711548
rect 501646 711312 501882 711548
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7612 501562 -7376
rect 501646 -7612 501882 -7376
rect 501326 -7932 501562 -7696
rect 501646 -7932 501882 -7696
rect 505826 704912 506062 705148
rect 506146 704912 506382 705148
rect 505826 704592 506062 704828
rect 506146 704592 506382 704828
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -892 506062 -656
rect 506146 -892 506382 -656
rect 505826 -1212 506062 -976
rect 506146 -1212 506382 -976
rect 510326 705872 510562 706108
rect 510646 705872 510882 706108
rect 510326 705552 510562 705788
rect 510646 705552 510882 705788
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1852 510562 -1616
rect 510646 -1852 510882 -1616
rect 510326 -2172 510562 -1936
rect 510646 -2172 510882 -1936
rect 514826 706832 515062 707068
rect 515146 706832 515382 707068
rect 514826 706512 515062 706748
rect 515146 706512 515382 706748
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2812 515062 -2576
rect 515146 -2812 515382 -2576
rect 514826 -3132 515062 -2896
rect 515146 -3132 515382 -2896
rect 519326 707792 519562 708028
rect 519646 707792 519882 708028
rect 519326 707472 519562 707708
rect 519646 707472 519882 707708
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3772 519562 -3536
rect 519646 -3772 519882 -3536
rect 519326 -4092 519562 -3856
rect 519646 -4092 519882 -3856
rect 523826 708752 524062 708988
rect 524146 708752 524382 708988
rect 523826 708432 524062 708668
rect 524146 708432 524382 708668
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4732 524062 -4496
rect 524146 -4732 524382 -4496
rect 523826 -5052 524062 -4816
rect 524146 -5052 524382 -4816
rect 528326 709712 528562 709948
rect 528646 709712 528882 709948
rect 528326 709392 528562 709628
rect 528646 709392 528882 709628
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5692 528562 -5456
rect 528646 -5692 528882 -5456
rect 528326 -6012 528562 -5776
rect 528646 -6012 528882 -5776
rect 532826 710672 533062 710908
rect 533146 710672 533382 710908
rect 532826 710352 533062 710588
rect 533146 710352 533382 710588
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6652 533062 -6416
rect 533146 -6652 533382 -6416
rect 532826 -6972 533062 -6736
rect 533146 -6972 533382 -6736
rect 537326 711632 537562 711868
rect 537646 711632 537882 711868
rect 537326 711312 537562 711548
rect 537646 711312 537882 711548
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7612 537562 -7376
rect 537646 -7612 537882 -7376
rect 537326 -7932 537562 -7696
rect 537646 -7932 537882 -7696
rect 541826 704912 542062 705148
rect 542146 704912 542382 705148
rect 541826 704592 542062 704828
rect 542146 704592 542382 704828
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -892 542062 -656
rect 542146 -892 542382 -656
rect 541826 -1212 542062 -976
rect 542146 -1212 542382 -976
rect 546326 705872 546562 706108
rect 546646 705872 546882 706108
rect 546326 705552 546562 705788
rect 546646 705552 546882 705788
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1852 546562 -1616
rect 546646 -1852 546882 -1616
rect 546326 -2172 546562 -1936
rect 546646 -2172 546882 -1936
rect 550826 706832 551062 707068
rect 551146 706832 551382 707068
rect 550826 706512 551062 706748
rect 551146 706512 551382 706748
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2812 551062 -2576
rect 551146 -2812 551382 -2576
rect 550826 -3132 551062 -2896
rect 551146 -3132 551382 -2896
rect 555326 707792 555562 708028
rect 555646 707792 555882 708028
rect 555326 707472 555562 707708
rect 555646 707472 555882 707708
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3772 555562 -3536
rect 555646 -3772 555882 -3536
rect 555326 -4092 555562 -3856
rect 555646 -4092 555882 -3856
rect 559826 708752 560062 708988
rect 560146 708752 560382 708988
rect 559826 708432 560062 708668
rect 560146 708432 560382 708668
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4732 560062 -4496
rect 560146 -4732 560382 -4496
rect 559826 -5052 560062 -4816
rect 560146 -5052 560382 -4816
rect 564326 709712 564562 709948
rect 564646 709712 564882 709948
rect 564326 709392 564562 709628
rect 564646 709392 564882 709628
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5692 564562 -5456
rect 564646 -5692 564882 -5456
rect 564326 -6012 564562 -5776
rect 564646 -6012 564882 -5776
rect 568826 710672 569062 710908
rect 569146 710672 569382 710908
rect 568826 710352 569062 710588
rect 569146 710352 569382 710588
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6652 569062 -6416
rect 569146 -6652 569382 -6416
rect 568826 -6972 569062 -6736
rect 569146 -6972 569382 -6736
rect 573326 711632 573562 711868
rect 573646 711632 573882 711868
rect 573326 711312 573562 711548
rect 573646 711312 573882 711548
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7612 573562 -7376
rect 573646 -7612 573882 -7376
rect 573326 -7932 573562 -7696
rect 573646 -7932 573882 -7696
rect 577826 704912 578062 705148
rect 578146 704912 578382 705148
rect 577826 704592 578062 704828
rect 578146 704592 578382 704828
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -892 578062 -656
rect 578146 -892 578382 -656
rect 577826 -1212 578062 -976
rect 578146 -1212 578382 -976
rect 592372 711632 592608 711868
rect 592692 711632 592928 711868
rect 592372 711312 592608 711548
rect 592692 711312 592928 711548
rect 591412 710672 591648 710908
rect 591732 710672 591968 710908
rect 591412 710352 591648 710588
rect 591732 710352 591968 710588
rect 590452 709712 590688 709948
rect 590772 709712 591008 709948
rect 590452 709392 590688 709628
rect 590772 709392 591008 709628
rect 589492 708752 589728 708988
rect 589812 708752 590048 708988
rect 589492 708432 589728 708668
rect 589812 708432 590048 708668
rect 588532 707792 588768 708028
rect 588852 707792 589088 708028
rect 588532 707472 588768 707708
rect 588852 707472 589088 707708
rect 587572 706832 587808 707068
rect 587892 706832 588128 707068
rect 587572 706512 587808 706748
rect 587892 706512 588128 706748
rect 582326 705872 582562 706108
rect 582646 705872 582882 706108
rect 582326 705552 582562 705788
rect 582646 705552 582882 705788
rect 586612 705872 586848 706108
rect 586932 705872 587168 706108
rect 586612 705552 586848 705788
rect 586932 705552 587168 705788
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585652 704912 585888 705148
rect 585972 704912 586208 705148
rect 585652 704592 585888 704828
rect 585972 704592 586208 704828
rect 585652 687218 585888 687454
rect 585972 687218 586208 687454
rect 585652 686898 585888 687134
rect 585972 686898 586208 687134
rect 585652 651218 585888 651454
rect 585972 651218 586208 651454
rect 585652 650898 585888 651134
rect 585972 650898 586208 651134
rect 585652 615218 585888 615454
rect 585972 615218 586208 615454
rect 585652 614898 585888 615134
rect 585972 614898 586208 615134
rect 585652 579218 585888 579454
rect 585972 579218 586208 579454
rect 585652 578898 585888 579134
rect 585972 578898 586208 579134
rect 585652 543218 585888 543454
rect 585972 543218 586208 543454
rect 585652 542898 585888 543134
rect 585972 542898 586208 543134
rect 585652 507218 585888 507454
rect 585972 507218 586208 507454
rect 585652 506898 585888 507134
rect 585972 506898 586208 507134
rect 585652 471218 585888 471454
rect 585972 471218 586208 471454
rect 585652 470898 585888 471134
rect 585972 470898 586208 471134
rect 585652 435218 585888 435454
rect 585972 435218 586208 435454
rect 585652 434898 585888 435134
rect 585972 434898 586208 435134
rect 585652 399218 585888 399454
rect 585972 399218 586208 399454
rect 585652 398898 585888 399134
rect 585972 398898 586208 399134
rect 585652 363218 585888 363454
rect 585972 363218 586208 363454
rect 585652 362898 585888 363134
rect 585972 362898 586208 363134
rect 585652 327218 585888 327454
rect 585972 327218 586208 327454
rect 585652 326898 585888 327134
rect 585972 326898 586208 327134
rect 585652 291218 585888 291454
rect 585972 291218 586208 291454
rect 585652 290898 585888 291134
rect 585972 290898 586208 291134
rect 585652 255218 585888 255454
rect 585972 255218 586208 255454
rect 585652 254898 585888 255134
rect 585972 254898 586208 255134
rect 585652 219218 585888 219454
rect 585972 219218 586208 219454
rect 585652 218898 585888 219134
rect 585972 218898 586208 219134
rect 585652 183218 585888 183454
rect 585972 183218 586208 183454
rect 585652 182898 585888 183134
rect 585972 182898 586208 183134
rect 585652 147218 585888 147454
rect 585972 147218 586208 147454
rect 585652 146898 585888 147134
rect 585972 146898 586208 147134
rect 585652 111218 585888 111454
rect 585972 111218 586208 111454
rect 585652 110898 585888 111134
rect 585972 110898 586208 111134
rect 585652 75218 585888 75454
rect 585972 75218 586208 75454
rect 585652 74898 585888 75134
rect 585972 74898 586208 75134
rect 585652 39218 585888 39454
rect 585972 39218 586208 39454
rect 585652 38898 585888 39134
rect 585972 38898 586208 39134
rect 585652 3218 585888 3454
rect 585972 3218 586208 3454
rect 585652 2898 585888 3134
rect 585972 2898 586208 3134
rect 585652 -892 585888 -656
rect 585972 -892 586208 -656
rect 585652 -1212 585888 -976
rect 585972 -1212 586208 -976
rect 586612 691718 586848 691954
rect 586932 691718 587168 691954
rect 586612 691398 586848 691634
rect 586932 691398 587168 691634
rect 586612 655718 586848 655954
rect 586932 655718 587168 655954
rect 586612 655398 586848 655634
rect 586932 655398 587168 655634
rect 586612 619718 586848 619954
rect 586932 619718 587168 619954
rect 586612 619398 586848 619634
rect 586932 619398 587168 619634
rect 586612 583718 586848 583954
rect 586932 583718 587168 583954
rect 586612 583398 586848 583634
rect 586932 583398 587168 583634
rect 586612 547718 586848 547954
rect 586932 547718 587168 547954
rect 586612 547398 586848 547634
rect 586932 547398 587168 547634
rect 586612 511718 586848 511954
rect 586932 511718 587168 511954
rect 586612 511398 586848 511634
rect 586932 511398 587168 511634
rect 586612 475718 586848 475954
rect 586932 475718 587168 475954
rect 586612 475398 586848 475634
rect 586932 475398 587168 475634
rect 586612 439718 586848 439954
rect 586932 439718 587168 439954
rect 586612 439398 586848 439634
rect 586932 439398 587168 439634
rect 586612 403718 586848 403954
rect 586932 403718 587168 403954
rect 586612 403398 586848 403634
rect 586932 403398 587168 403634
rect 586612 367718 586848 367954
rect 586932 367718 587168 367954
rect 586612 367398 586848 367634
rect 586932 367398 587168 367634
rect 586612 331718 586848 331954
rect 586932 331718 587168 331954
rect 586612 331398 586848 331634
rect 586932 331398 587168 331634
rect 586612 295718 586848 295954
rect 586932 295718 587168 295954
rect 586612 295398 586848 295634
rect 586932 295398 587168 295634
rect 586612 259718 586848 259954
rect 586932 259718 587168 259954
rect 586612 259398 586848 259634
rect 586932 259398 587168 259634
rect 586612 223718 586848 223954
rect 586932 223718 587168 223954
rect 586612 223398 586848 223634
rect 586932 223398 587168 223634
rect 586612 187718 586848 187954
rect 586932 187718 587168 187954
rect 586612 187398 586848 187634
rect 586932 187398 587168 187634
rect 586612 151718 586848 151954
rect 586932 151718 587168 151954
rect 586612 151398 586848 151634
rect 586932 151398 587168 151634
rect 586612 115718 586848 115954
rect 586932 115718 587168 115954
rect 586612 115398 586848 115634
rect 586932 115398 587168 115634
rect 586612 79718 586848 79954
rect 586932 79718 587168 79954
rect 586612 79398 586848 79634
rect 586932 79398 587168 79634
rect 586612 43718 586848 43954
rect 586932 43718 587168 43954
rect 586612 43398 586848 43634
rect 586932 43398 587168 43634
rect 586612 7718 586848 7954
rect 586932 7718 587168 7954
rect 586612 7398 586848 7634
rect 586932 7398 587168 7634
rect 582326 -1852 582562 -1616
rect 582646 -1852 582882 -1616
rect 582326 -2172 582562 -1936
rect 582646 -2172 582882 -1936
rect 586612 -1852 586848 -1616
rect 586932 -1852 587168 -1616
rect 586612 -2172 586848 -1936
rect 586932 -2172 587168 -1936
rect 587572 696218 587808 696454
rect 587892 696218 588128 696454
rect 587572 695898 587808 696134
rect 587892 695898 588128 696134
rect 587572 660218 587808 660454
rect 587892 660218 588128 660454
rect 587572 659898 587808 660134
rect 587892 659898 588128 660134
rect 587572 624218 587808 624454
rect 587892 624218 588128 624454
rect 587572 623898 587808 624134
rect 587892 623898 588128 624134
rect 587572 588218 587808 588454
rect 587892 588218 588128 588454
rect 587572 587898 587808 588134
rect 587892 587898 588128 588134
rect 587572 552218 587808 552454
rect 587892 552218 588128 552454
rect 587572 551898 587808 552134
rect 587892 551898 588128 552134
rect 587572 516218 587808 516454
rect 587892 516218 588128 516454
rect 587572 515898 587808 516134
rect 587892 515898 588128 516134
rect 587572 480218 587808 480454
rect 587892 480218 588128 480454
rect 587572 479898 587808 480134
rect 587892 479898 588128 480134
rect 587572 444218 587808 444454
rect 587892 444218 588128 444454
rect 587572 443898 587808 444134
rect 587892 443898 588128 444134
rect 587572 408218 587808 408454
rect 587892 408218 588128 408454
rect 587572 407898 587808 408134
rect 587892 407898 588128 408134
rect 587572 372218 587808 372454
rect 587892 372218 588128 372454
rect 587572 371898 587808 372134
rect 587892 371898 588128 372134
rect 587572 336218 587808 336454
rect 587892 336218 588128 336454
rect 587572 335898 587808 336134
rect 587892 335898 588128 336134
rect 587572 300218 587808 300454
rect 587892 300218 588128 300454
rect 587572 299898 587808 300134
rect 587892 299898 588128 300134
rect 587572 264218 587808 264454
rect 587892 264218 588128 264454
rect 587572 263898 587808 264134
rect 587892 263898 588128 264134
rect 587572 228218 587808 228454
rect 587892 228218 588128 228454
rect 587572 227898 587808 228134
rect 587892 227898 588128 228134
rect 587572 192218 587808 192454
rect 587892 192218 588128 192454
rect 587572 191898 587808 192134
rect 587892 191898 588128 192134
rect 587572 156218 587808 156454
rect 587892 156218 588128 156454
rect 587572 155898 587808 156134
rect 587892 155898 588128 156134
rect 587572 120218 587808 120454
rect 587892 120218 588128 120454
rect 587572 119898 587808 120134
rect 587892 119898 588128 120134
rect 587572 84218 587808 84454
rect 587892 84218 588128 84454
rect 587572 83898 587808 84134
rect 587892 83898 588128 84134
rect 587572 48218 587808 48454
rect 587892 48218 588128 48454
rect 587572 47898 587808 48134
rect 587892 47898 588128 48134
rect 587572 12218 587808 12454
rect 587892 12218 588128 12454
rect 587572 11898 587808 12134
rect 587892 11898 588128 12134
rect 587572 -2812 587808 -2576
rect 587892 -2812 588128 -2576
rect 587572 -3132 587808 -2896
rect 587892 -3132 588128 -2896
rect 588532 700718 588768 700954
rect 588852 700718 589088 700954
rect 588532 700398 588768 700634
rect 588852 700398 589088 700634
rect 588532 664718 588768 664954
rect 588852 664718 589088 664954
rect 588532 664398 588768 664634
rect 588852 664398 589088 664634
rect 588532 628718 588768 628954
rect 588852 628718 589088 628954
rect 588532 628398 588768 628634
rect 588852 628398 589088 628634
rect 588532 592718 588768 592954
rect 588852 592718 589088 592954
rect 588532 592398 588768 592634
rect 588852 592398 589088 592634
rect 588532 556718 588768 556954
rect 588852 556718 589088 556954
rect 588532 556398 588768 556634
rect 588852 556398 589088 556634
rect 588532 520718 588768 520954
rect 588852 520718 589088 520954
rect 588532 520398 588768 520634
rect 588852 520398 589088 520634
rect 588532 484718 588768 484954
rect 588852 484718 589088 484954
rect 588532 484398 588768 484634
rect 588852 484398 589088 484634
rect 588532 448718 588768 448954
rect 588852 448718 589088 448954
rect 588532 448398 588768 448634
rect 588852 448398 589088 448634
rect 588532 412718 588768 412954
rect 588852 412718 589088 412954
rect 588532 412398 588768 412634
rect 588852 412398 589088 412634
rect 588532 376718 588768 376954
rect 588852 376718 589088 376954
rect 588532 376398 588768 376634
rect 588852 376398 589088 376634
rect 588532 340718 588768 340954
rect 588852 340718 589088 340954
rect 588532 340398 588768 340634
rect 588852 340398 589088 340634
rect 588532 304718 588768 304954
rect 588852 304718 589088 304954
rect 588532 304398 588768 304634
rect 588852 304398 589088 304634
rect 588532 268718 588768 268954
rect 588852 268718 589088 268954
rect 588532 268398 588768 268634
rect 588852 268398 589088 268634
rect 588532 232718 588768 232954
rect 588852 232718 589088 232954
rect 588532 232398 588768 232634
rect 588852 232398 589088 232634
rect 588532 196718 588768 196954
rect 588852 196718 589088 196954
rect 588532 196398 588768 196634
rect 588852 196398 589088 196634
rect 588532 160718 588768 160954
rect 588852 160718 589088 160954
rect 588532 160398 588768 160634
rect 588852 160398 589088 160634
rect 588532 124718 588768 124954
rect 588852 124718 589088 124954
rect 588532 124398 588768 124634
rect 588852 124398 589088 124634
rect 588532 88718 588768 88954
rect 588852 88718 589088 88954
rect 588532 88398 588768 88634
rect 588852 88398 589088 88634
rect 588532 52718 588768 52954
rect 588852 52718 589088 52954
rect 588532 52398 588768 52634
rect 588852 52398 589088 52634
rect 588532 16718 588768 16954
rect 588852 16718 589088 16954
rect 588532 16398 588768 16634
rect 588852 16398 589088 16634
rect 588532 -3772 588768 -3536
rect 588852 -3772 589088 -3536
rect 588532 -4092 588768 -3856
rect 588852 -4092 589088 -3856
rect 589492 669218 589728 669454
rect 589812 669218 590048 669454
rect 589492 668898 589728 669134
rect 589812 668898 590048 669134
rect 589492 633218 589728 633454
rect 589812 633218 590048 633454
rect 589492 632898 589728 633134
rect 589812 632898 590048 633134
rect 589492 597218 589728 597454
rect 589812 597218 590048 597454
rect 589492 596898 589728 597134
rect 589812 596898 590048 597134
rect 589492 561218 589728 561454
rect 589812 561218 590048 561454
rect 589492 560898 589728 561134
rect 589812 560898 590048 561134
rect 589492 525218 589728 525454
rect 589812 525218 590048 525454
rect 589492 524898 589728 525134
rect 589812 524898 590048 525134
rect 589492 489218 589728 489454
rect 589812 489218 590048 489454
rect 589492 488898 589728 489134
rect 589812 488898 590048 489134
rect 589492 453218 589728 453454
rect 589812 453218 590048 453454
rect 589492 452898 589728 453134
rect 589812 452898 590048 453134
rect 589492 417218 589728 417454
rect 589812 417218 590048 417454
rect 589492 416898 589728 417134
rect 589812 416898 590048 417134
rect 589492 381218 589728 381454
rect 589812 381218 590048 381454
rect 589492 380898 589728 381134
rect 589812 380898 590048 381134
rect 589492 345218 589728 345454
rect 589812 345218 590048 345454
rect 589492 344898 589728 345134
rect 589812 344898 590048 345134
rect 589492 309218 589728 309454
rect 589812 309218 590048 309454
rect 589492 308898 589728 309134
rect 589812 308898 590048 309134
rect 589492 273218 589728 273454
rect 589812 273218 590048 273454
rect 589492 272898 589728 273134
rect 589812 272898 590048 273134
rect 589492 237218 589728 237454
rect 589812 237218 590048 237454
rect 589492 236898 589728 237134
rect 589812 236898 590048 237134
rect 589492 201218 589728 201454
rect 589812 201218 590048 201454
rect 589492 200898 589728 201134
rect 589812 200898 590048 201134
rect 589492 165218 589728 165454
rect 589812 165218 590048 165454
rect 589492 164898 589728 165134
rect 589812 164898 590048 165134
rect 589492 129218 589728 129454
rect 589812 129218 590048 129454
rect 589492 128898 589728 129134
rect 589812 128898 590048 129134
rect 589492 93218 589728 93454
rect 589812 93218 590048 93454
rect 589492 92898 589728 93134
rect 589812 92898 590048 93134
rect 589492 57218 589728 57454
rect 589812 57218 590048 57454
rect 589492 56898 589728 57134
rect 589812 56898 590048 57134
rect 589492 21218 589728 21454
rect 589812 21218 590048 21454
rect 589492 20898 589728 21134
rect 589812 20898 590048 21134
rect 589492 -4732 589728 -4496
rect 589812 -4732 590048 -4496
rect 589492 -5052 589728 -4816
rect 589812 -5052 590048 -4816
rect 590452 673718 590688 673954
rect 590772 673718 591008 673954
rect 590452 673398 590688 673634
rect 590772 673398 591008 673634
rect 590452 637718 590688 637954
rect 590772 637718 591008 637954
rect 590452 637398 590688 637634
rect 590772 637398 591008 637634
rect 590452 601718 590688 601954
rect 590772 601718 591008 601954
rect 590452 601398 590688 601634
rect 590772 601398 591008 601634
rect 590452 565718 590688 565954
rect 590772 565718 591008 565954
rect 590452 565398 590688 565634
rect 590772 565398 591008 565634
rect 590452 529718 590688 529954
rect 590772 529718 591008 529954
rect 590452 529398 590688 529634
rect 590772 529398 591008 529634
rect 590452 493718 590688 493954
rect 590772 493718 591008 493954
rect 590452 493398 590688 493634
rect 590772 493398 591008 493634
rect 590452 457718 590688 457954
rect 590772 457718 591008 457954
rect 590452 457398 590688 457634
rect 590772 457398 591008 457634
rect 590452 421718 590688 421954
rect 590772 421718 591008 421954
rect 590452 421398 590688 421634
rect 590772 421398 591008 421634
rect 590452 385718 590688 385954
rect 590772 385718 591008 385954
rect 590452 385398 590688 385634
rect 590772 385398 591008 385634
rect 590452 349718 590688 349954
rect 590772 349718 591008 349954
rect 590452 349398 590688 349634
rect 590772 349398 591008 349634
rect 590452 313718 590688 313954
rect 590772 313718 591008 313954
rect 590452 313398 590688 313634
rect 590772 313398 591008 313634
rect 590452 277718 590688 277954
rect 590772 277718 591008 277954
rect 590452 277398 590688 277634
rect 590772 277398 591008 277634
rect 590452 241718 590688 241954
rect 590772 241718 591008 241954
rect 590452 241398 590688 241634
rect 590772 241398 591008 241634
rect 590452 205718 590688 205954
rect 590772 205718 591008 205954
rect 590452 205398 590688 205634
rect 590772 205398 591008 205634
rect 590452 169718 590688 169954
rect 590772 169718 591008 169954
rect 590452 169398 590688 169634
rect 590772 169398 591008 169634
rect 590452 133718 590688 133954
rect 590772 133718 591008 133954
rect 590452 133398 590688 133634
rect 590772 133398 591008 133634
rect 590452 97718 590688 97954
rect 590772 97718 591008 97954
rect 590452 97398 590688 97634
rect 590772 97398 591008 97634
rect 590452 61718 590688 61954
rect 590772 61718 591008 61954
rect 590452 61398 590688 61634
rect 590772 61398 591008 61634
rect 590452 25718 590688 25954
rect 590772 25718 591008 25954
rect 590452 25398 590688 25634
rect 590772 25398 591008 25634
rect 590452 -5692 590688 -5456
rect 590772 -5692 591008 -5456
rect 590452 -6012 590688 -5776
rect 590772 -6012 591008 -5776
rect 591412 678218 591648 678454
rect 591732 678218 591968 678454
rect 591412 677898 591648 678134
rect 591732 677898 591968 678134
rect 591412 642218 591648 642454
rect 591732 642218 591968 642454
rect 591412 641898 591648 642134
rect 591732 641898 591968 642134
rect 591412 606218 591648 606454
rect 591732 606218 591968 606454
rect 591412 605898 591648 606134
rect 591732 605898 591968 606134
rect 591412 570218 591648 570454
rect 591732 570218 591968 570454
rect 591412 569898 591648 570134
rect 591732 569898 591968 570134
rect 591412 534218 591648 534454
rect 591732 534218 591968 534454
rect 591412 533898 591648 534134
rect 591732 533898 591968 534134
rect 591412 498218 591648 498454
rect 591732 498218 591968 498454
rect 591412 497898 591648 498134
rect 591732 497898 591968 498134
rect 591412 462218 591648 462454
rect 591732 462218 591968 462454
rect 591412 461898 591648 462134
rect 591732 461898 591968 462134
rect 591412 426218 591648 426454
rect 591732 426218 591968 426454
rect 591412 425898 591648 426134
rect 591732 425898 591968 426134
rect 591412 390218 591648 390454
rect 591732 390218 591968 390454
rect 591412 389898 591648 390134
rect 591732 389898 591968 390134
rect 591412 354218 591648 354454
rect 591732 354218 591968 354454
rect 591412 353898 591648 354134
rect 591732 353898 591968 354134
rect 591412 318218 591648 318454
rect 591732 318218 591968 318454
rect 591412 317898 591648 318134
rect 591732 317898 591968 318134
rect 591412 282218 591648 282454
rect 591732 282218 591968 282454
rect 591412 281898 591648 282134
rect 591732 281898 591968 282134
rect 591412 246218 591648 246454
rect 591732 246218 591968 246454
rect 591412 245898 591648 246134
rect 591732 245898 591968 246134
rect 591412 210218 591648 210454
rect 591732 210218 591968 210454
rect 591412 209898 591648 210134
rect 591732 209898 591968 210134
rect 591412 174218 591648 174454
rect 591732 174218 591968 174454
rect 591412 173898 591648 174134
rect 591732 173898 591968 174134
rect 591412 138218 591648 138454
rect 591732 138218 591968 138454
rect 591412 137898 591648 138134
rect 591732 137898 591968 138134
rect 591412 102218 591648 102454
rect 591732 102218 591968 102454
rect 591412 101898 591648 102134
rect 591732 101898 591968 102134
rect 591412 66218 591648 66454
rect 591732 66218 591968 66454
rect 591412 65898 591648 66134
rect 591732 65898 591968 66134
rect 591412 30218 591648 30454
rect 591732 30218 591968 30454
rect 591412 29898 591648 30134
rect 591732 29898 591968 30134
rect 591412 -6652 591648 -6416
rect 591732 -6652 591968 -6416
rect 591412 -6972 591648 -6736
rect 591732 -6972 591968 -6736
rect 592372 682718 592608 682954
rect 592692 682718 592928 682954
rect 592372 682398 592608 682634
rect 592692 682398 592928 682634
rect 592372 646718 592608 646954
rect 592692 646718 592928 646954
rect 592372 646398 592608 646634
rect 592692 646398 592928 646634
rect 592372 610718 592608 610954
rect 592692 610718 592928 610954
rect 592372 610398 592608 610634
rect 592692 610398 592928 610634
rect 592372 574718 592608 574954
rect 592692 574718 592928 574954
rect 592372 574398 592608 574634
rect 592692 574398 592928 574634
rect 592372 538718 592608 538954
rect 592692 538718 592928 538954
rect 592372 538398 592608 538634
rect 592692 538398 592928 538634
rect 592372 502718 592608 502954
rect 592692 502718 592928 502954
rect 592372 502398 592608 502634
rect 592692 502398 592928 502634
rect 592372 466718 592608 466954
rect 592692 466718 592928 466954
rect 592372 466398 592608 466634
rect 592692 466398 592928 466634
rect 592372 430718 592608 430954
rect 592692 430718 592928 430954
rect 592372 430398 592608 430634
rect 592692 430398 592928 430634
rect 592372 394718 592608 394954
rect 592692 394718 592928 394954
rect 592372 394398 592608 394634
rect 592692 394398 592928 394634
rect 592372 358718 592608 358954
rect 592692 358718 592928 358954
rect 592372 358398 592608 358634
rect 592692 358398 592928 358634
rect 592372 322718 592608 322954
rect 592692 322718 592928 322954
rect 592372 322398 592608 322634
rect 592692 322398 592928 322634
rect 592372 286718 592608 286954
rect 592692 286718 592928 286954
rect 592372 286398 592608 286634
rect 592692 286398 592928 286634
rect 592372 250718 592608 250954
rect 592692 250718 592928 250954
rect 592372 250398 592608 250634
rect 592692 250398 592928 250634
rect 592372 214718 592608 214954
rect 592692 214718 592928 214954
rect 592372 214398 592608 214634
rect 592692 214398 592928 214634
rect 592372 178718 592608 178954
rect 592692 178718 592928 178954
rect 592372 178398 592608 178634
rect 592692 178398 592928 178634
rect 592372 142718 592608 142954
rect 592692 142718 592928 142954
rect 592372 142398 592608 142634
rect 592692 142398 592928 142634
rect 592372 106718 592608 106954
rect 592692 106718 592928 106954
rect 592372 106398 592608 106634
rect 592692 106398 592928 106634
rect 592372 70718 592608 70954
rect 592692 70718 592928 70954
rect 592372 70398 592608 70634
rect 592692 70398 592928 70634
rect 592372 34718 592608 34954
rect 592692 34718 592928 34954
rect 592372 34398 592608 34634
rect 592692 34398 592928 34634
rect 592372 -7612 592608 -7376
rect 592692 -7612 592928 -7376
rect 592372 -7932 592608 -7696
rect 592692 -7932 592928 -7696
<< metal5 >>
rect -9036 711868 592960 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect -9036 711548 592960 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect -9036 711280 592960 711312
rect -8076 710908 592000 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect -8076 710588 592000 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect -8076 710320 592000 710352
rect -7116 709948 591040 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect -7116 709628 591040 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect -7116 709360 591040 709392
rect -6156 708988 590080 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect -6156 708668 590080 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect -6156 708400 590080 708432
rect -5196 708028 589120 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect -5196 707708 589120 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect -5196 707440 589120 707472
rect -4236 707068 588160 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect -4236 706748 588160 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect -4236 706480 588160 706512
rect -3276 706108 587200 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect -3276 705788 587200 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect -3276 705520 587200 705552
rect -2316 705148 586240 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect -2316 704828 586240 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect -2316 704560 586240 704592
rect -9036 700954 592960 700986
rect -9036 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 592960 700954
rect -9036 700634 592960 700718
rect -9036 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 592960 700634
rect -9036 700366 592960 700398
rect -9036 696454 592960 696486
rect -9036 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 592960 696454
rect -9036 696134 592960 696218
rect -9036 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 592960 696134
rect -9036 695866 592960 695898
rect -9036 691954 592960 691986
rect -9036 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 592960 691954
rect -9036 691634 592960 691718
rect -9036 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 592960 691634
rect -9036 691366 592960 691398
rect -9036 687454 592960 687486
rect -9036 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 592960 687454
rect -9036 687134 592960 687218
rect -9036 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 592960 687134
rect -9036 686866 592960 686898
rect -9036 682954 592960 682986
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect -9036 682634 592960 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect -9036 682366 592960 682398
rect -9036 678454 592960 678486
rect -9036 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592960 678454
rect -9036 678134 592960 678218
rect -9036 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592960 678134
rect -9036 677866 592960 677898
rect -9036 673954 592960 673986
rect -9036 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 592960 673954
rect -9036 673634 592960 673718
rect -9036 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 592960 673634
rect -9036 673366 592960 673398
rect -9036 669454 592960 669486
rect -9036 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 592960 669454
rect -9036 669134 592960 669218
rect -9036 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 592960 669134
rect -9036 668866 592960 668898
rect -9036 664954 592960 664986
rect -9036 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 592960 664954
rect -9036 664634 592960 664718
rect -9036 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 592960 664634
rect -9036 664366 592960 664398
rect -9036 660454 592960 660486
rect -9036 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 592960 660454
rect -9036 660134 592960 660218
rect -9036 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 592960 660134
rect -9036 659866 592960 659898
rect -9036 655954 592960 655986
rect -9036 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 592960 655954
rect -9036 655634 592960 655718
rect -9036 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 592960 655634
rect -9036 655366 592960 655398
rect -9036 651454 592960 651486
rect -9036 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 592960 651454
rect -9036 651134 592960 651218
rect -9036 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 592960 651134
rect -9036 650866 592960 650898
rect -9036 646954 592960 646986
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect -9036 646634 592960 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect -9036 646366 592960 646398
rect -9036 642454 592960 642486
rect -9036 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592960 642454
rect -9036 642134 592960 642218
rect -9036 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592960 642134
rect -9036 641866 592960 641898
rect -9036 637954 592960 637986
rect -9036 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 592960 637954
rect -9036 637634 592960 637718
rect -9036 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 592960 637634
rect -9036 637366 592960 637398
rect -9036 633454 592960 633486
rect -9036 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 592960 633454
rect -9036 633134 592960 633218
rect -9036 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 592960 633134
rect -9036 632866 592960 632898
rect -9036 628954 592960 628986
rect -9036 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 592960 628954
rect -9036 628634 592960 628718
rect -9036 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 592960 628634
rect -9036 628366 592960 628398
rect -9036 624454 592960 624486
rect -9036 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 592960 624454
rect -9036 624134 592960 624218
rect -9036 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 592960 624134
rect -9036 623866 592960 623898
rect -9036 619954 592960 619986
rect -9036 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 592960 619954
rect -9036 619634 592960 619718
rect -9036 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 592960 619634
rect -9036 619366 592960 619398
rect -9036 615454 592960 615486
rect -9036 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 592960 615454
rect -9036 615134 592960 615218
rect -9036 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 592960 615134
rect -9036 614866 592960 614898
rect -9036 610954 592960 610986
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect -9036 610634 592960 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect -9036 610366 592960 610398
rect -9036 606454 592960 606486
rect -9036 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592960 606454
rect -9036 606134 592960 606218
rect -9036 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592960 606134
rect -9036 605866 592960 605898
rect -9036 601954 592960 601986
rect -9036 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 592960 601954
rect -9036 601634 592960 601718
rect -9036 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 592960 601634
rect -9036 601366 592960 601398
rect -9036 597454 592960 597486
rect -9036 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 592960 597454
rect -9036 597134 592960 597218
rect -9036 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 592960 597134
rect -9036 596866 592960 596898
rect -9036 592954 592960 592986
rect -9036 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 592960 592954
rect -9036 592634 592960 592718
rect -9036 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 592960 592634
rect -9036 592366 592960 592398
rect -9036 588454 592960 588486
rect -9036 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 592960 588454
rect -9036 588134 592960 588218
rect -9036 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 592960 588134
rect -9036 587866 592960 587898
rect -9036 583954 592960 583986
rect -9036 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 592960 583954
rect -9036 583634 592960 583718
rect -9036 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 592960 583634
rect -9036 583366 592960 583398
rect -9036 579454 592960 579486
rect -9036 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 592960 579454
rect -9036 579134 592960 579218
rect -9036 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 592960 579134
rect -9036 578866 592960 578898
rect -9036 574954 592960 574986
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect -9036 574634 592960 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect -9036 574366 592960 574398
rect -9036 570454 592960 570486
rect -9036 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592960 570454
rect -9036 570134 592960 570218
rect -9036 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592960 570134
rect -9036 569866 592960 569898
rect -9036 565954 592960 565986
rect -9036 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 592960 565954
rect -9036 565634 592960 565718
rect -9036 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 592960 565634
rect -9036 565366 592960 565398
rect -9036 561454 592960 561486
rect -9036 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 592960 561454
rect -9036 561134 592960 561218
rect -9036 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 592960 561134
rect -9036 560866 592960 560898
rect -9036 556954 592960 556986
rect -9036 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 592960 556954
rect -9036 556634 592960 556718
rect -9036 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 592960 556634
rect -9036 556366 592960 556398
rect -9036 552454 592960 552486
rect -9036 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 592960 552454
rect -9036 552134 592960 552218
rect -9036 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 592960 552134
rect -9036 551866 592960 551898
rect -9036 547954 592960 547986
rect -9036 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 592960 547954
rect -9036 547634 592960 547718
rect -9036 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 592960 547634
rect -9036 547366 592960 547398
rect -9036 543454 592960 543486
rect -9036 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 592960 543454
rect -9036 543134 592960 543218
rect -9036 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 592960 543134
rect -9036 542866 592960 542898
rect -9036 538954 592960 538986
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect -9036 538634 592960 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect -9036 538366 592960 538398
rect -9036 534454 592960 534486
rect -9036 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592960 534454
rect -9036 534134 592960 534218
rect -9036 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592960 534134
rect -9036 533866 592960 533898
rect -9036 529954 592960 529986
rect -9036 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 592960 529954
rect -9036 529634 592960 529718
rect -9036 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 592960 529634
rect -9036 529366 592960 529398
rect -9036 525454 592960 525486
rect -9036 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 592960 525454
rect -9036 525134 592960 525218
rect -9036 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 592960 525134
rect -9036 524866 592960 524898
rect -9036 520954 592960 520986
rect -9036 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 592960 520954
rect -9036 520634 592960 520718
rect -9036 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 592960 520634
rect -9036 520366 592960 520398
rect -9036 516454 592960 516486
rect -9036 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 592960 516454
rect -9036 516134 592960 516218
rect -9036 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 592960 516134
rect -9036 515866 592960 515898
rect -9036 511954 592960 511986
rect -9036 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 592960 511954
rect -9036 511634 592960 511718
rect -9036 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 592960 511634
rect -9036 511366 592960 511398
rect -9036 507454 592960 507486
rect -9036 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 592960 507454
rect -9036 507134 592960 507218
rect -9036 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 592960 507134
rect -9036 506866 592960 506898
rect -9036 502954 592960 502986
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect -9036 502634 592960 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect -9036 502366 592960 502398
rect -9036 498454 592960 498486
rect -9036 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592960 498454
rect -9036 498134 592960 498218
rect -9036 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592960 498134
rect -9036 497866 592960 497898
rect -9036 493954 592960 493986
rect -9036 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 592960 493954
rect -9036 493634 592960 493718
rect -9036 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 592960 493634
rect -9036 493366 592960 493398
rect -9036 489454 592960 489486
rect -9036 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 592960 489454
rect -9036 489134 592960 489218
rect -9036 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 592960 489134
rect -9036 488866 592960 488898
rect -9036 484954 592960 484986
rect -9036 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 592960 484954
rect -9036 484634 592960 484718
rect -9036 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 592960 484634
rect -9036 484366 592960 484398
rect -9036 480454 592960 480486
rect -9036 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 592960 480454
rect -9036 480134 592960 480218
rect -9036 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 592960 480134
rect -9036 479866 592960 479898
rect -9036 475954 592960 475986
rect -9036 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 592960 475954
rect -9036 475634 592960 475718
rect -9036 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 592960 475634
rect -9036 475366 592960 475398
rect -9036 471454 592960 471486
rect -9036 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 592960 471454
rect -9036 471134 592960 471218
rect -9036 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 592960 471134
rect -9036 470866 592960 470898
rect -9036 466954 592960 466986
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect -9036 466634 592960 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect -9036 466366 592960 466398
rect -9036 462454 592960 462486
rect -9036 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592960 462454
rect -9036 462134 592960 462218
rect -9036 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592960 462134
rect -9036 461866 592960 461898
rect -9036 457954 592960 457986
rect -9036 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 592960 457954
rect -9036 457634 592960 457718
rect -9036 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 592960 457634
rect -9036 457366 592960 457398
rect -9036 453454 592960 453486
rect -9036 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 592960 453454
rect -9036 453134 592960 453218
rect -9036 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 592960 453134
rect -9036 452866 592960 452898
rect -9036 448954 592960 448986
rect -9036 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 592960 448954
rect -9036 448634 592960 448718
rect -9036 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 592960 448634
rect -9036 448366 592960 448398
rect -9036 444454 592960 444486
rect -9036 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 592960 444454
rect -9036 444134 592960 444218
rect -9036 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 592960 444134
rect -9036 443866 592960 443898
rect -9036 439954 592960 439986
rect -9036 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 252010 439954
rect 252246 439718 282730 439954
rect 282966 439718 313450 439954
rect 313686 439718 344170 439954
rect 344406 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 592960 439954
rect -9036 439634 592960 439718
rect -9036 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 252010 439634
rect 252246 439398 282730 439634
rect 282966 439398 313450 439634
rect 313686 439398 344170 439634
rect 344406 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 592960 439634
rect -9036 439366 592960 439398
rect -9036 435454 592960 435486
rect -9036 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 236650 435454
rect 236886 435218 267370 435454
rect 267606 435218 298090 435454
rect 298326 435218 328810 435454
rect 329046 435218 359530 435454
rect 359766 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 592960 435454
rect -9036 435134 592960 435218
rect -9036 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 236650 435134
rect 236886 434898 267370 435134
rect 267606 434898 298090 435134
rect 298326 434898 328810 435134
rect 329046 434898 359530 435134
rect 359766 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 592960 435134
rect -9036 434866 592960 434898
rect -9036 430954 592960 430986
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect -9036 430634 592960 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect -9036 430366 592960 430398
rect -9036 426454 592960 426486
rect -9036 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592960 426454
rect -9036 426134 592960 426218
rect -9036 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592960 426134
rect -9036 425866 592960 425898
rect -9036 421954 592960 421986
rect -9036 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 592960 421954
rect -9036 421634 592960 421718
rect -9036 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 592960 421634
rect -9036 421366 592960 421398
rect -9036 417454 592960 417486
rect -9036 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 592960 417454
rect -9036 417134 592960 417218
rect -9036 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 592960 417134
rect -9036 416866 592960 416898
rect -9036 412954 592960 412986
rect -9036 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 592960 412954
rect -9036 412634 592960 412718
rect -9036 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 592960 412634
rect -9036 412366 592960 412398
rect -9036 408454 592960 408486
rect -9036 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 592960 408454
rect -9036 408134 592960 408218
rect -9036 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 592960 408134
rect -9036 407866 592960 407898
rect -9036 403954 592960 403986
rect -9036 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 252010 403954
rect 252246 403718 282730 403954
rect 282966 403718 313450 403954
rect 313686 403718 344170 403954
rect 344406 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 592960 403954
rect -9036 403634 592960 403718
rect -9036 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 252010 403634
rect 252246 403398 282730 403634
rect 282966 403398 313450 403634
rect 313686 403398 344170 403634
rect 344406 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 592960 403634
rect -9036 403366 592960 403398
rect -9036 399454 592960 399486
rect -9036 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 236650 399454
rect 236886 399218 267370 399454
rect 267606 399218 298090 399454
rect 298326 399218 328810 399454
rect 329046 399218 359530 399454
rect 359766 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 592960 399454
rect -9036 399134 592960 399218
rect -9036 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 236650 399134
rect 236886 398898 267370 399134
rect 267606 398898 298090 399134
rect 298326 398898 328810 399134
rect 329046 398898 359530 399134
rect 359766 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 592960 399134
rect -9036 398866 592960 398898
rect -9036 394954 592960 394986
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect -9036 394634 592960 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect -9036 394366 592960 394398
rect -9036 390454 592960 390486
rect -9036 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592960 390454
rect -9036 390134 592960 390218
rect -9036 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592960 390134
rect -9036 389866 592960 389898
rect -9036 385954 592960 385986
rect -9036 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 592960 385954
rect -9036 385634 592960 385718
rect -9036 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 592960 385634
rect -9036 385366 592960 385398
rect -9036 381454 592960 381486
rect -9036 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 592960 381454
rect -9036 381134 592960 381218
rect -9036 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 592960 381134
rect -9036 380866 592960 380898
rect -9036 376954 592960 376986
rect -9036 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 592960 376954
rect -9036 376634 592960 376718
rect -9036 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 592960 376634
rect -9036 376366 592960 376398
rect -9036 372454 592960 372486
rect -9036 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 592960 372454
rect -9036 372134 592960 372218
rect -9036 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 592960 372134
rect -9036 371866 592960 371898
rect -9036 367954 592960 367986
rect -9036 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 252010 367954
rect 252246 367718 282730 367954
rect 282966 367718 313450 367954
rect 313686 367718 344170 367954
rect 344406 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 592960 367954
rect -9036 367634 592960 367718
rect -9036 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 252010 367634
rect 252246 367398 282730 367634
rect 282966 367398 313450 367634
rect 313686 367398 344170 367634
rect 344406 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 592960 367634
rect -9036 367366 592960 367398
rect -9036 363454 592960 363486
rect -9036 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 236650 363454
rect 236886 363218 267370 363454
rect 267606 363218 298090 363454
rect 298326 363218 328810 363454
rect 329046 363218 359530 363454
rect 359766 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 592960 363454
rect -9036 363134 592960 363218
rect -9036 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 236650 363134
rect 236886 362898 267370 363134
rect 267606 362898 298090 363134
rect 298326 362898 328810 363134
rect 329046 362898 359530 363134
rect 359766 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 592960 363134
rect -9036 362866 592960 362898
rect -9036 358954 592960 358986
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect -9036 358634 592960 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect -9036 358366 592960 358398
rect -9036 354454 592960 354486
rect -9036 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592960 354454
rect -9036 354134 592960 354218
rect -9036 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592960 354134
rect -9036 353866 592960 353898
rect -9036 349954 592960 349986
rect -9036 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 592960 349954
rect -9036 349634 592960 349718
rect -9036 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 592960 349634
rect -9036 349366 592960 349398
rect -9036 345454 592960 345486
rect -9036 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 592960 345454
rect -9036 345134 592960 345218
rect -9036 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 592960 345134
rect -9036 344866 592960 344898
rect -9036 340954 592960 340986
rect -9036 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 592960 340954
rect -9036 340634 592960 340718
rect -9036 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 592960 340634
rect -9036 340366 592960 340398
rect -9036 336454 592960 336486
rect -9036 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 592960 336454
rect -9036 336134 592960 336218
rect -9036 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 592960 336134
rect -9036 335866 592960 335898
rect -9036 331954 592960 331986
rect -9036 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 252010 331954
rect 252246 331718 282730 331954
rect 282966 331718 313450 331954
rect 313686 331718 344170 331954
rect 344406 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 592960 331954
rect -9036 331634 592960 331718
rect -9036 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 252010 331634
rect 252246 331398 282730 331634
rect 282966 331398 313450 331634
rect 313686 331398 344170 331634
rect 344406 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 592960 331634
rect -9036 331366 592960 331398
rect -9036 327454 592960 327486
rect -9036 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 236650 327454
rect 236886 327218 267370 327454
rect 267606 327218 298090 327454
rect 298326 327218 328810 327454
rect 329046 327218 359530 327454
rect 359766 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 592960 327454
rect -9036 327134 592960 327218
rect -9036 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 236650 327134
rect 236886 326898 267370 327134
rect 267606 326898 298090 327134
rect 298326 326898 328810 327134
rect 329046 326898 359530 327134
rect 359766 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 592960 327134
rect -9036 326866 592960 326898
rect -9036 322954 592960 322986
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect -9036 322634 592960 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect -9036 322366 592960 322398
rect -9036 318454 592960 318486
rect -9036 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592960 318454
rect -9036 318134 592960 318218
rect -9036 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592960 318134
rect -9036 317866 592960 317898
rect -9036 313954 592960 313986
rect -9036 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 592960 313954
rect -9036 313634 592960 313718
rect -9036 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 592960 313634
rect -9036 313366 592960 313398
rect -9036 309454 592960 309486
rect -9036 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 592960 309454
rect -9036 309134 592960 309218
rect -9036 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 592960 309134
rect -9036 308866 592960 308898
rect -9036 304954 592960 304986
rect -9036 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 592960 304954
rect -9036 304634 592960 304718
rect -9036 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 592960 304634
rect -9036 304366 592960 304398
rect -9036 300454 592960 300486
rect -9036 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 592960 300454
rect -9036 300134 592960 300218
rect -9036 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 592960 300134
rect -9036 299866 592960 299898
rect -9036 295954 592960 295986
rect -9036 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 592960 295954
rect -9036 295634 592960 295718
rect -9036 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 592960 295634
rect -9036 295366 592960 295398
rect -9036 291454 592960 291486
rect -9036 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 592960 291454
rect -9036 291134 592960 291218
rect -9036 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 592960 291134
rect -9036 290866 592960 290898
rect -9036 286954 592960 286986
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect -9036 286634 592960 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect -9036 286366 592960 286398
rect -9036 282454 592960 282486
rect -9036 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592960 282454
rect -9036 282134 592960 282218
rect -9036 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592960 282134
rect -9036 281866 592960 281898
rect -9036 277954 592960 277986
rect -9036 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 592960 277954
rect -9036 277634 592960 277718
rect -9036 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 592960 277634
rect -9036 277366 592960 277398
rect -9036 273454 592960 273486
rect -9036 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 592960 273454
rect -9036 273134 592960 273218
rect -9036 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 592960 273134
rect -9036 272866 592960 272898
rect -9036 268954 592960 268986
rect -9036 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 592960 268954
rect -9036 268634 592960 268718
rect -9036 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 592960 268634
rect -9036 268366 592960 268398
rect -9036 264454 592960 264486
rect -9036 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 592960 264454
rect -9036 264134 592960 264218
rect -9036 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 592960 264134
rect -9036 263866 592960 263898
rect -9036 259954 592960 259986
rect -9036 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 592960 259954
rect -9036 259634 592960 259718
rect -9036 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 592960 259634
rect -9036 259366 592960 259398
rect -9036 255454 592960 255486
rect -9036 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 592960 255454
rect -9036 255134 592960 255218
rect -9036 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 592960 255134
rect -9036 254866 592960 254898
rect -9036 250954 592960 250986
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect -9036 250634 592960 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect -9036 250366 592960 250398
rect -9036 246454 592960 246486
rect -9036 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592960 246454
rect -9036 246134 592960 246218
rect -9036 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592960 246134
rect -9036 245866 592960 245898
rect -9036 241954 592960 241986
rect -9036 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 592960 241954
rect -9036 241634 592960 241718
rect -9036 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 592960 241634
rect -9036 241366 592960 241398
rect -9036 237454 592960 237486
rect -9036 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 592960 237454
rect -9036 237134 592960 237218
rect -9036 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 592960 237134
rect -9036 236866 592960 236898
rect -9036 232954 592960 232986
rect -9036 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 592960 232954
rect -9036 232634 592960 232718
rect -9036 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 592960 232634
rect -9036 232366 592960 232398
rect -9036 228454 592960 228486
rect -9036 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 592960 228454
rect -9036 228134 592960 228218
rect -9036 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 592960 228134
rect -9036 227866 592960 227898
rect -9036 223954 592960 223986
rect -9036 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 220328 223954
rect 220564 223718 356056 223954
rect 356292 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 592960 223954
rect -9036 223634 592960 223718
rect -9036 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 220328 223634
rect 220564 223398 356056 223634
rect 356292 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 592960 223634
rect -9036 223366 592960 223398
rect -9036 219454 592960 219486
rect -9036 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 592960 219454
rect -9036 219134 592960 219218
rect -9036 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 592960 219134
rect -9036 218866 592960 218898
rect -9036 214954 592960 214986
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect -9036 214634 592960 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect -9036 214366 592960 214398
rect -9036 210454 592960 210486
rect -9036 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592960 210454
rect -9036 210134 592960 210218
rect -9036 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592960 210134
rect -9036 209866 592960 209898
rect -9036 205954 592960 205986
rect -9036 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 592960 205954
rect -9036 205634 592960 205718
rect -9036 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 592960 205634
rect -9036 205366 592960 205398
rect -9036 201454 592960 201486
rect -9036 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 592960 201454
rect -9036 201134 592960 201218
rect -9036 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 592960 201134
rect -9036 200866 592960 200898
rect -9036 196954 592960 196986
rect -9036 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 592960 196954
rect -9036 196634 592960 196718
rect -9036 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 592960 196634
rect -9036 196366 592960 196398
rect -9036 192454 592960 192486
rect -9036 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 592960 192454
rect -9036 192134 592960 192218
rect -9036 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 592960 192134
rect -9036 191866 592960 191898
rect -9036 187954 592960 187986
rect -9036 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 220328 187954
rect 220564 187718 356056 187954
rect 356292 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 592960 187954
rect -9036 187634 592960 187718
rect -9036 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 220328 187634
rect 220564 187398 356056 187634
rect 356292 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 592960 187634
rect -9036 187366 592960 187398
rect -9036 183454 592960 183486
rect -9036 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 592960 183454
rect -9036 183134 592960 183218
rect -9036 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 592960 183134
rect -9036 182866 592960 182898
rect -9036 178954 592960 178986
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect -9036 178634 592960 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect -9036 178366 592960 178398
rect -9036 174454 592960 174486
rect -9036 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592960 174454
rect -9036 174134 592960 174218
rect -9036 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592960 174134
rect -9036 173866 592960 173898
rect -9036 169954 592960 169986
rect -9036 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 592960 169954
rect -9036 169634 592960 169718
rect -9036 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 592960 169634
rect -9036 169366 592960 169398
rect -9036 165454 592960 165486
rect -9036 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 592960 165454
rect -9036 165134 592960 165218
rect -9036 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 592960 165134
rect -9036 164866 592960 164898
rect -9036 160954 592960 160986
rect -9036 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 592960 160954
rect -9036 160634 592960 160718
rect -9036 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 592960 160634
rect -9036 160366 592960 160398
rect -9036 156454 592960 156486
rect -9036 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 592960 156454
rect -9036 156134 592960 156218
rect -9036 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 592960 156134
rect -9036 155866 592960 155898
rect -9036 151954 592960 151986
rect -9036 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 592960 151954
rect -9036 151634 592960 151718
rect -9036 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 592960 151634
rect -9036 151366 592960 151398
rect -9036 147454 592960 147486
rect -9036 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 592960 147454
rect -9036 147134 592960 147218
rect -9036 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 592960 147134
rect -9036 146866 592960 146898
rect -9036 142954 592960 142986
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect -9036 142634 592960 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect -9036 142366 592960 142398
rect -9036 138454 592960 138486
rect -9036 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592960 138454
rect -9036 138134 592960 138218
rect -9036 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592960 138134
rect -9036 137866 592960 137898
rect -9036 133954 592960 133986
rect -9036 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 592960 133954
rect -9036 133634 592960 133718
rect -9036 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 592960 133634
rect -9036 133366 592960 133398
rect -9036 129454 592960 129486
rect -9036 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 592960 129454
rect -9036 129134 592960 129218
rect -9036 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 592960 129134
rect -9036 128866 592960 128898
rect -9036 124954 592960 124986
rect -9036 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 592960 124954
rect -9036 124634 592960 124718
rect -9036 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 592960 124634
rect -9036 124366 592960 124398
rect -9036 120454 592960 120486
rect -9036 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 592960 120454
rect -9036 120134 592960 120218
rect -9036 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 592960 120134
rect -9036 119866 592960 119898
rect -9036 115954 592960 115986
rect -9036 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 592960 115954
rect -9036 115634 592960 115718
rect -9036 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 592960 115634
rect -9036 115366 592960 115398
rect -9036 111454 592960 111486
rect -9036 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 592960 111454
rect -9036 111134 592960 111218
rect -9036 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 592960 111134
rect -9036 110866 592960 110898
rect -9036 106954 592960 106986
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect -9036 106634 592960 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect -9036 106366 592960 106398
rect -9036 102454 592960 102486
rect -9036 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592960 102454
rect -9036 102134 592960 102218
rect -9036 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592960 102134
rect -9036 101866 592960 101898
rect -9036 97954 592960 97986
rect -9036 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 592960 97954
rect -9036 97634 592960 97718
rect -9036 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 592960 97634
rect -9036 97366 592960 97398
rect -9036 93454 592960 93486
rect -9036 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 592960 93454
rect -9036 93134 592960 93218
rect -9036 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 592960 93134
rect -9036 92866 592960 92898
rect -9036 88954 592960 88986
rect -9036 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 592960 88954
rect -9036 88634 592960 88718
rect -9036 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 592960 88634
rect -9036 88366 592960 88398
rect -9036 84454 592960 84486
rect -9036 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 592960 84454
rect -9036 84134 592960 84218
rect -9036 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 592960 84134
rect -9036 83866 592960 83898
rect -9036 79954 592960 79986
rect -9036 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 592960 79954
rect -9036 79634 592960 79718
rect -9036 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 592960 79634
rect -9036 79366 592960 79398
rect -9036 75454 592960 75486
rect -9036 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 592960 75454
rect -9036 75134 592960 75218
rect -9036 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 592960 75134
rect -9036 74866 592960 74898
rect -9036 70954 592960 70986
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect -9036 70634 592960 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect -9036 70366 592960 70398
rect -9036 66454 592960 66486
rect -9036 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592960 66454
rect -9036 66134 592960 66218
rect -9036 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592960 66134
rect -9036 65866 592960 65898
rect -9036 61954 592960 61986
rect -9036 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 592960 61954
rect -9036 61634 592960 61718
rect -9036 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 592960 61634
rect -9036 61366 592960 61398
rect -9036 57454 592960 57486
rect -9036 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 592960 57454
rect -9036 57134 592960 57218
rect -9036 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 592960 57134
rect -9036 56866 592960 56898
rect -9036 52954 592960 52986
rect -9036 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 592960 52954
rect -9036 52634 592960 52718
rect -9036 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 592960 52634
rect -9036 52366 592960 52398
rect -9036 48454 592960 48486
rect -9036 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 592960 48454
rect -9036 48134 592960 48218
rect -9036 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 592960 48134
rect -9036 47866 592960 47898
rect -9036 43954 592960 43986
rect -9036 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 592960 43954
rect -9036 43634 592960 43718
rect -9036 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 592960 43634
rect -9036 43366 592960 43398
rect -9036 39454 592960 39486
rect -9036 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 592960 39454
rect -9036 39134 592960 39218
rect -9036 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 592960 39134
rect -9036 38866 592960 38898
rect -9036 34954 592960 34986
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect -9036 34634 592960 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect -9036 34366 592960 34398
rect -9036 30454 592960 30486
rect -9036 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592960 30454
rect -9036 30134 592960 30218
rect -9036 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592960 30134
rect -9036 29866 592960 29898
rect -9036 25954 592960 25986
rect -9036 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 592960 25954
rect -9036 25634 592960 25718
rect -9036 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 592960 25634
rect -9036 25366 592960 25398
rect -9036 21454 592960 21486
rect -9036 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 592960 21454
rect -9036 21134 592960 21218
rect -9036 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 592960 21134
rect -9036 20866 592960 20898
rect -9036 16954 592960 16986
rect -9036 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 592960 16954
rect -9036 16634 592960 16718
rect -9036 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 592960 16634
rect -9036 16366 592960 16398
rect -9036 12454 592960 12486
rect -9036 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 592960 12454
rect -9036 12134 592960 12218
rect -9036 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 592960 12134
rect -9036 11866 592960 11898
rect -9036 7954 592960 7986
rect -9036 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 592960 7954
rect -9036 7634 592960 7718
rect -9036 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 592960 7634
rect -9036 7366 592960 7398
rect -9036 3454 592960 3486
rect -9036 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 592960 3454
rect -9036 3134 592960 3218
rect -9036 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 592960 3134
rect -9036 2866 592960 2898
rect -2316 -656 586240 -624
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect -2316 -976 586240 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect -2316 -1244 586240 -1212
rect -3276 -1616 587200 -1584
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect -3276 -1936 587200 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect -3276 -2204 587200 -2172
rect -4236 -2576 588160 -2544
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect -4236 -2896 588160 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect -4236 -3164 588160 -3132
rect -5196 -3536 589120 -3504
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect -5196 -3856 589120 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect -5196 -4124 589120 -4092
rect -6156 -4496 590080 -4464
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect -6156 -4816 590080 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect -6156 -5084 590080 -5052
rect -7116 -5456 591040 -5424
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect -7116 -5776 591040 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect -7116 -6044 591040 -6012
rect -8076 -6416 592000 -6384
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect -8076 -6736 592000 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect -8076 -7004 592000 -6972
rect -9036 -7376 592960 -7344
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect -9036 -7696 592960 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect -9036 -7964 592960 -7932
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst
timestamp 0
transform 1 0 220000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 232400 0 1 310400
box 14 0 130166 132435
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2316 -1244 -1696 705180 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 -1244 586240 -624 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 704560 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585620 -1244 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7964 2414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7964 38414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7964 74414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7964 110414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7964 146414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7964 182414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7964 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7964 254414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 245308 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7964 290414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 245308 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7964 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7964 362414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 444835 362414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7964 398414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7964 434414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7964 470414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7964 506414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7964 542414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7964 578414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 2866 592960 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 38866 592960 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 74866 592960 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 110866 592960 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 146866 592960 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 182866 592960 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 218866 592960 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 254866 592960 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 290866 592960 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 326866 592960 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 362866 592960 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 398866 592960 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 434866 592960 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 470866 592960 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 506866 592960 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 542866 592960 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 578866 592960 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 614866 592960 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 650866 592960 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 686866 592960 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -4236 -3164 -3616 707100 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 -3164 588160 -2544 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 706480 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587540 -3164 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7964 11414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7964 47414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7964 83414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7964 119414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7964 155414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7964 191414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7964 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7964 263414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 245308 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7964 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7964 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7964 371414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7964 407414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7964 443414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7964 479414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7964 515414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7964 551414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 11866 592960 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 47866 592960 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 83866 592960 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 119866 592960 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 155866 592960 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 191866 592960 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 227866 592960 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 263866 592960 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 299866 592960 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 335866 592960 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 371866 592960 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 407866 592960 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 443866 592960 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 479866 592960 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 515866 592960 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 551866 592960 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 587866 592960 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 623866 592960 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 659866 592960 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 695866 592960 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5196 -4124 -4576 708060 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 -4124 589120 -3504 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 707440 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 588500 -4124 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 15294 -7964 15914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 51294 -7964 51914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 87294 -7964 87914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 -7964 123914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 -7964 159914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 195294 -7964 195914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 -7964 231914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 565308 231914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 -7964 267914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 245308 267914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 565308 267914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 -7964 303914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 565308 303914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 -7964 339914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 565308 339914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 375294 -7964 375914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 411294 -7964 411914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 447294 -7964 447914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 483294 -7964 483914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 519294 -7964 519914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 555294 -7964 555914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 16366 592960 16986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 52366 592960 52986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 88366 592960 88986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 124366 592960 124986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 160366 592960 160986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 196366 592960 196986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 232366 592960 232986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 268366 592960 268986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 304366 592960 304986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 340366 592960 340986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 376366 592960 376986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 412366 592960 412986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 448366 592960 448986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 484366 592960 484986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 520366 592960 520986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 556366 592960 556986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 592366 592960 592986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 628366 592960 628986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 664366 592960 664986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 700366 592960 700986 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -6156 -5084 -5536 709020 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 -5084 590080 -4464 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 708400 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 589460 -5084 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 19794 -7964 20414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 55794 -7964 56414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 91794 -7964 92414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 -7964 128414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 -7964 164414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 199794 -7964 200414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 -7964 236414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 -7964 272414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 -7964 308414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 -7964 344414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 379794 -7964 380414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 415794 -7964 416414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 451794 -7964 452414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 487794 -7964 488414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 523794 -7964 524414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 559794 -7964 560414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 20866 592960 21486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 56866 592960 57486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 92866 592960 93486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 128866 592960 129486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 164866 592960 165486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 200866 592960 201486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 236866 592960 237486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 272866 592960 273486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 308866 592960 309486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 344866 592960 345486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 380866 592960 381486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 416866 592960 417486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 452866 592960 453486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 488866 592960 489486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 524866 592960 525486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 560866 592960 561486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 596866 592960 597486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 632866 592960 633486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 668866 592960 669486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -8076 -7004 -7456 710940 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 -7004 592000 -6384 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 710320 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 591380 -7004 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 28794 -7964 29414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 64794 -7964 65414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 -7964 101414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 -7964 137414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 172794 -7964 173414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 208794 -7964 209414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 -7964 245414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 245308 245414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 565308 245414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 -7964 281414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 245308 281414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 565308 281414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 -7964 317414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 565308 317414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 -7964 353414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 565308 353414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 388794 -7964 389414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 424794 -7964 425414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 460794 -7964 461414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 496794 -7964 497414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 532794 -7964 533414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 568794 -7964 569414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 29866 592960 30486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 65866 592960 66486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 101866 592960 102486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 137866 592960 138486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 173866 592960 174486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 209866 592960 210486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 245866 592960 246486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 281866 592960 282486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 317866 592960 318486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 353866 592960 354486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 389866 592960 390486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 425866 592960 426486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 461866 592960 462486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 497866 592960 498486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 533866 592960 534486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 569866 592960 570486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 605866 592960 606486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 641866 592960 642486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 677866 592960 678486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -9036 -7964 -8416 711900 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 -7964 592960 -7344 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 711280 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592340 -7964 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7964 33914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7964 69914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7964 105914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7964 141914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7964 177914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7964 213914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7964 249914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 245308 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7964 285914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 245308 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7964 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7964 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7964 393914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7964 429914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7964 465914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7964 501914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7964 537914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7964 573914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 34366 592960 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 70366 592960 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 106366 592960 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 142366 592960 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 178366 592960 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 214366 592960 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 250366 592960 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 286366 592960 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 322366 592960 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 358366 592960 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 394366 592960 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 430366 592960 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 466366 592960 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 502366 592960 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 538366 592960 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 574366 592960 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 610366 592960 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 646366 592960 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 682366 592960 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -3276 -2204 -2656 706140 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 -2204 587200 -1584 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 705520 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586580 -2204 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7964 6914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7964 42914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7964 78914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7964 114914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7964 150914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7964 186914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7964 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7964 258914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 245308 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7964 294914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 245308 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7964 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7964 366914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7964 402914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7964 438914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7964 474914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7964 510914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7964 546914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7964 582914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 7366 592960 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 43366 592960 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 79366 592960 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 115366 592960 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 151366 592960 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 187366 592960 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 223366 592960 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 259366 592960 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 295366 592960 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 331366 592960 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 367366 592960 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 403366 592960 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 439366 592960 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 475366 592960 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 511366 592960 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 547366 592960 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 583366 592960 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 619366 592960 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 655366 592960 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 691366 592960 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -7116 -6044 -6496 709980 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 -6044 591040 -5424 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 709360 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 590420 -6044 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 24294 -7964 24914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 60294 -7964 60914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 96294 -7964 96914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 -7964 132914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 -7964 168914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 204294 -7964 204914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 -7964 240914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 -7964 276914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 -7964 312914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 -7964 348914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 384294 -7964 384914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 420294 -7964 420914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 456294 -7964 456914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 492294 -7964 492914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 528294 -7964 528914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 564294 -7964 564914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 25366 592960 25986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 61366 592960 61986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 97366 592960 97986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 133366 592960 133986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 169366 592960 169986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 205366 592960 205986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 241366 592960 241986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 277366 592960 277986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 313366 592960 313986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 349366 592960 349986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 385366 592960 385986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 421366 592960 421986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 457366 592960 457986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 493366 592960 493986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 529366 592960 529986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 565366 592960 565986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 601366 592960 601986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 637366 592960 637986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 673366 592960 673986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
