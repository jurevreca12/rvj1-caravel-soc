magic
tech sky130A
magscale 1 2
timestamp 1653482387
<< obsli1 >>
rect 1104 2159 68908 69649
<< obsm1 >>
rect 14 1980 69630 69680
<< metal2 >>
rect 662 71364 718 72164
rect 3238 71364 3294 72164
rect 5814 71364 5870 72164
rect 8390 71364 8446 72164
rect 10966 71364 11022 72164
rect 13542 71364 13598 72164
rect 16118 71364 16174 72164
rect 18694 71364 18750 72164
rect 21270 71364 21326 72164
rect 23846 71364 23902 72164
rect 26422 71364 26478 72164
rect 28998 71364 29054 72164
rect 31574 71364 31630 72164
rect 34150 71364 34206 72164
rect 36726 71364 36782 72164
rect 39302 71364 39358 72164
rect 41878 71364 41934 72164
rect 44454 71364 44510 72164
rect 47030 71364 47086 72164
rect 49606 71364 49662 72164
rect 52182 71364 52238 72164
rect 54758 71364 54814 72164
rect 57334 71364 57390 72164
rect 59910 71364 59966 72164
rect 62486 71364 62542 72164
rect 65062 71364 65118 72164
rect 67638 71364 67694 72164
rect 69570 71364 69626 72164
rect 18 0 74 800
rect 1950 0 2006 800
rect 4526 0 4582 800
rect 7102 0 7158 800
rect 9678 0 9734 800
rect 12254 0 12310 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 22558 0 22614 800
rect 25134 0 25190 800
rect 27710 0 27766 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 38014 0 38070 800
rect 40590 0 40646 800
rect 43166 0 43222 800
rect 45742 0 45798 800
rect 48318 0 48374 800
rect 50894 0 50950 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 58622 0 58678 800
rect 61198 0 61254 800
rect 63774 0 63830 800
rect 66350 0 66406 800
rect 68926 0 68982 800
<< obsm2 >>
rect 20 71308 606 71482
rect 774 71308 3182 71482
rect 3350 71308 5758 71482
rect 5926 71308 8334 71482
rect 8502 71308 10910 71482
rect 11078 71308 13486 71482
rect 13654 71308 16062 71482
rect 16230 71308 18638 71482
rect 18806 71308 21214 71482
rect 21382 71308 23790 71482
rect 23958 71308 26366 71482
rect 26534 71308 28942 71482
rect 29110 71308 31518 71482
rect 31686 71308 34094 71482
rect 34262 71308 36670 71482
rect 36838 71308 39246 71482
rect 39414 71308 41822 71482
rect 41990 71308 44398 71482
rect 44566 71308 46974 71482
rect 47142 71308 49550 71482
rect 49718 71308 52126 71482
rect 52294 71308 54702 71482
rect 54870 71308 57278 71482
rect 57446 71308 59854 71482
rect 60022 71308 62430 71482
rect 62598 71308 65006 71482
rect 65174 71308 67582 71482
rect 67750 71308 69514 71482
rect 20 856 69624 71308
rect 130 734 1894 856
rect 2062 734 4470 856
rect 4638 734 7046 856
rect 7214 734 9622 856
rect 9790 734 12198 856
rect 12366 734 14774 856
rect 14942 734 17350 856
rect 17518 734 19926 856
rect 20094 734 22502 856
rect 22670 734 25078 856
rect 25246 734 27654 856
rect 27822 734 30230 856
rect 30398 734 32806 856
rect 32974 734 35382 856
rect 35550 734 37958 856
rect 38126 734 40534 856
rect 40702 734 43110 856
rect 43278 734 45686 856
rect 45854 734 48262 856
rect 48430 734 50838 856
rect 51006 734 53414 856
rect 53582 734 55990 856
rect 56158 734 58566 856
rect 58734 734 61142 856
rect 61310 734 63718 856
rect 63886 734 66294 856
rect 66462 734 68870 856
rect 69038 734 69624 856
<< metal3 >>
rect 0 70048 800 70168
rect 69220 69368 70020 69488
rect 0 67328 800 67448
rect 69220 66648 70020 66768
rect 0 64608 800 64728
rect 69220 63928 70020 64048
rect 0 61888 800 62008
rect 69220 61208 70020 61328
rect 0 59168 800 59288
rect 69220 58488 70020 58608
rect 0 56448 800 56568
rect 69220 55768 70020 55888
rect 0 53728 800 53848
rect 69220 53048 70020 53168
rect 0 51008 800 51128
rect 69220 50328 70020 50448
rect 0 48288 800 48408
rect 69220 47608 70020 47728
rect 0 45568 800 45688
rect 69220 44888 70020 45008
rect 0 42848 800 42968
rect 69220 42168 70020 42288
rect 0 40128 800 40248
rect 69220 39448 70020 39568
rect 0 37408 800 37528
rect 69220 36728 70020 36848
rect 0 34688 800 34808
rect 69220 34008 70020 34128
rect 0 31968 800 32088
rect 69220 31288 70020 31408
rect 0 29248 800 29368
rect 69220 28568 70020 28688
rect 0 26528 800 26648
rect 69220 25848 70020 25968
rect 0 23808 800 23928
rect 69220 23128 70020 23248
rect 0 21088 800 21208
rect 69220 20408 70020 20528
rect 0 18368 800 18488
rect 69220 17688 70020 17808
rect 0 15648 800 15768
rect 69220 14968 70020 15088
rect 0 12928 800 13048
rect 69220 12248 70020 12368
rect 0 10208 800 10328
rect 69220 9528 70020 9648
rect 0 7488 800 7608
rect 69220 6808 70020 6928
rect 0 4768 800 4888
rect 69220 4088 70020 4208
rect 0 2048 800 2168
rect 69220 1368 70020 1488
<< obsm3 >>
rect 880 69968 69220 70141
rect 800 69568 69220 69968
rect 800 69288 69140 69568
rect 800 67528 69220 69288
rect 880 67248 69220 67528
rect 800 66848 69220 67248
rect 800 66568 69140 66848
rect 800 64808 69220 66568
rect 880 64528 69220 64808
rect 800 64128 69220 64528
rect 800 63848 69140 64128
rect 800 62088 69220 63848
rect 880 61808 69220 62088
rect 800 61408 69220 61808
rect 800 61128 69140 61408
rect 800 59368 69220 61128
rect 880 59088 69220 59368
rect 800 58688 69220 59088
rect 800 58408 69140 58688
rect 800 56648 69220 58408
rect 880 56368 69220 56648
rect 800 55968 69220 56368
rect 800 55688 69140 55968
rect 800 53928 69220 55688
rect 880 53648 69220 53928
rect 800 53248 69220 53648
rect 800 52968 69140 53248
rect 800 51208 69220 52968
rect 880 50928 69220 51208
rect 800 50528 69220 50928
rect 800 50248 69140 50528
rect 800 48488 69220 50248
rect 880 48208 69220 48488
rect 800 47808 69220 48208
rect 800 47528 69140 47808
rect 800 45768 69220 47528
rect 880 45488 69220 45768
rect 800 45088 69220 45488
rect 800 44808 69140 45088
rect 800 43048 69220 44808
rect 880 42768 69220 43048
rect 800 42368 69220 42768
rect 800 42088 69140 42368
rect 800 40328 69220 42088
rect 880 40048 69220 40328
rect 800 39648 69220 40048
rect 800 39368 69140 39648
rect 800 37608 69220 39368
rect 880 37328 69220 37608
rect 800 36928 69220 37328
rect 800 36648 69140 36928
rect 800 34888 69220 36648
rect 880 34608 69220 34888
rect 800 34208 69220 34608
rect 800 33928 69140 34208
rect 800 32168 69220 33928
rect 880 31888 69220 32168
rect 800 31488 69220 31888
rect 800 31208 69140 31488
rect 800 29448 69220 31208
rect 880 29168 69220 29448
rect 800 28768 69220 29168
rect 800 28488 69140 28768
rect 800 26728 69220 28488
rect 880 26448 69220 26728
rect 800 26048 69220 26448
rect 800 25768 69140 26048
rect 800 24008 69220 25768
rect 880 23728 69220 24008
rect 800 23328 69220 23728
rect 800 23048 69140 23328
rect 800 21288 69220 23048
rect 880 21008 69220 21288
rect 800 20608 69220 21008
rect 800 20328 69140 20608
rect 800 18568 69220 20328
rect 880 18288 69220 18568
rect 800 17888 69220 18288
rect 800 17608 69140 17888
rect 800 15848 69220 17608
rect 880 15568 69220 15848
rect 800 15168 69220 15568
rect 800 14888 69140 15168
rect 800 13128 69220 14888
rect 880 12848 69220 13128
rect 800 12448 69220 12848
rect 800 12168 69140 12448
rect 800 10408 69220 12168
rect 880 10128 69220 10408
rect 800 9728 69220 10128
rect 800 9448 69140 9728
rect 800 7688 69220 9448
rect 880 7408 69220 7688
rect 800 7008 69220 7408
rect 800 6728 69140 7008
rect 800 4968 69220 6728
rect 880 4688 69220 4968
rect 800 4288 69220 4688
rect 800 4008 69140 4288
rect 800 2248 69220 4008
rect 880 1968 69220 2248
rect 800 1568 69220 1968
rect 800 1395 69140 1568
<< metal4 >>
rect 4208 2128 4528 69680
rect 19568 2128 19888 69680
rect 34928 2128 35248 69680
rect 50288 2128 50608 69680
rect 65648 2128 65968 69680
<< obsm4 >>
rect 15147 2347 19488 68781
rect 19968 2347 34848 68781
rect 35328 2347 50208 68781
rect 50688 2347 65568 68781
rect 66048 2347 66181 68781
<< labels >>
rlabel metal3 s 69220 50328 70020 50448 6 clk_i
port 1 nsew signal input
rlabel metal2 s 65062 71364 65118 72164 6 rst_i
port 2 nsew signal input
rlabel metal2 s 41878 71364 41934 72164 6 uart_rx_i
port 3 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 uart_tx_o
port 4 nsew signal output
rlabel metal4 s 4208 2128 4528 69680 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 69680 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 69680 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 69680 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 69680 6 vssd1
port 6 nsew ground bidirectional
rlabel metal2 s 39302 71364 39358 72164 6 wbs_ack_o
port 7 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 wbs_adr_i[0]
port 8 nsew signal input
rlabel metal3 s 69220 1368 70020 1488 6 wbs_adr_i[10]
port 9 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_adr_i[11]
port 10 nsew signal input
rlabel metal3 s 69220 61208 70020 61328 6 wbs_adr_i[12]
port 11 nsew signal input
rlabel metal2 s 28998 71364 29054 72164 6 wbs_adr_i[13]
port 12 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 wbs_adr_i[14]
port 13 nsew signal input
rlabel metal2 s 34150 71364 34206 72164 6 wbs_adr_i[15]
port 14 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 wbs_adr_i[16]
port 15 nsew signal input
rlabel metal3 s 69220 25848 70020 25968 6 wbs_adr_i[17]
port 16 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[18]
port 17 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 wbs_adr_i[19]
port 18 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 wbs_adr_i[1]
port 19 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_adr_i[20]
port 20 nsew signal input
rlabel metal2 s 49606 71364 49662 72164 6 wbs_adr_i[21]
port 21 nsew signal input
rlabel metal2 s 59910 71364 59966 72164 6 wbs_adr_i[22]
port 22 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[23]
port 23 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[24]
port 24 nsew signal input
rlabel metal3 s 69220 69368 70020 69488 6 wbs_adr_i[25]
port 25 nsew signal input
rlabel metal3 s 69220 17688 70020 17808 6 wbs_adr_i[26]
port 26 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wbs_adr_i[27]
port 27 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_adr_i[28]
port 28 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_adr_i[29]
port 29 nsew signal input
rlabel metal3 s 69220 14968 70020 15088 6 wbs_adr_i[2]
port 30 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wbs_adr_i[30]
port 31 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 wbs_adr_i[31]
port 32 nsew signal input
rlabel metal3 s 69220 12248 70020 12368 6 wbs_adr_i[3]
port 33 nsew signal input
rlabel metal2 s 36726 71364 36782 72164 6 wbs_adr_i[4]
port 34 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 wbs_adr_i[5]
port 35 nsew signal input
rlabel metal2 s 44454 71364 44510 72164 6 wbs_adr_i[6]
port 36 nsew signal input
rlabel metal3 s 69220 55768 70020 55888 6 wbs_adr_i[7]
port 37 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[8]
port 38 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 wbs_adr_i[9]
port 39 nsew signal input
rlabel metal3 s 69220 63928 70020 64048 6 wbs_cyc_i
port 40 nsew signal input
rlabel metal2 s 69570 71364 69626 72164 6 wbs_dat_i[0]
port 41 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 wbs_dat_i[10]
port 42 nsew signal input
rlabel metal2 s 21270 71364 21326 72164 6 wbs_dat_i[11]
port 43 nsew signal input
rlabel metal3 s 69220 31288 70020 31408 6 wbs_dat_i[12]
port 44 nsew signal input
rlabel metal2 s 23846 71364 23902 72164 6 wbs_dat_i[13]
port 45 nsew signal input
rlabel metal3 s 69220 58488 70020 58608 6 wbs_dat_i[14]
port 46 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_dat_i[15]
port 47 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[16]
port 48 nsew signal input
rlabel metal2 s 26422 71364 26478 72164 6 wbs_dat_i[17]
port 49 nsew signal input
rlabel metal3 s 69220 4088 70020 4208 6 wbs_dat_i[18]
port 50 nsew signal input
rlabel metal3 s 69220 39448 70020 39568 6 wbs_dat_i[19]
port 51 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[1]
port 52 nsew signal input
rlabel metal2 s 16118 71364 16174 72164 6 wbs_dat_i[20]
port 53 nsew signal input
rlabel metal3 s 69220 6808 70020 6928 6 wbs_dat_i[21]
port 54 nsew signal input
rlabel metal3 s 69220 66648 70020 66768 6 wbs_dat_i[22]
port 55 nsew signal input
rlabel metal2 s 57334 71364 57390 72164 6 wbs_dat_i[23]
port 56 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_i[24]
port 57 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[25]
port 58 nsew signal input
rlabel metal3 s 69220 20408 70020 20528 6 wbs_dat_i[26]
port 59 nsew signal input
rlabel metal2 s 18694 71364 18750 72164 6 wbs_dat_i[27]
port 60 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 wbs_dat_i[28]
port 61 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_dat_i[29]
port 62 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 wbs_dat_i[2]
port 63 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[30]
port 64 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 wbs_dat_i[31]
port 65 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[3]
port 66 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[4]
port 67 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wbs_dat_i[5]
port 68 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_i[6]
port 69 nsew signal input
rlabel metal3 s 69220 36728 70020 36848 6 wbs_dat_i[7]
port 70 nsew signal input
rlabel metal3 s 69220 23128 70020 23248 6 wbs_dat_i[8]
port 71 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_i[9]
port 72 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 wbs_dat_o[0]
port 73 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 wbs_dat_o[10]
port 74 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_o[11]
port 75 nsew signal output
rlabel metal3 s 69220 28568 70020 28688 6 wbs_dat_o[12]
port 76 nsew signal output
rlabel metal3 s 69220 47608 70020 47728 6 wbs_dat_o[13]
port 77 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_o[14]
port 78 nsew signal output
rlabel metal3 s 69220 53048 70020 53168 6 wbs_dat_o[15]
port 79 nsew signal output
rlabel metal2 s 5814 71364 5870 72164 6 wbs_dat_o[16]
port 80 nsew signal output
rlabel metal2 s 8390 71364 8446 72164 6 wbs_dat_o[17]
port 81 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[18]
port 82 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 83 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_o[1]
port 84 nsew signal output
rlabel metal2 s 10966 71364 11022 72164 6 wbs_dat_o[20]
port 85 nsew signal output
rlabel metal2 s 31574 71364 31630 72164 6 wbs_dat_o[21]
port 86 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 wbs_dat_o[22]
port 87 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 wbs_dat_o[23]
port 88 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[24]
port 89 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[25]
port 90 nsew signal output
rlabel metal2 s 62486 71364 62542 72164 6 wbs_dat_o[26]
port 91 nsew signal output
rlabel metal2 s 47030 71364 47086 72164 6 wbs_dat_o[27]
port 92 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[28]
port 93 nsew signal output
rlabel metal2 s 67638 71364 67694 72164 6 wbs_dat_o[29]
port 94 nsew signal output
rlabel metal3 s 69220 9528 70020 9648 6 wbs_dat_o[2]
port 95 nsew signal output
rlabel metal2 s 662 71364 718 72164 6 wbs_dat_o[30]
port 96 nsew signal output
rlabel metal3 s 69220 42168 70020 42288 6 wbs_dat_o[31]
port 97 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[3]
port 98 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[4]
port 99 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 wbs_dat_o[5]
port 100 nsew signal output
rlabel metal3 s 69220 44888 70020 45008 6 wbs_dat_o[6]
port 101 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[7]
port 102 nsew signal output
rlabel metal2 s 54758 71364 54814 72164 6 wbs_dat_o[8]
port 103 nsew signal output
rlabel metal2 s 52182 71364 52238 72164 6 wbs_dat_o[9]
port 104 nsew signal output
rlabel metal2 s 3238 71364 3294 72164 6 wbs_sel_i[0]
port 105 nsew signal input
rlabel metal2 s 13542 71364 13598 72164 6 wbs_sel_i[1]
port 106 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_sel_i[2]
port 107 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 wbs_sel_i[3]
port 108 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 wbs_stb_i
port 109 nsew signal input
rlabel metal3 s 69220 34008 70020 34128 6 wbs_we_i
port 110 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70020 72164
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11385362
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/wbuart32/runs/wbuart32/results/signoff/wbuart_wrap.magic.gds
string GDS_START 1122860
<< end >>

