magic
tech sky130A
magscale 1 2
timestamp 1654713702
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 348786 700544 348792 700596
rect 348844 700584 348850 700596
rect 357618 700584 357624 700596
rect 348844 700556 357624 700584
rect 348844 700544 348850 700556
rect 357618 700544 357624 700556
rect 357676 700544 357682 700596
rect 332502 700476 332508 700528
rect 332560 700516 332566 700528
rect 358814 700516 358820 700528
rect 332560 700488 358820 700516
rect 332560 700476 332566 700488
rect 358814 700476 358820 700488
rect 358872 700476 358878 700528
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 357526 700448 357532 700460
rect 300176 700420 357532 700448
rect 300176 700408 300182 700420
rect 357526 700408 357532 700420
rect 357584 700408 357590 700460
rect 283834 700340 283840 700392
rect 283892 700380 283898 700392
rect 358906 700380 358912 700392
rect 283892 700352 358912 700380
rect 283892 700340 283898 700352
rect 358906 700340 358912 700352
rect 358964 700340 358970 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 21358 700312 21364 700324
rect 8168 700284 21364 700312
rect 8168 700272 8174 700284
rect 21358 700272 21364 700284
rect 21416 700272 21422 700324
rect 217962 700272 217968 700324
rect 218020 700312 218026 700324
rect 235166 700312 235172 700324
rect 218020 700284 235172 700312
rect 218020 700272 218026 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 357434 700312 357440 700324
rect 267700 700284 357440 700312
rect 267700 700272 267706 700284
rect 357434 700272 357440 700284
rect 357492 700272 357498 700324
rect 359458 700272 359464 700324
rect 359516 700312 359522 700324
rect 397454 700312 397460 700324
rect 359516 700284 397460 700312
rect 359516 700272 359522 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 467098 700272 467104 700324
rect 467156 700312 467162 700324
rect 527174 700312 527180 700324
rect 467156 700284 527180 700312
rect 467156 700272 467162 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 527818 700272 527824 700324
rect 527876 700312 527882 700324
rect 559650 700312 559656 700324
rect 527876 700284 559656 700312
rect 527876 700272 527882 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 371878 696940 371884 696992
rect 371936 696980 371942 696992
rect 580166 696980 580172 696992
rect 371936 696952 580172 696980
rect 371936 696940 371942 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 18598 670732 18604 670744
rect 3568 670704 18604 670732
rect 3568 670692 3574 670704
rect 18598 670692 18604 670704
rect 18656 670692 18662 670744
rect 360838 670692 360844 670744
rect 360896 670732 360902 670744
rect 580166 670732 580172 670744
rect 360896 670704 580172 670732
rect 360896 670692 360902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 17218 656928 17224 656940
rect 3476 656900 17224 656928
rect 3476 656888 3482 656900
rect 17218 656888 17224 656900
rect 17276 656888 17282 656940
rect 367738 643084 367744 643136
rect 367796 643124 367802 643136
rect 580166 643124 580172 643136
rect 367796 643096 580172 643124
rect 367796 643084 367802 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 13078 632108 13084 632120
rect 3476 632080 13084 632108
rect 3476 632068 3482 632080
rect 13078 632068 13084 632080
rect 13136 632068 13142 632120
rect 373258 630640 373264 630692
rect 373316 630680 373322 630692
rect 579982 630680 579988 630692
rect 373316 630652 579988 630680
rect 373316 630640 373322 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 378778 616836 378784 616888
rect 378836 616876 378842 616888
rect 580166 616876 580172 616888
rect 378836 616848 580172 616876
rect 378836 616836 378842 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 606024 3516 606076
rect 3568 606064 3574 606076
rect 7558 606064 7564 606076
rect 3568 606036 7564 606064
rect 3568 606024 3574 606036
rect 7558 606024 7564 606036
rect 7616 606024 7622 606076
rect 363598 590656 363604 590708
rect 363656 590696 363662 590708
rect 580166 590696 580172 590708
rect 363656 590668 580172 590696
rect 363656 590656 363662 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 10318 579680 10324 579692
rect 3384 579652 10324 579680
rect 3384 579640 3390 579652
rect 10318 579640 10324 579652
rect 10376 579640 10382 579692
rect 369118 576852 369124 576904
rect 369176 576892 369182 576904
rect 580166 576892 580172 576904
rect 369176 576864 580172 576892
rect 369176 576852 369182 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 381538 563048 381544 563100
rect 381596 563088 381602 563100
rect 580166 563088 580172 563100
rect 381596 563060 580172 563088
rect 381596 563048 381602 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3602 553392 3608 553444
rect 3660 553432 3666 553444
rect 22738 553432 22744 553444
rect 3660 553404 22744 553432
rect 3660 553392 3666 553404
rect 22738 553392 22744 553404
rect 22796 553392 22802 553444
rect 498838 536800 498844 536852
rect 498896 536840 498902 536852
rect 579890 536840 579896 536852
rect 498896 536812 579896 536840
rect 498896 536800 498902 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 14458 527184 14464 527196
rect 3016 527156 14464 527184
rect 3016 527144 3022 527156
rect 14458 527144 14464 527156
rect 14516 527144 14522 527196
rect 3326 501304 3332 501356
rect 3384 501344 3390 501356
rect 8938 501344 8944 501356
rect 3384 501316 8944 501344
rect 3384 501304 3390 501316
rect 8938 501304 8944 501316
rect 8996 501304 9002 501356
rect 480898 484372 480904 484424
rect 480956 484412 480962 484424
rect 580166 484412 580172 484424
rect 480956 484384 580172 484412
rect 480956 484372 480962 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 217318 478864 217324 478916
rect 217376 478904 217382 478916
rect 220078 478904 220084 478916
rect 217376 478876 220084 478904
rect 217376 478864 217382 478876
rect 220078 478864 220084 478876
rect 220136 478864 220142 478916
rect 219066 478252 219072 478304
rect 219124 478292 219130 478304
rect 238754 478292 238760 478304
rect 219124 478264 238760 478292
rect 219124 478252 219130 478264
rect 238754 478252 238760 478264
rect 238812 478252 238818 478304
rect 217594 478184 217600 478236
rect 217652 478224 217658 478236
rect 248506 478224 248512 478236
rect 217652 478196 248512 478224
rect 217652 478184 217658 478196
rect 248506 478184 248512 478196
rect 248564 478184 248570 478236
rect 309134 478184 309140 478236
rect 309192 478224 309198 478236
rect 357618 478224 357624 478236
rect 309192 478196 357624 478224
rect 309192 478184 309198 478196
rect 357618 478184 357624 478196
rect 357676 478184 357682 478236
rect 218054 478116 218060 478168
rect 218112 478156 218118 478168
rect 314746 478156 314752 478168
rect 218112 478128 314752 478156
rect 218112 478116 218118 478128
rect 314746 478116 314752 478128
rect 314804 478116 314810 478168
rect 245746 476960 245752 477012
rect 245804 477000 245810 477012
rect 247034 477000 247040 477012
rect 245804 476972 247040 477000
rect 245804 476960 245810 476972
rect 247034 476960 247040 476972
rect 247092 476960 247098 477012
rect 258074 476960 258080 477012
rect 258132 477000 258138 477012
rect 262214 477000 262220 477012
rect 258132 476972 262220 477000
rect 258132 476960 258138 476972
rect 262214 476960 262220 476972
rect 262272 476960 262278 477012
rect 217502 476756 217508 476808
rect 217560 476796 217566 476808
rect 230474 476796 230480 476808
rect 217560 476768 230480 476796
rect 217560 476756 217566 476768
rect 230474 476756 230480 476768
rect 230532 476756 230538 476808
rect 233234 476688 233240 476740
rect 233292 476728 233298 476740
rect 242894 476728 242900 476740
rect 233292 476700 242900 476728
rect 233292 476688 233298 476700
rect 242894 476688 242900 476700
rect 242952 476688 242958 476740
rect 247310 476688 247316 476740
rect 247368 476728 247374 476740
rect 248414 476728 248420 476740
rect 247368 476700 248420 476728
rect 247368 476688 247374 476700
rect 248414 476688 248420 476700
rect 248472 476688 248478 476740
rect 258074 476688 258080 476740
rect 258132 476728 258138 476740
rect 258718 476728 258724 476740
rect 258132 476700 258724 476728
rect 258132 476688 258138 476700
rect 258718 476688 258724 476700
rect 258776 476688 258782 476740
rect 291194 476688 291200 476740
rect 291252 476728 291258 476740
rect 325786 476728 325792 476740
rect 291252 476700 325792 476728
rect 291252 476688 291258 476700
rect 325786 476688 325792 476700
rect 325844 476688 325850 476740
rect 278774 476620 278780 476672
rect 278832 476660 278838 476672
rect 304994 476660 305000 476672
rect 278832 476632 305000 476660
rect 278832 476620 278838 476632
rect 304994 476620 305000 476632
rect 305052 476620 305058 476672
rect 240134 476552 240140 476604
rect 240192 476592 240198 476604
rect 252554 476592 252560 476604
rect 240192 476564 252560 476592
rect 240192 476552 240198 476564
rect 252554 476552 252560 476564
rect 252612 476552 252618 476604
rect 252646 476552 252652 476604
rect 252704 476592 252710 476604
rect 264974 476592 264980 476604
rect 252704 476564 264980 476592
rect 252704 476552 252710 476564
rect 264974 476552 264980 476564
rect 265032 476552 265038 476604
rect 280154 476552 280160 476604
rect 280212 476592 280218 476604
rect 307754 476592 307760 476604
rect 280212 476564 307760 476592
rect 280212 476552 280218 476564
rect 307754 476552 307760 476564
rect 307812 476552 307818 476604
rect 233326 476484 233332 476536
rect 233384 476524 233390 476536
rect 247034 476524 247040 476536
rect 233384 476496 247040 476524
rect 233384 476484 233390 476496
rect 247034 476484 247040 476496
rect 247092 476484 247098 476536
rect 248506 476484 248512 476536
rect 248564 476524 248570 476536
rect 260834 476524 260840 476536
rect 248564 476496 260840 476524
rect 248564 476484 248570 476496
rect 260834 476484 260840 476496
rect 260892 476484 260898 476536
rect 260926 476484 260932 476536
rect 260984 476524 260990 476536
rect 277946 476524 277952 476536
rect 260984 476496 277952 476524
rect 260984 476484 260990 476496
rect 277946 476484 277952 476496
rect 278004 476484 278010 476536
rect 281534 476484 281540 476536
rect 281592 476524 281598 476536
rect 310514 476524 310520 476536
rect 281592 476496 310520 476524
rect 281592 476484 281598 476496
rect 310514 476484 310520 476496
rect 310572 476484 310578 476536
rect 237466 476416 237472 476468
rect 237524 476456 237530 476468
rect 239122 476456 239128 476468
rect 237524 476428 239128 476456
rect 237524 476416 237530 476428
rect 239122 476416 239128 476428
rect 239180 476416 239186 476468
rect 241422 476416 241428 476468
rect 241480 476456 241486 476468
rect 244274 476456 244280 476468
rect 241480 476428 244280 476456
rect 241480 476416 241486 476428
rect 244274 476416 244280 476428
rect 244332 476416 244338 476468
rect 255314 476416 255320 476468
rect 255372 476456 255378 476468
rect 268010 476456 268016 476468
rect 255372 476428 268016 476456
rect 255372 476416 255378 476428
rect 268010 476416 268016 476428
rect 268068 476416 268074 476468
rect 282914 476416 282920 476468
rect 282972 476456 282978 476468
rect 313274 476456 313280 476468
rect 282972 476428 313280 476456
rect 282972 476416 282978 476428
rect 313274 476416 313280 476428
rect 313332 476416 313338 476468
rect 249794 476388 249800 476400
rect 238726 476360 249800 476388
rect 231854 476280 231860 476332
rect 231912 476320 231918 476332
rect 235994 476320 236000 476332
rect 231912 476292 236000 476320
rect 231912 476280 231918 476292
rect 235994 476280 236000 476292
rect 236052 476280 236058 476332
rect 236178 476280 236184 476332
rect 236236 476320 236242 476332
rect 238726 476320 238754 476360
rect 249794 476348 249800 476360
rect 249852 476348 249858 476400
rect 251266 476348 251272 476400
rect 251324 476388 251330 476400
rect 263594 476388 263600 476400
rect 251324 476360 263600 476388
rect 251324 476348 251330 476360
rect 263594 476348 263600 476360
rect 263652 476348 263658 476400
rect 284294 476348 284300 476400
rect 284352 476388 284358 476400
rect 314654 476388 314660 476400
rect 284352 476360 314660 476388
rect 284352 476348 284358 476360
rect 314654 476348 314660 476360
rect 314712 476348 314718 476400
rect 236236 476292 238754 476320
rect 236236 476280 236242 476292
rect 242894 476280 242900 476332
rect 242952 476320 242958 476332
rect 242952 476292 253934 476320
rect 242952 476280 242958 476292
rect 236086 476212 236092 476264
rect 236144 476252 236150 476264
rect 236144 476224 238754 476252
rect 236144 476212 236150 476224
rect 234614 476144 234620 476196
rect 234672 476184 234678 476196
rect 237374 476184 237380 476196
rect 234672 476156 237380 476184
rect 234672 476144 234678 476156
rect 237374 476144 237380 476156
rect 237432 476144 237438 476196
rect 238726 476184 238754 476224
rect 238846 476212 238852 476264
rect 238904 476252 238910 476264
rect 244642 476252 244648 476264
rect 238904 476224 244648 476252
rect 238904 476212 238910 476224
rect 244642 476212 244648 476224
rect 244700 476212 244706 476264
rect 253906 476252 253934 476292
rect 256786 476280 256792 476332
rect 256844 476320 256850 476332
rect 270494 476320 270500 476332
rect 256844 476292 270500 476320
rect 256844 476280 256850 476292
rect 270494 476280 270500 476292
rect 270552 476280 270558 476332
rect 285674 476280 285680 476332
rect 285732 476320 285738 476332
rect 317414 476320 317420 476332
rect 285732 476292 317420 476320
rect 285732 476280 285738 476292
rect 317414 476280 317420 476292
rect 317472 476280 317478 476332
rect 255406 476252 255412 476264
rect 253906 476224 255412 476252
rect 255406 476212 255412 476224
rect 255464 476212 255470 476264
rect 258166 476212 258172 476264
rect 258224 476252 258230 476264
rect 273254 476252 273260 476264
rect 258224 476224 273260 476252
rect 258224 476212 258230 476224
rect 273254 476212 273260 476224
rect 273312 476212 273318 476264
rect 288434 476212 288440 476264
rect 288492 476252 288498 476264
rect 320174 476252 320180 476264
rect 288492 476224 320180 476252
rect 288492 476212 288498 476224
rect 320174 476212 320180 476224
rect 320232 476212 320238 476264
rect 241422 476184 241428 476196
rect 238726 476156 241428 476184
rect 241422 476144 241428 476156
rect 241480 476144 241486 476196
rect 241514 476144 241520 476196
rect 241572 476184 241578 476196
rect 245654 476184 245660 476196
rect 241572 476156 245660 476184
rect 241572 476144 241578 476156
rect 245654 476144 245660 476156
rect 245712 476144 245718 476196
rect 252370 476144 252376 476196
rect 252428 476184 252434 476196
rect 253934 476184 253940 476196
rect 252428 476156 253940 476184
rect 252428 476144 252434 476156
rect 253934 476144 253940 476156
rect 253992 476144 253998 476196
rect 259546 476144 259552 476196
rect 259604 476184 259610 476196
rect 276014 476184 276020 476196
rect 259604 476156 276020 476184
rect 259604 476144 259610 476156
rect 276014 476144 276020 476156
rect 276072 476144 276078 476196
rect 289814 476144 289820 476196
rect 289872 476184 289878 476196
rect 322934 476184 322940 476196
rect 289872 476156 322940 476184
rect 289872 476144 289878 476156
rect 322934 476144 322940 476156
rect 322992 476144 322998 476196
rect 234706 476076 234712 476128
rect 234764 476116 234770 476128
rect 235994 476116 236000 476128
rect 234764 476088 236000 476116
rect 234764 476076 234770 476088
rect 235994 476076 236000 476088
rect 236052 476076 236058 476128
rect 236178 476116 236184 476128
rect 236104 476088 236184 476116
rect 235994 475940 236000 475992
rect 236052 475980 236058 475992
rect 236104 475980 236132 476088
rect 236178 476076 236184 476088
rect 236236 476076 236242 476128
rect 242802 476076 242808 476128
rect 242860 476116 242866 476128
rect 244274 476116 244280 476128
rect 242860 476088 244280 476116
rect 242860 476076 242866 476088
rect 244274 476076 244280 476088
rect 244332 476076 244338 476128
rect 245838 476076 245844 476128
rect 245896 476116 245902 476128
rect 258258 476116 258264 476128
rect 245896 476088 258264 476116
rect 245896 476076 245902 476088
rect 258258 476076 258264 476088
rect 258316 476076 258322 476128
rect 277578 476076 277584 476128
rect 277636 476116 277642 476128
rect 302234 476116 302240 476128
rect 277636 476088 302240 476116
rect 277636 476076 277642 476088
rect 302234 476076 302240 476088
rect 302292 476076 302298 476128
rect 236052 475952 236132 475980
rect 236052 475940 236058 475952
rect 219158 475328 219164 475380
rect 219216 475368 219222 475380
rect 247126 475368 247132 475380
rect 219216 475340 247132 475368
rect 219216 475328 219222 475340
rect 247126 475328 247132 475340
rect 247184 475328 247190 475380
rect 267550 475328 267556 475380
rect 267608 475368 267614 475380
rect 274634 475368 274640 475380
rect 267608 475340 274640 475368
rect 267608 475328 267614 475340
rect 274634 475328 274640 475340
rect 274692 475328 274698 475380
rect 301038 475328 301044 475380
rect 301096 475368 301102 475380
rect 580258 475368 580264 475380
rect 301096 475340 580264 475368
rect 301096 475328 301102 475340
rect 580258 475328 580264 475340
rect 580316 475328 580322 475380
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 331214 474756 331220 474768
rect 3384 474728 331220 474756
rect 3384 474716 3390 474728
rect 331214 474716 331220 474728
rect 331272 474716 331278 474768
rect 217778 474036 217784 474088
rect 217836 474076 217842 474088
rect 250438 474076 250444 474088
rect 217836 474048 250444 474076
rect 217836 474036 217842 474048
rect 250438 474036 250444 474048
rect 250496 474036 250502 474088
rect 276014 474036 276020 474088
rect 276072 474076 276078 474088
rect 300854 474076 300860 474088
rect 276072 474048 300860 474076
rect 276072 474036 276078 474048
rect 300854 474036 300860 474048
rect 300912 474036 300918 474088
rect 320174 474036 320180 474088
rect 320232 474076 320238 474088
rect 498838 474076 498844 474088
rect 320232 474048 498844 474076
rect 320232 474036 320238 474048
rect 498838 474036 498844 474048
rect 498896 474036 498902 474088
rect 21358 473968 21364 474020
rect 21416 474008 21422 474020
rect 347866 474008 347872 474020
rect 21416 473980 347872 474008
rect 21416 473968 21422 473980
rect 347866 473968 347872 473980
rect 347924 473968 347930 474020
rect 217870 472676 217876 472728
rect 217928 472716 217934 472728
rect 254026 472716 254032 472728
rect 217928 472688 254032 472716
rect 217928 472676 217934 472688
rect 254026 472676 254032 472688
rect 254084 472676 254090 472728
rect 269206 472676 269212 472728
rect 269264 472716 269270 472728
rect 289906 472716 289912 472728
rect 269264 472688 289912 472716
rect 269264 472676 269270 472688
rect 289906 472676 289912 472688
rect 289964 472676 289970 472728
rect 71774 472608 71780 472660
rect 71832 472648 71838 472660
rect 346486 472648 346492 472660
rect 71832 472620 346492 472648
rect 71832 472608 71838 472620
rect 346486 472608 346492 472620
rect 346544 472608 346550 472660
rect 298094 471316 298100 471368
rect 298152 471356 298158 471368
rect 373258 471356 373264 471368
rect 298152 471328 373264 471356
rect 298152 471316 298158 471328
rect 373258 471316 373264 471328
rect 373316 471316 373322 471368
rect 14458 471248 14464 471300
rect 14516 471288 14522 471300
rect 328454 471288 328460 471300
rect 14516 471260 328460 471288
rect 14516 471248 14522 471260
rect 328454 471248 328460 471260
rect 328512 471248 328518 471300
rect 267734 469888 267740 469940
rect 267792 469928 267798 469940
rect 287054 469928 287060 469940
rect 267792 469900 287060 469928
rect 267792 469888 267798 469900
rect 287054 469888 287060 469900
rect 287112 469888 287118 469940
rect 10318 469820 10324 469872
rect 10376 469860 10382 469872
rect 327074 469860 327080 469872
rect 10376 469832 327080 469860
rect 10376 469820 10382 469832
rect 327074 469820 327080 469832
rect 327132 469820 327138 469872
rect 334066 469820 334072 469872
rect 334124 469860 334130 469872
rect 359458 469860 359464 469872
rect 334124 469832 359464 469860
rect 334124 469820 334130 469832
rect 359458 469820 359464 469832
rect 359516 469820 359522 469872
rect 266446 468528 266452 468580
rect 266504 468568 266510 468580
rect 285766 468568 285772 468580
rect 266504 468540 285772 468568
rect 266504 468528 266510 468540
rect 285766 468528 285772 468540
rect 285824 468528 285830 468580
rect 13078 468460 13084 468512
rect 13136 468500 13142 468512
rect 324314 468500 324320 468512
rect 13136 468472 324320 468500
rect 13136 468460 13142 468472
rect 324314 468460 324320 468472
rect 324372 468460 324378 468512
rect 329834 468460 329840 468512
rect 329892 468500 329898 468512
rect 467098 468500 467104 468512
rect 329892 468472 467104 468500
rect 329892 468460 329898 468472
rect 467098 468460 467104 468472
rect 467156 468460 467162 468512
rect 295334 467168 295340 467220
rect 295392 467208 295398 467220
rect 369118 467208 369124 467220
rect 295392 467180 369124 467208
rect 295392 467168 295398 467180
rect 369118 467168 369124 467180
rect 369176 467168 369182 467220
rect 4798 467100 4804 467152
rect 4856 467140 4862 467152
rect 321554 467140 321560 467152
rect 4856 467112 321560 467140
rect 4856 467100 4862 467112
rect 321554 467100 321560 467112
rect 321612 467100 321618 467152
rect 169754 465672 169760 465724
rect 169812 465712 169818 465724
rect 314746 465712 314752 465724
rect 169812 465684 314752 465712
rect 169812 465672 169818 465684
rect 314746 465672 314752 465684
rect 314804 465672 314810 465724
rect 327166 465672 327172 465724
rect 327224 465712 327230 465724
rect 371878 465712 371884 465724
rect 327224 465684 371884 465712
rect 327224 465672 327230 465684
rect 371878 465672 371884 465684
rect 371936 465672 371942 465724
rect 304994 464380 305000 464432
rect 305052 464420 305058 464432
rect 428458 464420 428464 464432
rect 305052 464392 428464 464420
rect 305052 464380 305058 464392
rect 428458 464380 428464 464392
rect 428516 464380 428522 464432
rect 22738 464312 22744 464364
rect 22796 464352 22802 464364
rect 351914 464352 351920 464364
rect 22796 464324 351920 464352
rect 22796 464312 22802 464324
rect 351914 464312 351920 464324
rect 351972 464312 351978 464364
rect 271874 462952 271880 463004
rect 271932 462992 271938 463004
rect 295426 462992 295432 463004
rect 271932 462964 295432 462992
rect 271932 462952 271938 462964
rect 295426 462952 295432 462964
rect 295484 462952 295490 463004
rect 332594 462952 332600 463004
rect 332652 462992 332658 463004
rect 462314 462992 462320 463004
rect 332652 462964 462320 462992
rect 332652 462952 332658 462964
rect 462314 462952 462320 462964
rect 462372 462952 462378 463004
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 332686 462380 332692 462392
rect 3384 462352 332692 462380
rect 3384 462340 3390 462352
rect 332686 462340 332692 462352
rect 332744 462340 332750 462392
rect 273162 461728 273168 461780
rect 273220 461768 273226 461780
rect 280338 461768 280344 461780
rect 273220 461740 280344 461768
rect 273220 461728 273226 461740
rect 280338 461728 280344 461740
rect 280396 461728 280402 461780
rect 277302 461660 277308 461712
rect 277360 461700 277366 461712
rect 287054 461700 287060 461712
rect 277360 461672 287060 461700
rect 277360 461660 277366 461672
rect 287054 461660 287060 461672
rect 287112 461660 287118 461712
rect 219250 461592 219256 461644
rect 219308 461632 219314 461644
rect 241606 461632 241612 461644
rect 219308 461604 241612 461632
rect 219308 461592 219314 461604
rect 241606 461592 241612 461604
rect 241664 461592 241670 461644
rect 263686 461592 263692 461644
rect 263744 461632 263750 461644
rect 280246 461632 280252 461644
rect 263744 461604 280252 461632
rect 263744 461592 263750 461604
rect 280246 461592 280252 461604
rect 280304 461592 280310 461644
rect 317414 461592 317420 461644
rect 317472 461632 317478 461644
rect 480898 461632 480904 461644
rect 317472 461604 480904 461632
rect 317472 461592 317478 461604
rect 480898 461592 480904 461604
rect 480956 461592 480962 461644
rect 322934 460232 322940 460284
rect 322992 460272 322998 460284
rect 363598 460272 363604 460284
rect 322992 460244 363604 460272
rect 322992 460232 322998 460244
rect 363598 460232 363604 460244
rect 363656 460232 363662 460284
rect 17218 460164 17224 460216
rect 17276 460204 17282 460216
rect 350074 460204 350080 460216
rect 17276 460176 350080 460204
rect 17276 460164 17282 460176
rect 350074 460164 350080 460176
rect 350132 460164 350138 460216
rect 308122 458872 308128 458924
rect 308180 458912 308186 458924
rect 364334 458912 364340 458924
rect 308180 458884 364340 458912
rect 308180 458872 308186 458884
rect 364334 458872 364340 458884
rect 364392 458872 364398 458924
rect 7558 458804 7564 458856
rect 7616 458844 7622 458856
rect 350810 458844 350816 458856
rect 7616 458816 350816 458844
rect 7616 458804 7622 458816
rect 350810 458804 350816 458816
rect 350868 458804 350874 458856
rect 303614 457512 303620 457564
rect 303672 457552 303678 457564
rect 494054 457552 494060 457564
rect 303672 457524 494060 457552
rect 303672 457512 303678 457524
rect 494054 457512 494060 457524
rect 494112 457512 494118 457564
rect 8938 457444 8944 457496
rect 8996 457484 9002 457496
rect 352282 457484 352288 457496
rect 8996 457456 352288 457484
rect 8996 457444 9002 457456
rect 352282 457444 352288 457456
rect 352340 457444 352346 457496
rect 270954 456084 270960 456136
rect 271012 456124 271018 456136
rect 292574 456124 292580 456136
rect 271012 456096 292580 456124
rect 271012 456084 271018 456096
rect 292574 456084 292580 456096
rect 292632 456084 292638 456136
rect 300946 456084 300952 456136
rect 301004 456124 301010 456136
rect 527818 456124 527824 456136
rect 301004 456096 527824 456124
rect 301004 456084 301010 456096
rect 527818 456084 527824 456096
rect 527876 456084 527882 456136
rect 18598 456016 18604 456068
rect 18656 456056 18662 456068
rect 323578 456056 323584 456068
rect 18656 456028 323584 456056
rect 18656 456016 18662 456028
rect 323578 456016 323584 456028
rect 323636 456016 323642 456068
rect 269022 455336 269028 455388
rect 269080 455376 269086 455388
rect 276474 455376 276480 455388
rect 269080 455348 276480 455376
rect 269080 455336 269086 455348
rect 276474 455336 276480 455348
rect 276532 455336 276538 455388
rect 274450 454724 274456 454776
rect 274508 454764 274514 454776
rect 283006 454764 283012 454776
rect 274508 454736 283012 454764
rect 274508 454724 274514 454736
rect 283006 454724 283012 454736
rect 283064 454724 283070 454776
rect 278682 454656 278688 454708
rect 278740 454696 278746 454708
rect 288802 454696 288808 454708
rect 278740 454668 288808 454696
rect 278740 454656 278746 454668
rect 288802 454656 288808 454668
rect 288860 454656 288866 454708
rect 298922 454656 298928 454708
rect 298980 454696 298986 454708
rect 360838 454696 360844 454708
rect 298980 454668 360844 454696
rect 298980 454656 298986 454668
rect 360838 454656 360844 454668
rect 360896 454656 360902 454708
rect 274082 453364 274088 453416
rect 274140 453404 274146 453416
rect 298186 453404 298192 453416
rect 274140 453376 298192 453404
rect 274140 453364 274146 453376
rect 298186 453364 298192 453376
rect 298244 453364 298250 453416
rect 217686 453296 217692 453348
rect 217744 453336 217750 453348
rect 231946 453336 231952 453348
rect 217744 453308 231952 453336
rect 217744 453296 217750 453308
rect 231946 453296 231952 453308
rect 232004 453296 232010 453348
rect 267642 453296 267648 453348
rect 267700 453336 267706 453348
rect 273254 453336 273260 453348
rect 267700 453308 273260 453336
rect 267700 453296 267706 453308
rect 273254 453296 273260 453308
rect 273312 453296 273318 453348
rect 275922 453296 275928 453348
rect 275980 453336 275986 453348
rect 285766 453336 285772 453348
rect 275980 453308 285772 453336
rect 275980 453296 275986 453308
rect 285766 453296 285772 453308
rect 285824 453296 285830 453348
rect 296714 453296 296720 453348
rect 296772 453336 296778 453348
rect 378778 453336 378784 453348
rect 296772 453308 378784 453336
rect 296772 453296 296778 453308
rect 378778 453296 378784 453308
rect 378836 453296 378842 453348
rect 271782 452752 271788 452804
rect 271840 452792 271846 452804
rect 279418 452792 279424 452804
rect 271840 452764 279424 452792
rect 271840 452752 271846 452764
rect 279418 452752 279424 452764
rect 279476 452752 279482 452804
rect 270402 451936 270408 451988
rect 270460 451976 270466 451988
rect 277486 451976 277492 451988
rect 270460 451948 277492 451976
rect 270460 451936 270466 451948
rect 277486 451936 277492 451948
rect 277544 451936 277550 451988
rect 280062 451936 280068 451988
rect 280120 451976 280126 451988
rect 290274 451976 290280 451988
rect 280120 451948 290280 451976
rect 280120 451936 280126 451948
rect 290274 451936 290280 451948
rect 290332 451936 290338 451988
rect 219342 451868 219348 451920
rect 219400 451908 219406 451920
rect 244642 451908 244648 451920
rect 219400 451880 244648 451908
rect 219400 451868 219406 451880
rect 244642 451868 244648 451880
rect 244700 451868 244706 451920
rect 266262 451868 266268 451920
rect 266320 451908 266326 451920
rect 271966 451908 271972 451920
rect 266320 451880 271972 451908
rect 266320 451868 266326 451880
rect 271966 451868 271972 451880
rect 272024 451868 272030 451920
rect 274542 451868 274548 451920
rect 274600 451908 274606 451920
rect 284386 451908 284392 451920
rect 274600 451880 284392 451908
rect 274600 451868 274606 451880
rect 284386 451868 284392 451880
rect 284444 451868 284450 451920
rect 294138 451868 294144 451920
rect 294196 451908 294202 451920
rect 381538 451908 381544 451920
rect 294196 451880 381544 451908
rect 294196 451868 294202 451880
rect 381538 451868 381544 451880
rect 381596 451868 381602 451920
rect 265158 450576 265164 450628
rect 265216 450616 265222 450628
rect 283098 450616 283104 450628
rect 265216 450588 283104 450616
rect 265216 450576 265222 450588
rect 283098 450576 283104 450588
rect 283156 450576 283162 450628
rect 325602 450576 325608 450628
rect 325660 450616 325666 450628
rect 367738 450616 367744 450628
rect 325660 450588 367744 450616
rect 325660 450576 325666 450588
rect 367738 450576 367744 450588
rect 367796 450576 367802 450628
rect 3602 450508 3608 450560
rect 3660 450548 3666 450560
rect 331030 450548 331036 450560
rect 3660 450520 331036 450548
rect 3660 450508 3666 450520
rect 331030 450508 331036 450520
rect 331088 450508 331094 450560
rect 307846 449624 307852 449676
rect 307904 449664 307910 449676
rect 412634 449664 412640 449676
rect 307904 449636 412640 449664
rect 307904 449624 307910 449636
rect 412634 449624 412640 449636
rect 412692 449624 412698 449676
rect 153194 449556 153200 449608
rect 153252 449596 153258 449608
rect 317138 449596 317144 449608
rect 153252 449568 317144 449596
rect 153252 449556 153258 449568
rect 317138 449556 317144 449568
rect 317196 449556 317202 449608
rect 305454 449488 305460 449540
rect 305512 449528 305518 449540
rect 477494 449528 477500 449540
rect 305512 449500 477500 449528
rect 305512 449488 305518 449500
rect 477494 449488 477500 449500
rect 477552 449488 477558 449540
rect 88334 449420 88340 449472
rect 88392 449460 88398 449472
rect 319438 449460 319444 449472
rect 88392 449432 319444 449460
rect 88392 449420 88398 449432
rect 319438 449420 319444 449432
rect 319496 449420 319502 449472
rect 303154 449352 303160 449404
rect 303212 449392 303218 449404
rect 542354 449392 542360 449404
rect 303212 449364 542360 449392
rect 303212 449352 303218 449364
rect 542354 449352 542360 449364
rect 542412 449352 542418 449404
rect 23474 449284 23480 449336
rect 23532 449324 23538 449336
rect 321738 449324 321744 449336
rect 23532 449296 321744 449324
rect 23532 449284 23538 449296
rect 321738 449284 321744 449296
rect 321796 449284 321802 449336
rect 3418 449216 3424 449268
rect 3476 449256 3482 449268
rect 326430 449256 326436 449268
rect 3476 449228 326436 449256
rect 3476 449216 3482 449228
rect 326430 449216 326436 449228
rect 326488 449216 326494 449268
rect 3510 449148 3516 449200
rect 3568 449188 3574 449200
rect 328730 449188 328736 449200
rect 3568 449160 328736 449188
rect 3568 449148 3574 449160
rect 328730 449148 328736 449160
rect 328788 449148 328794 449200
rect 201494 448060 201500 448112
rect 201552 448100 201558 448112
rect 341886 448100 341892 448112
rect 201552 448072 341892 448100
rect 201552 448060 201558 448072
rect 341886 448060 341892 448072
rect 341944 448060 341950 448112
rect 136634 447992 136640 448044
rect 136692 448032 136698 448044
rect 344186 448032 344192 448044
rect 136692 448004 344192 448032
rect 136692 447992 136698 448004
rect 344186 447992 344192 448004
rect 344244 447992 344250 448044
rect 104894 447924 104900 447976
rect 104952 447964 104958 447976
rect 317874 447964 317880 447976
rect 104952 447936 317880 447964
rect 104952 447924 104958 447936
rect 317874 447924 317880 447936
rect 317932 447924 317938 447976
rect 40034 447856 40040 447908
rect 40092 447896 40098 447908
rect 320174 447896 320180 447908
rect 40092 447868 320180 447896
rect 40092 447856 40098 447868
rect 320174 447856 320180 447868
rect 320232 447856 320238 447908
rect 2866 447788 2872 447840
rect 2924 447828 2930 447840
rect 353478 447828 353484 447840
rect 2924 447800 353484 447828
rect 2924 447788 2930 447800
rect 353478 447788 353484 447800
rect 353536 447788 353542 447840
rect 255958 447040 255964 447092
rect 256016 447080 256022 447092
rect 258258 447080 258264 447092
rect 256016 447052 258264 447080
rect 256016 447040 256022 447052
rect 258258 447040 258264 447052
rect 258316 447040 258322 447092
rect 262858 447040 262864 447092
rect 262916 447080 262922 447092
rect 267550 447080 267556 447092
rect 262916 447052 267556 447080
rect 262916 447040 262922 447052
rect 267550 447040 267556 447052
rect 267608 447040 267614 447092
rect 231854 446972 231860 447024
rect 231912 447012 231918 447024
rect 232406 447012 232412 447024
rect 231912 446984 232412 447012
rect 231912 446972 231918 446984
rect 232406 446972 232412 446984
rect 232464 446972 232470 447024
rect 235994 446972 236000 447024
rect 236052 447012 236058 447024
rect 237006 447012 237012 447024
rect 236052 446984 237012 447012
rect 236052 446972 236058 446984
rect 237006 446972 237012 446984
rect 237064 446972 237070 447024
rect 241514 446972 241520 447024
rect 241572 447012 241578 447024
rect 242342 447012 242348 447024
rect 241572 446984 242348 447012
rect 241572 446972 241578 446984
rect 242342 446972 242348 446984
rect 242400 446972 242406 447024
rect 248414 446972 248420 447024
rect 248472 447012 248478 447024
rect 249334 447012 249340 447024
rect 248472 446984 249340 447012
rect 248472 446972 248478 446984
rect 249334 446972 249340 446984
rect 249392 446972 249398 447024
rect 250438 446972 250444 447024
rect 250496 447012 250502 447024
rect 252002 447012 252008 447024
rect 250496 446984 252008 447012
rect 250496 446972 250502 446984
rect 252002 446972 252008 446984
rect 252060 446972 252066 447024
rect 253934 446972 253940 447024
rect 253992 447012 253998 447024
rect 254854 447012 254860 447024
rect 253992 446984 254860 447012
rect 253992 446972 253998 446984
rect 254854 446972 254860 446984
rect 254912 446972 254918 447024
rect 256602 446972 256608 447024
rect 256660 447012 256666 447024
rect 259730 447012 259736 447024
rect 256660 446984 259736 447012
rect 256660 446972 256666 446984
rect 259730 446972 259736 446984
rect 259788 446972 259794 447024
rect 261478 446972 261484 447024
rect 261536 447012 261542 447024
rect 265986 447012 265992 447024
rect 261536 446984 265992 447012
rect 261536 446972 261542 446984
rect 265986 446972 265992 446984
rect 266044 446972 266050 447024
rect 271874 446972 271880 447024
rect 271932 447012 271938 447024
rect 272702 447012 272708 447024
rect 271932 446984 272708 447012
rect 271932 446972 271938 446984
rect 272702 446972 272708 446984
rect 272760 446972 272766 447024
rect 277486 446972 277492 447024
rect 277544 447012 277550 447024
rect 278038 447012 278044 447024
rect 277544 446984 278044 447012
rect 277544 446972 277550 446984
rect 278038 446972 278044 446984
rect 278096 446972 278102 447024
rect 282914 446972 282920 447024
rect 282972 447012 282978 447024
rect 283374 447012 283380 447024
rect 282972 446984 283380 447012
rect 282972 446972 282978 446984
rect 283374 446972 283380 446984
rect 283432 446972 283438 447024
rect 284294 446972 284300 447024
rect 284352 447012 284358 447024
rect 285030 447012 285036 447024
rect 284352 446984 285036 447012
rect 284352 446972 284358 446984
rect 285030 446972 285036 446984
rect 285088 446972 285094 447024
rect 285674 446972 285680 447024
rect 285732 447012 285738 447024
rect 286502 447012 286508 447024
rect 285732 446984 286508 447012
rect 285732 446972 285738 446984
rect 286502 446972 286508 446984
rect 286560 446972 286566 447024
rect 300946 446972 300952 447024
rect 301004 447012 301010 447024
rect 301222 447012 301228 447024
rect 301004 446984 301228 447012
rect 301004 446972 301010 446984
rect 301222 446972 301228 446984
rect 301280 446972 301286 447024
rect 264238 446904 264244 446956
rect 264296 446944 264302 446956
rect 269114 446944 269120 446956
rect 264296 446916 269120 446944
rect 264296 446904 264302 446916
rect 269114 446904 269120 446916
rect 269172 446904 269178 446956
rect 217962 446632 217968 446684
rect 218020 446672 218026 446684
rect 313182 446672 313188 446684
rect 218020 446644 313188 446672
rect 218020 446632 218026 446644
rect 313182 446632 313188 446644
rect 313240 446632 313246 446684
rect 339586 446632 339592 446684
rect 339644 446672 339650 446684
rect 357434 446672 357440 446684
rect 339644 446644 357440 446672
rect 339644 446632 339650 446644
rect 357434 446632 357440 446644
rect 357492 446632 357498 446684
rect 260742 446564 260748 446616
rect 260800 446604 260806 446616
rect 264422 446604 264428 446616
rect 260800 446576 264428 446604
rect 260800 446564 260806 446576
rect 264422 446564 264428 446576
rect 264480 446564 264486 446616
rect 302418 446564 302424 446616
rect 302476 446604 302482 446616
rect 333974 446604 333980 446616
rect 302476 446576 333980 446604
rect 302476 446564 302482 446576
rect 333974 446564 333980 446576
rect 334032 446564 334038 446616
rect 337194 446564 337200 446616
rect 337252 446604 337258 446616
rect 358814 446604 358820 446616
rect 337252 446576 358820 446604
rect 337252 446564 337258 446576
rect 358814 446564 358820 446576
rect 358872 446564 358878 446616
rect 312446 446496 312452 446548
rect 312504 446536 312510 446548
rect 358906 446536 358912 446548
rect 312504 446508 358912 446536
rect 312504 446496 312510 446508
rect 358906 446496 358912 446508
rect 358964 446496 358970 446548
rect 220078 446428 220084 446480
rect 220136 446468 220142 446480
rect 230382 446468 230388 446480
rect 220136 446440 230388 446468
rect 220136 446428 220142 446440
rect 230382 446428 230388 446440
rect 230440 446428 230446 446480
rect 265618 446428 265624 446480
rect 265676 446468 265682 446480
rect 270586 446468 270592 446480
rect 265676 446440 270592 446468
rect 265676 446428 265682 446440
rect 270586 446428 270592 446440
rect 270644 446428 270650 446480
rect 310882 446428 310888 446480
rect 310940 446468 310946 446480
rect 357526 446468 357532 446480
rect 310940 446440 357532 446468
rect 310940 446428 310946 446440
rect 357526 446428 357532 446440
rect 357584 446428 357590 446480
rect 311710 446360 311716 446412
rect 311768 446400 311774 446412
rect 362218 446400 362224 446412
rect 311768 446372 362224 446400
rect 311768 446360 311774 446372
rect 362218 446360 362224 446372
rect 362276 446360 362282 446412
rect 307018 446292 307024 446344
rect 307076 446332 307082 446344
rect 364978 446332 364984 446344
rect 307076 446304 364984 446332
rect 307076 446292 307082 446304
rect 364978 446292 364984 446304
rect 365036 446292 365042 446344
rect 253842 446224 253848 446276
rect 253900 446264 253906 446276
rect 256694 446264 256700 446276
rect 253900 446236 256700 446264
rect 253900 446224 253906 446236
rect 256694 446224 256700 446236
rect 256752 446224 256758 446276
rect 258718 446224 258724 446276
rect 258776 446264 258782 446276
rect 261294 446264 261300 446276
rect 258776 446236 261300 446264
rect 258776 446224 258782 446236
rect 261294 446224 261300 446236
rect 261352 446224 261358 446276
rect 304718 446224 304724 446276
rect 304776 446264 304782 446276
rect 363598 446264 363604 446276
rect 304776 446236 363604 446264
rect 304776 446224 304782 446236
rect 363598 446224 363604 446236
rect 363656 446224 363662 446276
rect 293126 446156 293132 446208
rect 293184 446196 293190 446208
rect 361022 446196 361028 446208
rect 293184 446168 361028 446196
rect 293184 446156 293190 446168
rect 361022 446156 361028 446168
rect 361080 446156 361086 446208
rect 292298 446088 292304 446140
rect 292356 446128 292362 446140
rect 373258 446128 373264 446140
rect 292356 446100 373264 446128
rect 292356 446088 292362 446100
rect 373258 446088 373264 446100
rect 373316 446088 373322 446140
rect 243538 446020 243544 446072
rect 243596 446060 243602 446072
rect 345014 446060 345020 446072
rect 243596 446032 345020 446060
rect 243596 446020 243602 446032
rect 345014 446020 345020 446032
rect 345072 446020 345078 446072
rect 229830 445952 229836 446004
rect 229888 445992 229894 446004
rect 338022 445992 338028 446004
rect 229888 445964 338028 445992
rect 229888 445952 229894 445964
rect 338022 445952 338028 445964
rect 338080 445952 338086 446004
rect 229738 445884 229744 445936
rect 229796 445924 229802 445936
rect 347314 445924 347320 445936
rect 229796 445896 347320 445924
rect 229796 445884 229802 445896
rect 347314 445884 347320 445896
rect 347372 445884 347378 445936
rect 228358 445816 228364 445868
rect 228416 445856 228422 445868
rect 349614 445856 349620 445868
rect 228416 445828 349620 445856
rect 228416 445816 228422 445828
rect 349614 445816 349620 445828
rect 349672 445816 349678 445868
rect 293862 445748 293868 445800
rect 293920 445788 293926 445800
rect 458818 445788 458824 445800
rect 293920 445760 458824 445788
rect 293920 445748 293926 445760
rect 458818 445748 458824 445760
rect 458876 445748 458882 445800
rect 228542 445204 228548 445256
rect 228600 445244 228606 445256
rect 336458 445244 336464 445256
rect 228600 445216 336464 445244
rect 228600 445204 228606 445216
rect 336458 445204 336464 445216
rect 336516 445204 336522 445256
rect 7558 445136 7564 445188
rect 7616 445176 7622 445188
rect 334158 445176 334164 445188
rect 7616 445148 334164 445176
rect 7616 445136 7622 445148
rect 334158 445136 334164 445148
rect 334216 445136 334222 445188
rect 225690 445068 225696 445120
rect 225748 445108 225754 445120
rect 338758 445108 338764 445120
rect 225748 445080 338764 445108
rect 225748 445068 225754 445080
rect 338758 445068 338764 445080
rect 338816 445068 338822 445120
rect 333974 445000 333980 445052
rect 334032 445040 334038 445052
rect 580258 445040 580264 445052
rect 334032 445012 580264 445040
rect 334032 445000 334038 445012
rect 580258 445000 580264 445012
rect 580316 445000 580322 445052
rect 224218 444932 224224 444984
rect 224276 444972 224282 444984
rect 341150 444972 341156 444984
rect 224276 444944 341156 444972
rect 224276 444932 224282 444944
rect 341150 444932 341156 444944
rect 341208 444932 341214 444984
rect 228450 444864 228456 444916
rect 228508 444904 228514 444916
rect 355870 444904 355876 444916
rect 228508 444876 355876 444904
rect 228508 444864 228514 444876
rect 355870 444864 355876 444876
rect 355928 444864 355934 444916
rect 300026 444796 300032 444848
rect 300084 444836 300090 444848
rect 442258 444836 442264 444848
rect 300084 444808 442264 444836
rect 300084 444796 300090 444808
rect 442258 444796 442264 444808
rect 442316 444796 442322 444848
rect 295426 444728 295432 444780
rect 295484 444768 295490 444780
rect 526438 444768 526444 444780
rect 295484 444740 526444 444768
rect 295484 444728 295490 444740
rect 526438 444728 526444 444740
rect 526496 444728 526502 444780
rect 93210 444660 93216 444712
rect 93268 444700 93274 444712
rect 343450 444700 343456 444712
rect 93268 444672 343456 444700
rect 93268 444660 93274 444672
rect 343450 444660 343456 444672
rect 343508 444660 343514 444712
rect 86218 444592 86224 444644
rect 86276 444632 86282 444644
rect 345750 444632 345756 444644
rect 86276 444604 345756 444632
rect 86276 444592 86282 444604
rect 345750 444592 345756 444604
rect 345808 444592 345814 444644
rect 84838 444524 84844 444576
rect 84896 444564 84902 444576
rect 348050 444564 348056 444576
rect 84896 444536 348056 444564
rect 84896 444524 84902 444536
rect 348050 444524 348056 444536
rect 348108 444524 348114 444576
rect 82078 444456 82084 444508
rect 82136 444496 82142 444508
rect 358170 444496 358176 444508
rect 82136 444468 358176 444496
rect 82136 444456 82142 444468
rect 358170 444456 358176 444468
rect 358228 444456 358234 444508
rect 314010 444388 314016 444440
rect 314068 444428 314074 444440
rect 369118 444428 369124 444440
rect 314068 444400 369124 444428
rect 314068 444388 314074 444400
rect 369118 444388 369124 444400
rect 369176 444388 369182 444440
rect 3510 443640 3516 443692
rect 3568 443680 3574 443692
rect 243538 443680 243544 443692
rect 3568 443652 243544 443680
rect 3568 443640 3574 443652
rect 243538 443640 243544 443652
rect 243596 443640 243602 443692
rect 309318 443640 309324 443692
rect 309376 443680 309382 443692
rect 309376 443652 316034 443680
rect 309376 443640 309382 443652
rect 316006 443544 316034 443652
rect 316310 443572 316316 443624
rect 316368 443612 316374 443624
rect 362310 443612 362316 443624
rect 316368 443584 362316 443612
rect 316368 443572 316374 443584
rect 362310 443572 362316 443584
rect 362368 443572 362374 443624
rect 367738 443544 367744 443556
rect 316006 443516 367744 443544
rect 367738 443504 367744 443516
rect 367796 443504 367802 443556
rect 226978 443436 226984 443488
rect 227036 443476 227042 443488
rect 335538 443476 335544 443488
rect 227036 443448 335544 443476
rect 227036 443436 227042 443448
rect 335538 443436 335544 443448
rect 335596 443436 335602 443488
rect 225598 443368 225604 443420
rect 225656 443408 225662 443420
rect 342254 443408 342260 443420
rect 225656 443380 342260 443408
rect 225656 443368 225662 443380
rect 342254 443368 342260 443380
rect 342312 443368 342318 443420
rect 221458 443300 221464 443352
rect 221516 443340 221522 443352
rect 340046 443340 340052 443352
rect 221516 443312 340052 443340
rect 221516 443300 221522 443312
rect 340046 443300 340052 443312
rect 340104 443300 340110 443352
rect 228634 443232 228640 443284
rect 228692 443272 228698 443284
rect 354030 443272 354036 443284
rect 228692 443244 354036 443272
rect 228692 443232 228698 443244
rect 354030 443232 354036 443244
rect 354088 443232 354094 443284
rect 220078 443164 220084 443216
rect 220136 443204 220142 443216
rect 354766 443204 354772 443216
rect 220136 443176 354772 443204
rect 220136 443164 220142 443176
rect 354766 443164 354772 443176
rect 354824 443164 354830 443216
rect 98638 443096 98644 443148
rect 98696 443136 98702 443148
rect 356238 443136 356244 443148
rect 98696 443108 356244 443136
rect 98696 443096 98702 443108
rect 356238 443096 356244 443108
rect 356296 443096 356302 443148
rect 95970 443028 95976 443080
rect 96028 443068 96034 443080
rect 356974 443068 356980 443080
rect 96028 443040 356980 443068
rect 96028 443028 96034 443040
rect 356974 443028 356980 443040
rect 357032 443028 357038 443080
rect 80698 442960 80704 443012
rect 80756 443000 80762 443012
rect 358814 443000 358820 443012
rect 80756 442972 358820 443000
rect 80756 442960 80762 442972
rect 358814 442960 358820 442972
rect 358872 442960 358878 443012
rect 3602 442212 3608 442264
rect 3660 442252 3666 442264
rect 229830 442252 229836 442264
rect 3660 442224 229836 442252
rect 3660 442212 3666 442224
rect 229830 442212 229836 442224
rect 229888 442212 229894 442264
rect 361022 442212 361028 442264
rect 361080 442252 361086 442264
rect 580994 442252 581000 442264
rect 361080 442224 581000 442252
rect 361080 442212 361086 442224
rect 580994 442212 581000 442224
rect 581052 442212 581058 442264
rect 3418 440852 3424 440904
rect 3476 440892 3482 440904
rect 229738 440892 229744 440904
rect 3476 440864 229744 440892
rect 3476 440852 3482 440864
rect 229738 440852 229744 440864
rect 229796 440852 229802 440904
rect 458818 439492 458824 439544
rect 458876 439532 458882 439544
rect 582374 439532 582380 439544
rect 458876 439504 582380 439532
rect 458876 439492 458882 439504
rect 582374 439492 582380 439504
rect 582432 439492 582438 439544
rect 362310 431876 362316 431928
rect 362368 431916 362374 431928
rect 580166 431916 580172 431928
rect 362368 431888 580172 431916
rect 362368 431876 362374 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 7558 423620 7564 423632
rect 3384 423592 7564 423620
rect 3384 423580 3390 423592
rect 7558 423580 7564 423592
rect 7616 423580 7622 423632
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 226978 411244 226984 411256
rect 3384 411216 226984 411244
rect 3384 411204 3390 411216
rect 226978 411204 226984 411216
rect 227036 411204 227042 411256
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 228634 398800 228640 398812
rect 3384 398772 228640 398800
rect 3384 398760 3390 398772
rect 228634 398760 228640 398772
rect 228692 398760 228698 398812
rect 369118 379448 369124 379500
rect 369176 379488 369182 379500
rect 580166 379488 580172 379500
rect 369176 379460 580172 379488
rect 369176 379448 369182 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3050 372512 3056 372564
rect 3108 372552 3114 372564
rect 228542 372552 228548 372564
rect 3108 372524 228548 372552
rect 3108 372512 3114 372524
rect 228542 372512 228548 372524
rect 228600 372512 228606 372564
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 220078 346372 220084 346384
rect 3384 346344 220084 346372
rect 3384 346332 3390 346344
rect 220078 346332 220084 346344
rect 220136 346332 220142 346384
rect 362218 325592 362224 325644
rect 362276 325632 362282 325644
rect 579890 325632 579896 325644
rect 362276 325604 579896 325632
rect 362276 325592 362282 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 225690 320124 225696 320136
rect 3384 320096 225696 320124
rect 3384 320084 3390 320096
rect 225690 320084 225696 320096
rect 225748 320084 225754 320136
rect 224954 309068 224960 309120
rect 225012 309108 225018 309120
rect 237190 309108 237196 309120
rect 225012 309080 237196 309108
rect 225012 309068 225018 309080
rect 237190 309068 237196 309080
rect 237248 309068 237254 309120
rect 290550 309068 290556 309120
rect 290608 309108 290614 309120
rect 349430 309108 349436 309120
rect 290608 309080 349436 309108
rect 290608 309068 290614 309080
rect 349430 309068 349436 309080
rect 349488 309068 349494 309120
rect 354858 309068 354864 309120
rect 354916 309108 354922 309120
rect 354916 309080 369854 309108
rect 354916 309068 354922 309080
rect 97258 309000 97264 309052
rect 97316 309040 97322 309052
rect 247678 309040 247684 309052
rect 97316 309012 247684 309040
rect 97316 309000 97322 309012
rect 247678 309000 247684 309012
rect 247736 309000 247742 309052
rect 281442 309000 281448 309052
rect 281500 309040 281506 309052
rect 281500 309012 287652 309040
rect 281500 309000 281506 309012
rect 68278 308932 68284 308984
rect 68336 308972 68342 308984
rect 234614 308972 234620 308984
rect 68336 308944 234620 308972
rect 68336 308932 68342 308944
rect 234614 308932 234620 308944
rect 234672 308932 234678 308984
rect 242250 308932 242256 308984
rect 242308 308972 242314 308984
rect 252186 308972 252192 308984
rect 242308 308944 252192 308972
rect 242308 308932 242314 308944
rect 252186 308932 252192 308944
rect 252244 308932 252250 308984
rect 263566 308944 278084 308972
rect 50338 308864 50344 308916
rect 50396 308904 50402 308916
rect 232866 308904 232872 308916
rect 50396 308876 232872 308904
rect 50396 308864 50402 308876
rect 232866 308864 232872 308876
rect 232924 308864 232930 308916
rect 64138 308796 64144 308848
rect 64196 308836 64202 308848
rect 233786 308836 233792 308848
rect 64196 308808 233792 308836
rect 64196 308796 64202 308808
rect 233786 308796 233792 308808
rect 233844 308796 233850 308848
rect 249334 308796 249340 308848
rect 249392 308836 249398 308848
rect 258258 308836 258264 308848
rect 249392 308808 258264 308836
rect 249392 308796 249398 308808
rect 258258 308796 258264 308808
rect 258316 308796 258322 308848
rect 46198 308728 46204 308780
rect 46256 308768 46262 308780
rect 232038 308768 232044 308780
rect 46256 308740 232044 308768
rect 46256 308728 46262 308740
rect 232038 308728 232044 308740
rect 232096 308728 232102 308780
rect 252002 308728 252008 308780
rect 252060 308768 252066 308780
rect 252060 308740 253888 308768
rect 252060 308728 252066 308740
rect 43438 308660 43444 308712
rect 43496 308700 43502 308712
rect 224954 308700 224960 308712
rect 43496 308672 224960 308700
rect 43496 308660 43502 308672
rect 224954 308660 224960 308672
rect 225012 308660 225018 308712
rect 236546 308700 236552 308712
rect 233620 308672 236552 308700
rect 39298 308592 39304 308644
rect 39356 308632 39362 308644
rect 233510 308632 233516 308644
rect 39356 308604 233516 308632
rect 39356 308592 39362 308604
rect 233510 308592 233516 308604
rect 233568 308592 233574 308644
rect 35894 308524 35900 308576
rect 35952 308564 35958 308576
rect 233620 308564 233648 308672
rect 236546 308660 236552 308672
rect 236604 308660 236610 308712
rect 252646 308700 252652 308712
rect 244246 308672 252652 308700
rect 241790 308632 241796 308644
rect 238726 308604 241796 308632
rect 235258 308564 235264 308576
rect 35952 308536 233648 308564
rect 234586 308536 235264 308564
rect 35952 308524 35958 308536
rect 27614 308456 27620 308508
rect 27672 308496 27678 308508
rect 234586 308496 234614 308536
rect 235258 308524 235264 308536
rect 235316 308524 235322 308576
rect 237098 308524 237104 308576
rect 237156 308564 237162 308576
rect 238726 308564 238754 308604
rect 241790 308592 241796 308604
rect 241848 308592 241854 308644
rect 243538 308592 243544 308644
rect 243596 308632 243602 308644
rect 244246 308632 244274 308672
rect 252646 308660 252652 308672
rect 252704 308660 252710 308712
rect 252738 308660 252744 308712
rect 252796 308700 252802 308712
rect 253566 308700 253572 308712
rect 252796 308672 253572 308700
rect 252796 308660 252802 308672
rect 253566 308660 253572 308672
rect 253624 308660 253630 308712
rect 253860 308700 253888 308740
rect 263566 308700 263594 308944
rect 268378 308728 268384 308780
rect 268436 308768 268442 308780
rect 275646 308768 275652 308780
rect 268436 308740 275652 308768
rect 268436 308728 268442 308740
rect 275646 308728 275652 308740
rect 275704 308728 275710 308780
rect 253860 308672 263594 308700
rect 264238 308660 264244 308712
rect 264296 308700 264302 308712
rect 276934 308700 276940 308712
rect 264296 308672 276940 308700
rect 264296 308660 264302 308672
rect 276934 308660 276940 308672
rect 276992 308660 276998 308712
rect 278056 308700 278084 308944
rect 281350 308932 281356 308984
rect 281408 308972 281414 308984
rect 287624 308972 287652 309012
rect 287698 309000 287704 309052
rect 287756 309040 287762 309052
rect 350810 309040 350816 309052
rect 287756 309012 350816 309040
rect 287756 309000 287762 309012
rect 350810 309000 350816 309012
rect 350868 309000 350874 309052
rect 354646 309012 360194 309040
rect 347314 308972 347320 308984
rect 281408 308944 284432 308972
rect 287624 308944 347320 308972
rect 281408 308932 281414 308944
rect 281166 308864 281172 308916
rect 281224 308904 281230 308916
rect 284404 308904 284432 308944
rect 347314 308932 347320 308944
rect 347372 308932 347378 308984
rect 347958 308904 347964 308916
rect 281224 308876 284340 308904
rect 284404 308876 347964 308904
rect 281224 308864 281230 308876
rect 284312 308836 284340 308876
rect 347958 308864 347964 308876
rect 348016 308864 348022 308916
rect 348602 308836 348608 308848
rect 284312 308808 348608 308836
rect 348602 308796 348608 308808
rect 348660 308796 348666 308848
rect 354214 308796 354220 308848
rect 354272 308836 354278 308848
rect 354646 308836 354674 309012
rect 354272 308808 354674 308836
rect 354272 308796 354278 308808
rect 355594 308796 355600 308848
rect 355652 308836 355658 308848
rect 360166 308836 360194 309012
rect 369826 308904 369854 309080
rect 438118 308904 438124 308916
rect 369826 308876 438124 308904
rect 438118 308864 438124 308876
rect 438176 308864 438182 308916
rect 436830 308836 436836 308848
rect 355652 308808 359872 308836
rect 360166 308808 436836 308836
rect 355652 308796 355658 308808
rect 282730 308728 282736 308780
rect 282788 308768 282794 308780
rect 353202 308768 353208 308780
rect 282788 308740 353208 308768
rect 282788 308728 282794 308740
rect 353202 308728 353208 308740
rect 353260 308728 353266 308780
rect 354674 308728 354680 308780
rect 354732 308768 354738 308780
rect 355410 308768 355416 308780
rect 354732 308740 355416 308768
rect 354732 308728 354738 308740
rect 355410 308728 355416 308740
rect 355468 308728 355474 308780
rect 356238 308728 356244 308780
rect 356296 308768 356302 308780
rect 356514 308768 356520 308780
rect 356296 308740 356520 308768
rect 356296 308728 356302 308740
rect 356514 308728 356520 308740
rect 356572 308728 356578 308780
rect 357434 308728 357440 308780
rect 357492 308768 357498 308780
rect 357894 308768 357900 308780
rect 357492 308740 357900 308768
rect 357492 308728 357498 308740
rect 357894 308728 357900 308740
rect 357952 308728 357958 308780
rect 359844 308768 359872 308808
rect 436830 308796 436836 308808
rect 436888 308796 436894 308848
rect 439498 308768 439504 308780
rect 359844 308740 439504 308768
rect 439498 308728 439504 308740
rect 439556 308728 439562 308780
rect 348786 308700 348792 308712
rect 278056 308672 348792 308700
rect 348786 308660 348792 308672
rect 348844 308660 348850 308712
rect 352926 308660 352932 308712
rect 352984 308700 352990 308712
rect 438026 308700 438032 308712
rect 352984 308672 438032 308700
rect 352984 308660 352990 308672
rect 438026 308660 438032 308672
rect 438084 308660 438090 308712
rect 243596 308604 244274 308632
rect 243596 308592 243602 308604
rect 253750 308592 253756 308644
rect 253808 308632 253814 308644
rect 254394 308632 254400 308644
rect 253808 308604 254400 308632
rect 253808 308592 253814 308604
rect 254394 308592 254400 308604
rect 254452 308592 254458 308644
rect 256050 308592 256056 308644
rect 256108 308632 256114 308644
rect 262858 308632 262864 308644
rect 256108 308604 262864 308632
rect 256108 308592 256114 308604
rect 262858 308592 262864 308604
rect 262916 308592 262922 308644
rect 283926 308592 283932 308644
rect 283984 308632 283990 308644
rect 341058 308632 341064 308644
rect 283984 308604 341064 308632
rect 283984 308592 283990 308604
rect 341058 308592 341064 308604
rect 341116 308592 341122 308644
rect 353570 308592 353576 308644
rect 353628 308632 353634 308644
rect 439406 308632 439412 308644
rect 353628 308604 439412 308632
rect 353628 308592 353634 308604
rect 439406 308592 439412 308604
rect 439464 308592 439470 308644
rect 237156 308536 238754 308564
rect 237156 308524 237162 308536
rect 238938 308524 238944 308576
rect 238996 308564 239002 308576
rect 239582 308564 239588 308576
rect 238996 308536 239588 308564
rect 238996 308524 239002 308536
rect 239582 308524 239588 308536
rect 239640 308524 239646 308576
rect 253566 308524 253572 308576
rect 253624 308564 253630 308576
rect 262214 308564 262220 308576
rect 253624 308536 262220 308564
rect 253624 308524 253630 308536
rect 262214 308524 262220 308536
rect 262272 308524 262278 308576
rect 262490 308524 262496 308576
rect 262548 308564 262554 308576
rect 348142 308564 348148 308576
rect 262548 308536 348148 308564
rect 262548 308524 262554 308536
rect 348142 308524 348148 308536
rect 348200 308524 348206 308576
rect 352282 308524 352288 308576
rect 352340 308564 352346 308576
rect 440418 308564 440424 308576
rect 352340 308536 440424 308564
rect 352340 308524 352346 308536
rect 440418 308524 440424 308536
rect 440476 308524 440482 308576
rect 27672 308468 234614 308496
rect 27672 308456 27678 308468
rect 234706 308456 234712 308508
rect 234764 308496 234770 308508
rect 235902 308496 235908 308508
rect 234764 308468 235908 308496
rect 234764 308456 234770 308468
rect 235902 308456 235908 308468
rect 235960 308456 235966 308508
rect 238110 308456 238116 308508
rect 238168 308496 238174 308508
rect 350166 308496 350172 308508
rect 238168 308468 262720 308496
rect 238168 308456 238174 308468
rect 23474 308388 23480 308440
rect 23532 308428 23538 308440
rect 23532 308400 219434 308428
rect 23532 308388 23538 308400
rect 219406 308292 219434 308400
rect 234982 308388 234988 308440
rect 235040 308428 235046 308440
rect 235534 308428 235540 308440
rect 235040 308400 235540 308428
rect 235040 308388 235046 308400
rect 235534 308388 235540 308400
rect 235592 308388 235598 308440
rect 236086 308388 236092 308440
rect 236144 308428 236150 308440
rect 236638 308428 236644 308440
rect 236144 308400 236644 308428
rect 236144 308388 236150 308400
rect 236638 308388 236644 308400
rect 236696 308388 236702 308440
rect 237558 308388 237564 308440
rect 237616 308428 237622 308440
rect 237926 308428 237932 308440
rect 237616 308400 237932 308428
rect 237616 308388 237622 308400
rect 237926 308388 237932 308400
rect 237984 308388 237990 308440
rect 238754 308388 238760 308440
rect 238812 308428 238818 308440
rect 239122 308428 239128 308440
rect 238812 308400 239128 308428
rect 238812 308388 238818 308400
rect 239122 308388 239128 308400
rect 239180 308388 239186 308440
rect 240318 308388 240324 308440
rect 240376 308428 240382 308440
rect 240962 308428 240968 308440
rect 240376 308400 240968 308428
rect 240376 308388 240382 308400
rect 240962 308388 240968 308400
rect 241020 308388 241026 308440
rect 242894 308388 242900 308440
rect 242952 308428 242958 308440
rect 243446 308428 243452 308440
rect 242952 308400 243452 308428
rect 242952 308388 242958 308400
rect 243446 308388 243452 308400
rect 243504 308388 243510 308440
rect 247678 308388 247684 308440
rect 247736 308428 247742 308440
rect 258902 308428 258908 308440
rect 247736 308400 258908 308428
rect 247736 308388 247742 308400
rect 258902 308388 258908 308400
rect 258960 308388 258966 308440
rect 260190 308388 260196 308440
rect 260248 308428 260254 308440
rect 262582 308428 262588 308440
rect 260248 308400 262588 308428
rect 260248 308388 260254 308400
rect 262582 308388 262588 308400
rect 262640 308388 262646 308440
rect 262692 308428 262720 308468
rect 263566 308468 350172 308496
rect 263566 308428 263594 308468
rect 350166 308456 350172 308468
rect 350224 308456 350230 308508
rect 351638 308456 351644 308508
rect 351696 308496 351702 308508
rect 439590 308496 439596 308508
rect 351696 308468 439596 308496
rect 351696 308456 351702 308468
rect 439590 308456 439596 308468
rect 439648 308456 439654 308508
rect 262692 308400 263594 308428
rect 312078 308388 312084 308440
rect 312136 308428 312142 308440
rect 312998 308428 313004 308440
rect 312136 308400 313004 308428
rect 312136 308388 312142 308400
rect 312998 308388 313004 308400
rect 313056 308388 313062 308440
rect 313366 308388 313372 308440
rect 313424 308428 313430 308440
rect 313642 308428 313648 308440
rect 313424 308400 313648 308428
rect 313424 308388 313430 308400
rect 313642 308388 313648 308400
rect 313700 308388 313706 308440
rect 314654 308388 314660 308440
rect 314712 308428 314718 308440
rect 315666 308428 315672 308440
rect 314712 308400 315672 308428
rect 314712 308388 314718 308400
rect 315666 308388 315672 308400
rect 315724 308388 315730 308440
rect 315758 308388 315764 308440
rect 315816 308428 315822 308440
rect 437474 308428 437480 308440
rect 315816 308400 345704 308428
rect 315816 308388 315822 308400
rect 234798 308320 234804 308372
rect 234856 308360 234862 308372
rect 235442 308360 235448 308372
rect 234856 308332 235448 308360
rect 234856 308320 234862 308332
rect 235442 308320 235448 308332
rect 235500 308320 235506 308372
rect 237466 308320 237472 308372
rect 237524 308360 237530 308372
rect 238386 308360 238392 308372
rect 237524 308332 238392 308360
rect 237524 308320 237530 308332
rect 238386 308320 238392 308332
rect 238444 308320 238450 308372
rect 238846 308320 238852 308372
rect 238904 308360 238910 308372
rect 239398 308360 239404 308372
rect 238904 308332 239404 308360
rect 238904 308320 238910 308332
rect 239398 308320 239404 308332
rect 239456 308320 239462 308372
rect 242986 308320 242992 308372
rect 243044 308360 243050 308372
rect 243722 308360 243728 308372
rect 243044 308332 243728 308360
rect 243044 308320 243050 308332
rect 243722 308320 243728 308332
rect 243780 308320 243786 308372
rect 251910 308320 251916 308372
rect 251968 308360 251974 308372
rect 253750 308360 253756 308372
rect 251968 308332 253756 308360
rect 251968 308320 251974 308332
rect 253750 308320 253756 308332
rect 253808 308320 253814 308372
rect 262306 308320 262312 308372
rect 262364 308360 262370 308372
rect 263042 308360 263048 308372
rect 262364 308332 263048 308360
rect 262364 308320 262370 308332
rect 263042 308320 263048 308332
rect 263100 308320 263106 308372
rect 284202 308320 284208 308372
rect 284260 308360 284266 308372
rect 338390 308360 338396 308372
rect 284260 308332 338396 308360
rect 284260 308320 284266 308332
rect 338390 308320 338396 308332
rect 338448 308320 338454 308372
rect 234430 308292 234436 308304
rect 219406 308264 234436 308292
rect 234430 308252 234436 308264
rect 234488 308252 234494 308304
rect 237650 308252 237656 308304
rect 237708 308292 237714 308304
rect 238294 308292 238300 308304
rect 237708 308264 238300 308292
rect 237708 308252 237714 308264
rect 238294 308252 238300 308264
rect 238352 308252 238358 308304
rect 239214 308252 239220 308304
rect 239272 308292 239278 308304
rect 239674 308292 239680 308304
rect 239272 308264 239680 308292
rect 239272 308252 239278 308264
rect 239674 308252 239680 308264
rect 239732 308252 239738 308304
rect 241606 308252 241612 308304
rect 241664 308292 241670 308304
rect 242618 308292 242624 308304
rect 241664 308264 242624 308292
rect 241664 308252 241670 308264
rect 242618 308252 242624 308264
rect 242676 308252 242682 308304
rect 243078 308252 243084 308304
rect 243136 308292 243142 308304
rect 243814 308292 243820 308304
rect 243136 308264 243820 308292
rect 243136 308252 243142 308264
rect 243814 308252 243820 308264
rect 243872 308252 243878 308304
rect 274818 308252 274824 308304
rect 274876 308292 274882 308304
rect 276290 308292 276296 308304
rect 274876 308264 276296 308292
rect 274876 308252 274882 308264
rect 276290 308252 276296 308264
rect 276348 308252 276354 308304
rect 285490 308252 285496 308304
rect 285548 308292 285554 308304
rect 337286 308292 337292 308304
rect 285548 308264 337292 308292
rect 285548 308252 285554 308264
rect 337286 308252 337292 308264
rect 337344 308252 337350 308304
rect 345676 308292 345704 308400
rect 350368 308400 437480 308428
rect 350368 308292 350396 308400
rect 437474 308388 437480 308400
rect 437532 308388 437538 308440
rect 350718 308320 350724 308372
rect 350776 308360 350782 308372
rect 351822 308360 351828 308372
rect 350776 308332 351828 308360
rect 350776 308320 350782 308332
rect 351822 308320 351828 308332
rect 351880 308320 351886 308372
rect 352006 308320 352012 308372
rect 352064 308360 352070 308372
rect 352558 308360 352564 308372
rect 352064 308332 352564 308360
rect 352064 308320 352070 308332
rect 352558 308320 352564 308332
rect 352616 308320 352622 308372
rect 356054 308320 356060 308372
rect 356112 308360 356118 308372
rect 356606 308360 356612 308372
rect 356112 308332 356612 308360
rect 356112 308320 356118 308332
rect 356606 308320 356612 308332
rect 356664 308320 356670 308372
rect 358906 308320 358912 308372
rect 358964 308360 358970 308372
rect 359734 308360 359740 308372
rect 358964 308332 359740 308360
rect 358964 308320 358970 308332
rect 359734 308320 359740 308332
rect 359792 308320 359798 308372
rect 345676 308264 350396 308292
rect 350994 308252 351000 308304
rect 351052 308292 351058 308304
rect 351270 308292 351276 308304
rect 351052 308264 351276 308292
rect 351052 308252 351058 308264
rect 351270 308252 351276 308264
rect 351328 308252 351334 308304
rect 353662 308252 353668 308304
rect 353720 308292 353726 308304
rect 354306 308292 354312 308304
rect 353720 308264 354312 308292
rect 353720 308252 353726 308264
rect 354306 308252 354312 308264
rect 354364 308252 354370 308304
rect 355134 308252 355140 308304
rect 355192 308292 355198 308304
rect 355962 308292 355968 308304
rect 355192 308264 355968 308292
rect 355192 308252 355198 308264
rect 355962 308252 355968 308264
rect 356020 308252 356026 308304
rect 356146 308252 356152 308304
rect 356204 308292 356210 308304
rect 357250 308292 357256 308304
rect 356204 308264 357256 308292
rect 356204 308252 356210 308264
rect 357250 308252 357256 308264
rect 357308 308252 357314 308304
rect 357802 308252 357808 308304
rect 357860 308292 357866 308304
rect 358354 308292 358360 308304
rect 357860 308264 358360 308292
rect 357860 308252 357866 308264
rect 358354 308252 358360 308264
rect 358412 308252 358418 308304
rect 358998 308252 359004 308304
rect 359056 308292 359062 308304
rect 360102 308292 360108 308304
rect 359056 308264 360108 308292
rect 359056 308252 359062 308264
rect 360102 308252 360108 308264
rect 360160 308252 360166 308304
rect 238754 308184 238760 308236
rect 238812 308224 238818 308236
rect 240042 308224 240048 308236
rect 238812 308196 240048 308224
rect 238812 308184 238818 308196
rect 240042 308184 240048 308196
rect 240100 308184 240106 308236
rect 250990 308184 250996 308236
rect 251048 308224 251054 308236
rect 262490 308224 262496 308236
rect 251048 308196 262496 308224
rect 251048 308184 251054 308196
rect 262490 308184 262496 308196
rect 262548 308184 262554 308236
rect 337562 308224 337568 308236
rect 292546 308196 337568 308224
rect 234246 308116 234252 308168
rect 234304 308156 234310 308168
rect 243170 308156 243176 308168
rect 234304 308128 243176 308156
rect 234304 308116 234310 308128
rect 243170 308116 243176 308128
rect 243228 308116 243234 308168
rect 262858 308116 262864 308168
rect 262916 308156 262922 308168
rect 268378 308156 268384 308168
rect 262916 308128 268384 308156
rect 262916 308116 262922 308128
rect 268378 308116 268384 308128
rect 268436 308116 268442 308168
rect 242526 308048 242532 308100
rect 242584 308088 242590 308100
rect 249794 308088 249800 308100
rect 242584 308060 249800 308088
rect 242584 308048 242590 308060
rect 249794 308048 249800 308060
rect 249852 308048 249858 308100
rect 282638 308048 282644 308100
rect 282696 308088 282702 308100
rect 283558 308088 283564 308100
rect 282696 308060 283564 308088
rect 282696 308048 282702 308060
rect 283558 308048 283564 308060
rect 283616 308048 283622 308100
rect 243722 307980 243728 308032
rect 243780 308020 243786 308032
rect 249150 308020 249156 308032
rect 243780 307992 249156 308020
rect 243780 307980 243786 307992
rect 249150 307980 249156 307992
rect 249208 307980 249214 308032
rect 278774 307980 278780 308032
rect 278832 308020 278838 308032
rect 281258 308020 281264 308032
rect 278832 307992 281264 308020
rect 278832 307980 278838 307992
rect 281258 307980 281264 307992
rect 281316 307980 281322 308032
rect 244918 307912 244924 307964
rect 244976 307952 244982 307964
rect 250438 307952 250444 307964
rect 244976 307924 250444 307952
rect 244976 307912 244982 307924
rect 250438 307912 250444 307924
rect 250496 307912 250502 307964
rect 276658 307912 276664 307964
rect 276716 307952 276722 307964
rect 278866 307952 278872 307964
rect 276716 307924 278872 307952
rect 276716 307912 276722 307924
rect 278866 307912 278872 307924
rect 278924 307912 278930 307964
rect 291010 307912 291016 307964
rect 291068 307952 291074 307964
rect 292546 307952 292574 308196
rect 337562 308184 337568 308196
rect 337620 308184 337626 308236
rect 353386 308184 353392 308236
rect 353444 308224 353450 308236
rect 354030 308224 354036 308236
rect 353444 308196 354036 308224
rect 353444 308184 353450 308196
rect 354030 308184 354036 308196
rect 354088 308184 354094 308236
rect 312170 308116 312176 308168
rect 312228 308156 312234 308168
rect 312354 308156 312360 308168
rect 312228 308128 312360 308156
rect 312228 308116 312234 308128
rect 312354 308116 312360 308128
rect 312412 308116 312418 308168
rect 313550 308116 313556 308168
rect 313608 308156 313614 308168
rect 314286 308156 314292 308168
rect 313608 308128 314292 308156
rect 313608 308116 313614 308128
rect 314286 308116 314292 308128
rect 314344 308116 314350 308168
rect 314746 308116 314752 308168
rect 314804 308156 314810 308168
rect 314930 308156 314936 308168
rect 314804 308128 314936 308156
rect 314804 308116 314810 308128
rect 314930 308116 314936 308128
rect 314988 308116 314994 308168
rect 316310 308116 316316 308168
rect 316368 308156 316374 308168
rect 316862 308156 316868 308168
rect 316368 308128 316868 308156
rect 316368 308116 316374 308128
rect 316862 308116 316868 308128
rect 316920 308116 316926 308168
rect 317598 308116 317604 308168
rect 317656 308156 317662 308168
rect 317782 308156 317788 308168
rect 317656 308128 317788 308156
rect 317656 308116 317662 308128
rect 317782 308116 317788 308128
rect 317840 308116 317846 308168
rect 319070 308116 319076 308168
rect 319128 308156 319134 308168
rect 319714 308156 319720 308168
rect 319128 308128 319720 308156
rect 319128 308116 319134 308128
rect 319714 308116 319720 308128
rect 319772 308116 319778 308168
rect 320266 308116 320272 308168
rect 320324 308156 320330 308168
rect 321002 308156 321008 308168
rect 320324 308128 321008 308156
rect 320324 308116 320330 308128
rect 321002 308116 321008 308128
rect 321060 308116 321066 308168
rect 341058 308116 341064 308168
rect 341116 308156 341122 308168
rect 353846 308156 353852 308168
rect 341116 308128 353852 308156
rect 341116 308116 341122 308128
rect 353846 308116 353852 308128
rect 353904 308116 353910 308168
rect 356330 308116 356336 308168
rect 356388 308156 356394 308168
rect 357066 308156 357072 308168
rect 356388 308128 357072 308156
rect 356388 308116 356394 308128
rect 357066 308116 357072 308128
rect 357124 308116 357130 308168
rect 357618 308116 357624 308168
rect 357676 308156 357682 308168
rect 357986 308156 357992 308168
rect 357676 308128 357992 308156
rect 357676 308116 357682 308128
rect 357986 308116 357992 308128
rect 358044 308116 358050 308168
rect 358814 308116 358820 308168
rect 358872 308156 358878 308168
rect 359274 308156 359280 308168
rect 358872 308128 359280 308156
rect 358872 308116 358878 308128
rect 359274 308116 359280 308128
rect 359332 308116 359338 308168
rect 311894 308048 311900 308100
rect 311952 308088 311958 308100
rect 312538 308088 312544 308100
rect 311952 308060 312544 308088
rect 311952 308048 311958 308060
rect 312538 308048 312544 308060
rect 312596 308048 312602 308100
rect 313274 308048 313280 308100
rect 313332 308088 313338 308100
rect 314470 308088 314476 308100
rect 313332 308060 314476 308088
rect 313332 308048 313338 308060
rect 314470 308048 314476 308060
rect 314528 308048 314534 308100
rect 316218 308048 316224 308100
rect 316276 308088 316282 308100
rect 316954 308088 316960 308100
rect 316276 308060 316960 308088
rect 316276 308048 316282 308060
rect 316954 308048 316960 308060
rect 317012 308048 317018 308100
rect 317506 308048 317512 308100
rect 317564 308088 317570 308100
rect 318426 308088 318432 308100
rect 317564 308060 318432 308088
rect 317564 308048 317570 308060
rect 318426 308048 318432 308060
rect 318484 308048 318490 308100
rect 357526 308048 357532 308100
rect 357584 308088 357590 308100
rect 358446 308088 358452 308100
rect 357584 308060 358452 308088
rect 357584 308048 357590 308060
rect 358446 308048 358452 308060
rect 358504 308048 358510 308100
rect 359182 308048 359188 308100
rect 359240 308088 359246 308100
rect 359458 308088 359464 308100
rect 359240 308060 359464 308088
rect 359240 308048 359246 308060
rect 359458 308048 359464 308060
rect 359516 308048 359522 308100
rect 312170 307980 312176 308032
rect 312228 308020 312234 308032
rect 313182 308020 313188 308032
rect 312228 307992 313188 308020
rect 312228 307980 312234 307992
rect 313182 307980 313188 307992
rect 313240 307980 313246 308032
rect 314746 307980 314752 308032
rect 314804 308020 314810 308032
rect 315574 308020 315580 308032
rect 314804 307992 315580 308020
rect 314804 307980 314810 307992
rect 315574 307980 315580 307992
rect 315632 307980 315638 308032
rect 316126 307980 316132 308032
rect 316184 308020 316190 308032
rect 317322 308020 317328 308032
rect 316184 307992 317328 308020
rect 316184 307980 316190 307992
rect 317322 307980 317328 307992
rect 317380 307980 317386 308032
rect 317414 307980 317420 308032
rect 317472 308020 317478 308032
rect 318610 308020 318616 308032
rect 317472 307992 318616 308020
rect 317472 307980 317478 307992
rect 318610 307980 318616 307992
rect 318668 307980 318674 308032
rect 318794 307980 318800 308032
rect 318852 308020 318858 308032
rect 319254 308020 319260 308032
rect 318852 307992 319260 308020
rect 318852 307980 318858 307992
rect 319254 307980 319260 307992
rect 319312 307980 319318 308032
rect 354766 307980 354772 308032
rect 354824 308020 354830 308032
rect 355778 308020 355784 308032
rect 354824 307992 355784 308020
rect 354824 307980 354830 307992
rect 355778 307980 355784 307992
rect 355836 307980 355842 308032
rect 291068 307924 292574 307952
rect 291068 307912 291074 307924
rect 308030 307912 308036 307964
rect 308088 307952 308094 307964
rect 315758 307952 315764 307964
rect 308088 307924 315764 307952
rect 308088 307912 308094 307924
rect 315758 307912 315764 307924
rect 315816 307912 315822 307964
rect 358814 307912 358820 307964
rect 358872 307952 358878 307964
rect 359642 307952 359648 307964
rect 358872 307924 359648 307952
rect 358872 307912 358878 307924
rect 359642 307912 359648 307924
rect 359700 307912 359706 307964
rect 246482 307844 246488 307896
rect 246540 307884 246546 307896
rect 248966 307884 248972 307896
rect 246540 307856 248972 307884
rect 246540 307844 246546 307856
rect 248966 307844 248972 307856
rect 249024 307844 249030 307896
rect 278130 307844 278136 307896
rect 278188 307884 278194 307896
rect 279786 307884 279792 307896
rect 278188 307856 279792 307884
rect 278188 307844 278194 307856
rect 279786 307844 279792 307856
rect 279844 307844 279850 307896
rect 282822 307844 282828 307896
rect 282880 307884 282886 307896
rect 285122 307884 285128 307896
rect 282880 307856 285128 307884
rect 282880 307844 282886 307856
rect 285122 307844 285128 307856
rect 285180 307844 285186 307896
rect 286042 307844 286048 307896
rect 286100 307884 286106 307896
rect 291838 307884 291844 307896
rect 286100 307856 291844 307884
rect 286100 307844 286106 307856
rect 291838 307844 291844 307856
rect 291896 307844 291902 307896
rect 318794 307844 318800 307896
rect 318852 307884 318858 307896
rect 319898 307884 319904 307896
rect 318852 307856 319904 307884
rect 318852 307844 318858 307856
rect 319898 307844 319904 307856
rect 319956 307844 319962 307896
rect 236638 307776 236644 307828
rect 236696 307816 236702 307828
rect 237098 307816 237104 307828
rect 236696 307788 237104 307816
rect 236696 307776 236702 307788
rect 237098 307776 237104 307788
rect 237156 307776 237162 307828
rect 245010 307816 245016 307828
rect 242176 307788 245016 307816
rect 242176 307624 242204 307788
rect 245010 307776 245016 307788
rect 245068 307776 245074 307828
rect 246850 307776 246856 307828
rect 246908 307816 246914 307828
rect 248506 307816 248512 307828
rect 246908 307788 248512 307816
rect 246908 307776 246914 307788
rect 248506 307776 248512 307788
rect 248564 307776 248570 307828
rect 249058 307776 249064 307828
rect 249116 307816 249122 307828
rect 251358 307816 251364 307828
rect 249116 307788 251364 307816
rect 249116 307776 249122 307788
rect 251358 307776 251364 307788
rect 251416 307776 251422 307828
rect 257338 307776 257344 307828
rect 257396 307816 257402 307828
rect 258074 307816 258080 307828
rect 257396 307788 258080 307816
rect 257396 307776 257402 307788
rect 258074 307776 258080 307788
rect 258132 307776 258138 307828
rect 265618 307776 265624 307828
rect 265676 307816 265682 307828
rect 266722 307816 266728 307828
rect 265676 307788 266728 307816
rect 265676 307776 265682 307788
rect 266722 307776 266728 307788
rect 266780 307776 266786 307828
rect 271138 307776 271144 307828
rect 271196 307816 271202 307828
rect 271966 307816 271972 307828
rect 271196 307788 271972 307816
rect 271196 307776 271202 307788
rect 271966 307776 271972 307788
rect 272024 307776 272030 307828
rect 275370 307776 275376 307828
rect 275428 307816 275434 307828
rect 276750 307816 276756 307828
rect 275428 307788 276756 307816
rect 275428 307776 275434 307788
rect 276750 307776 276756 307788
rect 276808 307776 276814 307828
rect 277118 307776 277124 307828
rect 277176 307816 277182 307828
rect 278038 307816 278044 307828
rect 277176 307788 278044 307816
rect 277176 307776 277182 307788
rect 278038 307776 278044 307788
rect 278096 307776 278102 307828
rect 279510 307776 279516 307828
rect 279568 307816 279574 307828
rect 281074 307816 281080 307828
rect 279568 307788 281080 307816
rect 279568 307776 279574 307788
rect 281074 307776 281080 307788
rect 281132 307776 281138 307828
rect 284110 307776 284116 307828
rect 284168 307816 284174 307828
rect 284938 307816 284944 307828
rect 284168 307788 284944 307816
rect 284168 307776 284174 307788
rect 284938 307776 284944 307788
rect 284996 307776 285002 307828
rect 285030 307776 285036 307828
rect 285088 307816 285094 307828
rect 286318 307816 286324 307828
rect 285088 307788 286324 307816
rect 285088 307776 285094 307788
rect 286318 307776 286324 307788
rect 286376 307776 286382 307828
rect 293218 307776 293224 307828
rect 293276 307816 293282 307828
rect 294690 307816 294696 307828
rect 293276 307788 294696 307816
rect 293276 307776 293282 307788
rect 294690 307776 294696 307788
rect 294748 307776 294754 307828
rect 295150 307776 295156 307828
rect 295208 307816 295214 307828
rect 296438 307816 296444 307828
rect 295208 307788 296444 307816
rect 295208 307776 295214 307788
rect 296438 307776 296444 307788
rect 296496 307776 296502 307828
rect 328638 307708 328644 307760
rect 328696 307748 328702 307760
rect 329374 307748 329380 307760
rect 328696 307720 329380 307748
rect 328696 307708 328702 307720
rect 329374 307708 329380 307720
rect 329432 307708 329438 307760
rect 243262 307640 243268 307692
rect 243320 307680 243326 307692
rect 244182 307680 244188 307692
rect 243320 307652 244188 307680
rect 243320 307640 243326 307652
rect 244182 307640 244188 307652
rect 244240 307640 244246 307692
rect 320358 307640 320364 307692
rect 320416 307680 320422 307692
rect 320542 307680 320548 307692
rect 320416 307652 320548 307680
rect 320416 307640 320422 307652
rect 320542 307640 320548 307652
rect 320600 307640 320606 307692
rect 242158 307572 242164 307624
rect 242216 307572 242222 307624
rect 320542 307504 320548 307556
rect 320600 307544 320606 307556
rect 321462 307544 321468 307556
rect 320600 307516 321468 307544
rect 320600 307504 320606 307516
rect 321462 307504 321468 307516
rect 321520 307504 321526 307556
rect 326706 307232 326712 307284
rect 326764 307272 326770 307284
rect 445018 307272 445024 307284
rect 326764 307244 445024 307272
rect 326764 307232 326770 307244
rect 445018 307232 445024 307244
rect 445076 307232 445082 307284
rect 80054 307164 80060 307216
rect 80112 307204 80118 307216
rect 244826 307204 244832 307216
rect 80112 307176 244832 307204
rect 80112 307164 80118 307176
rect 244826 307164 244832 307176
rect 244884 307164 244890 307216
rect 316494 307164 316500 307216
rect 316552 307204 316558 307216
rect 467098 307204 467104 307216
rect 316552 307176 467104 307204
rect 316552 307164 316558 307176
rect 467098 307164 467104 307176
rect 467156 307164 467162 307216
rect 57974 307096 57980 307148
rect 58032 307136 58038 307148
rect 240686 307136 240692 307148
rect 58032 307108 240692 307136
rect 58032 307096 58038 307108
rect 240686 307096 240692 307108
rect 240744 307096 240750 307148
rect 318242 307096 318248 307148
rect 318300 307136 318306 307148
rect 476758 307136 476764 307148
rect 318300 307108 476764 307136
rect 318300 307096 318306 307108
rect 476758 307096 476764 307108
rect 476816 307096 476822 307148
rect 25498 307028 25504 307080
rect 25556 307068 25562 307080
rect 230106 307068 230112 307080
rect 25556 307040 230112 307068
rect 25556 307028 25562 307040
rect 230106 307028 230112 307040
rect 230164 307028 230170 307080
rect 251174 307028 251180 307080
rect 251232 307068 251238 307080
rect 274818 307068 274824 307080
rect 251232 307040 274824 307068
rect 251232 307028 251238 307040
rect 274818 307028 274824 307040
rect 274876 307028 274882 307080
rect 284294 307028 284300 307080
rect 284352 307068 284358 307080
rect 293218 307068 293224 307080
rect 284352 307040 293224 307068
rect 284352 307028 284358 307040
rect 293218 307028 293224 307040
rect 293276 307028 293282 307080
rect 322106 307028 322112 307080
rect 322164 307068 322170 307080
rect 500218 307068 500224 307080
rect 322164 307040 500224 307068
rect 322164 307028 322170 307040
rect 500218 307028 500224 307040
rect 500276 307028 500282 307080
rect 272150 306960 272156 307012
rect 272208 306960 272214 307012
rect 288894 306960 288900 307012
rect 288952 306960 288958 307012
rect 245838 306824 245844 306876
rect 245896 306824 245902 306876
rect 245856 306604 245884 306824
rect 266354 306756 266360 306808
rect 266412 306796 266418 306808
rect 266630 306796 266636 306808
rect 266412 306768 266636 306796
rect 266412 306756 266418 306768
rect 266630 306756 266636 306768
rect 266688 306756 266694 306808
rect 272058 306756 272064 306808
rect 272116 306796 272122 306808
rect 272168 306796 272196 306960
rect 272116 306768 272196 306796
rect 288912 306796 288940 306960
rect 288986 306796 288992 306808
rect 288912 306768 288992 306796
rect 272116 306756 272122 306768
rect 288986 306756 288992 306768
rect 289044 306756 289050 306808
rect 299474 306688 299480 306740
rect 299532 306728 299538 306740
rect 299934 306728 299940 306740
rect 299532 306700 299940 306728
rect 299532 306688 299538 306700
rect 299934 306688 299940 306700
rect 299992 306688 299998 306740
rect 320174 306688 320180 306740
rect 320232 306728 320238 306740
rect 320726 306728 320732 306740
rect 320232 306700 320732 306728
rect 320232 306688 320238 306700
rect 320726 306688 320732 306700
rect 320784 306688 320790 306740
rect 329834 306688 329840 306740
rect 329892 306728 329898 306740
rect 330202 306728 330208 306740
rect 329892 306700 330208 306728
rect 329892 306688 329898 306700
rect 330202 306688 330208 306700
rect 330260 306688 330266 306740
rect 335814 306688 335820 306740
rect 335872 306728 335878 306740
rect 336090 306728 336096 306740
rect 335872 306700 336096 306728
rect 335872 306688 335878 306700
rect 336090 306688 336096 306700
rect 336148 306688 336154 306740
rect 273438 306620 273444 306672
rect 273496 306660 273502 306672
rect 273622 306660 273628 306672
rect 273496 306632 273628 306660
rect 273496 306620 273502 306632
rect 273622 306620 273628 306632
rect 273680 306620 273686 306672
rect 322934 306620 322940 306672
rect 322992 306660 322998 306672
rect 323486 306660 323492 306672
rect 322992 306632 323492 306660
rect 322992 306620 322998 306632
rect 323486 306620 323492 306632
rect 323544 306620 323550 306672
rect 230934 306552 230940 306604
rect 230992 306552 230998 306604
rect 245838 306552 245844 306604
rect 245896 306552 245902 306604
rect 263870 306552 263876 306604
rect 263928 306552 263934 306604
rect 283006 306552 283012 306604
rect 283064 306552 283070 306604
rect 291654 306552 291660 306604
rect 291712 306552 291718 306604
rect 320174 306552 320180 306604
rect 320232 306592 320238 306604
rect 321094 306592 321100 306604
rect 320232 306564 321100 306592
rect 320232 306552 320238 306564
rect 321094 306552 321100 306564
rect 321152 306552 321158 306604
rect 323210 306552 323216 306604
rect 323268 306552 323274 306604
rect 343634 306552 343640 306604
rect 343692 306592 343698 306604
rect 344002 306592 344008 306604
rect 343692 306564 344008 306592
rect 343692 306552 343698 306564
rect 344002 306552 344008 306564
rect 344060 306552 344066 306604
rect 230952 306400 230980 306552
rect 245930 306484 245936 306536
rect 245988 306524 245994 306536
rect 246390 306524 246396 306536
rect 245988 306496 246396 306524
rect 245988 306484 245994 306496
rect 246390 306484 246396 306496
rect 246448 306484 246454 306536
rect 250070 306484 250076 306536
rect 250128 306524 250134 306536
rect 250530 306524 250536 306536
rect 250128 306496 250536 306524
rect 250128 306484 250134 306496
rect 250530 306484 250536 306496
rect 250588 306484 250594 306536
rect 241514 306416 241520 306468
rect 241572 306456 241578 306468
rect 241790 306456 241796 306468
rect 241572 306428 241796 306456
rect 241572 306416 241578 306428
rect 241790 306416 241796 306428
rect 241848 306416 241854 306468
rect 245746 306416 245752 306468
rect 245804 306456 245810 306468
rect 246298 306456 246304 306468
rect 245804 306428 246304 306456
rect 245804 306416 245810 306428
rect 246298 306416 246304 306428
rect 246356 306416 246362 306468
rect 247310 306416 247316 306468
rect 247368 306456 247374 306468
rect 248138 306456 248144 306468
rect 247368 306428 248144 306456
rect 247368 306416 247374 306428
rect 248138 306416 248144 306428
rect 248196 306416 248202 306468
rect 249886 306416 249892 306468
rect 249944 306456 249950 306468
rect 250254 306456 250260 306468
rect 249944 306428 250260 306456
rect 249944 306416 249950 306428
rect 250254 306416 250260 306428
rect 250312 306416 250318 306468
rect 256970 306416 256976 306468
rect 257028 306456 257034 306468
rect 257154 306456 257160 306468
rect 257028 306428 257160 306456
rect 257028 306416 257034 306428
rect 257154 306416 257160 306428
rect 257212 306416 257218 306468
rect 260834 306416 260840 306468
rect 260892 306456 260898 306468
rect 261294 306456 261300 306468
rect 260892 306428 261300 306456
rect 260892 306416 260898 306428
rect 261294 306416 261300 306428
rect 261352 306416 261358 306468
rect 263888 306400 263916 306552
rect 270678 306416 270684 306468
rect 270736 306456 270742 306468
rect 270954 306456 270960 306468
rect 270736 306428 270960 306456
rect 270736 306416 270742 306428
rect 270954 306416 270960 306428
rect 271012 306416 271018 306468
rect 277578 306416 277584 306468
rect 277636 306456 277642 306468
rect 278222 306456 278228 306468
rect 277636 306428 278228 306456
rect 277636 306416 277642 306428
rect 278222 306416 278228 306428
rect 278280 306416 278286 306468
rect 281534 306416 281540 306468
rect 281592 306456 281598 306468
rect 281902 306456 281908 306468
rect 281592 306428 281908 306456
rect 281592 306416 281598 306428
rect 281902 306416 281908 306428
rect 281960 306416 281966 306468
rect 230934 306348 230940 306400
rect 230992 306348 230998 306400
rect 232038 306348 232044 306400
rect 232096 306388 232102 306400
rect 232958 306388 232964 306400
rect 232096 306360 232964 306388
rect 232096 306348 232102 306360
rect 232958 306348 232964 306360
rect 233016 306348 233022 306400
rect 247402 306348 247408 306400
rect 247460 306388 247466 306400
rect 248046 306388 248052 306400
rect 247460 306360 248052 306388
rect 247460 306348 247466 306360
rect 248046 306348 248052 306360
rect 248104 306348 248110 306400
rect 248506 306348 248512 306400
rect 248564 306388 248570 306400
rect 249242 306388 249248 306400
rect 248564 306360 249248 306388
rect 248564 306348 248570 306360
rect 249242 306348 249248 306360
rect 249300 306348 249306 306400
rect 252646 306348 252652 306400
rect 252704 306388 252710 306400
rect 253290 306388 253296 306400
rect 252704 306360 253296 306388
rect 252704 306348 252710 306360
rect 253290 306348 253296 306360
rect 253348 306348 253354 306400
rect 255406 306348 255412 306400
rect 255464 306388 255470 306400
rect 256510 306388 256516 306400
rect 255464 306360 256516 306388
rect 255464 306348 255470 306360
rect 256510 306348 256516 306360
rect 256568 306348 256574 306400
rect 256878 306348 256884 306400
rect 256936 306388 256942 306400
rect 257706 306388 257712 306400
rect 256936 306360 257712 306388
rect 256936 306348 256942 306360
rect 257706 306348 257712 306360
rect 257764 306348 257770 306400
rect 258258 306348 258264 306400
rect 258316 306388 258322 306400
rect 258994 306388 259000 306400
rect 258316 306360 259000 306388
rect 258316 306348 258322 306360
rect 258994 306348 259000 306360
rect 259052 306348 259058 306400
rect 259638 306348 259644 306400
rect 259696 306388 259702 306400
rect 260006 306388 260012 306400
rect 259696 306360 260012 306388
rect 259696 306348 259702 306360
rect 260006 306348 260012 306360
rect 260064 306348 260070 306400
rect 263870 306348 263876 306400
rect 263928 306348 263934 306400
rect 265342 306348 265348 306400
rect 265400 306388 265406 306400
rect 266078 306388 266084 306400
rect 265400 306360 266084 306388
rect 265400 306348 265406 306360
rect 266078 306348 266084 306360
rect 266136 306348 266142 306400
rect 268102 306348 268108 306400
rect 268160 306388 268166 306400
rect 268562 306388 268568 306400
rect 268160 306360 268568 306388
rect 268160 306348 268166 306360
rect 268562 306348 268568 306360
rect 268620 306348 268626 306400
rect 270494 306348 270500 306400
rect 270552 306388 270558 306400
rect 271598 306388 271604 306400
rect 270552 306360 271604 306388
rect 270552 306348 270558 306360
rect 271598 306348 271604 306360
rect 271656 306348 271662 306400
rect 273346 306348 273352 306400
rect 273404 306388 273410 306400
rect 274358 306388 274364 306400
rect 273404 306360 274364 306388
rect 273404 306348 273410 306360
rect 274358 306348 274364 306360
rect 274416 306348 274422 306400
rect 278958 306348 278964 306400
rect 279016 306388 279022 306400
rect 279326 306388 279332 306400
rect 279016 306360 279332 306388
rect 279016 306348 279022 306360
rect 279326 306348 279332 306360
rect 279384 306348 279390 306400
rect 283024 306332 283052 306552
rect 289814 306416 289820 306468
rect 289872 306456 289878 306468
rect 290642 306456 290648 306468
rect 289872 306428 290648 306456
rect 289872 306416 289878 306428
rect 290642 306416 290648 306428
rect 290700 306416 290706 306468
rect 284386 306348 284392 306400
rect 284444 306388 284450 306400
rect 285214 306388 285220 306400
rect 284444 306360 285220 306388
rect 284444 306348 284450 306360
rect 285214 306348 285220 306360
rect 285272 306348 285278 306400
rect 287238 306348 287244 306400
rect 287296 306388 287302 306400
rect 287790 306388 287796 306400
rect 287296 306360 287796 306388
rect 287296 306348 287302 306360
rect 287790 306348 287796 306360
rect 287848 306348 287854 306400
rect 288618 306348 288624 306400
rect 288676 306388 288682 306400
rect 289722 306388 289728 306400
rect 288676 306360 289728 306388
rect 288676 306348 288682 306360
rect 289722 306348 289728 306360
rect 289780 306348 289786 306400
rect 290090 306348 290096 306400
rect 290148 306388 290154 306400
rect 290826 306388 290832 306400
rect 290148 306360 290832 306388
rect 290148 306348 290154 306360
rect 290826 306348 290832 306360
rect 290884 306348 290890 306400
rect 291672 306332 291700 306552
rect 295610 306484 295616 306536
rect 295668 306524 295674 306536
rect 296346 306524 296352 306536
rect 295668 306496 296352 306524
rect 295668 306484 295674 306496
rect 296346 306484 296352 306496
rect 296404 306484 296410 306536
rect 307754 306484 307760 306536
rect 307812 306524 307818 306536
rect 308398 306524 308404 306536
rect 307812 306496 308404 306524
rect 307812 306484 307818 306496
rect 308398 306484 308404 306496
rect 308456 306484 308462 306536
rect 295426 306416 295432 306468
rect 295484 306456 295490 306468
rect 296070 306456 296076 306468
rect 295484 306428 296076 306456
rect 295484 306416 295490 306428
rect 296070 306416 296076 306428
rect 296128 306416 296134 306468
rect 302234 306416 302240 306468
rect 302292 306456 302298 306468
rect 302510 306456 302516 306468
rect 302292 306428 302516 306456
rect 302292 306416 302298 306428
rect 302510 306416 302516 306428
rect 302568 306416 302574 306468
rect 308030 306416 308036 306468
rect 308088 306456 308094 306468
rect 308490 306456 308496 306468
rect 308088 306428 308496 306456
rect 308088 306416 308094 306428
rect 308490 306416 308496 306428
rect 308548 306416 308554 306468
rect 310514 306416 310520 306468
rect 310572 306456 310578 306468
rect 311250 306456 311256 306468
rect 310572 306428 311256 306456
rect 310572 306416 310578 306428
rect 311250 306416 311256 306428
rect 311308 306416 311314 306468
rect 295702 306348 295708 306400
rect 295760 306388 295766 306400
rect 296254 306388 296260 306400
rect 295760 306360 296260 306388
rect 295760 306348 295766 306360
rect 296254 306348 296260 306360
rect 296312 306348 296318 306400
rect 298278 306348 298284 306400
rect 298336 306388 298342 306400
rect 299290 306388 299296 306400
rect 298336 306360 299296 306388
rect 298336 306348 298342 306360
rect 299290 306348 299296 306360
rect 299348 306348 299354 306400
rect 301038 306348 301044 306400
rect 301096 306388 301102 306400
rect 302142 306388 302148 306400
rect 301096 306360 302148 306388
rect 301096 306348 301102 306360
rect 302142 306348 302148 306360
rect 302200 306348 302206 306400
rect 306650 306348 306656 306400
rect 306708 306388 306714 306400
rect 307110 306388 307116 306400
rect 306708 306360 307116 306388
rect 306708 306348 306714 306360
rect 307110 306348 307116 306360
rect 307168 306348 307174 306400
rect 308122 306348 308128 306400
rect 308180 306388 308186 306400
rect 308858 306388 308864 306400
rect 308180 306360 308864 306388
rect 308180 306348 308186 306360
rect 308858 306348 308864 306360
rect 308916 306348 308922 306400
rect 309318 306348 309324 306400
rect 309376 306388 309382 306400
rect 309962 306388 309968 306400
rect 309376 306360 309968 306388
rect 309376 306348 309382 306360
rect 309962 306348 309968 306360
rect 310020 306348 310026 306400
rect 310698 306348 310704 306400
rect 310756 306388 310762 306400
rect 311434 306388 311440 306400
rect 310756 306360 311440 306388
rect 310756 306348 310762 306360
rect 311434 306348 311440 306360
rect 311492 306348 311498 306400
rect 323118 306348 323124 306400
rect 323176 306388 323182 306400
rect 323228 306388 323256 306552
rect 325786 306484 325792 306536
rect 325844 306524 325850 306536
rect 326890 306524 326896 306536
rect 325844 306496 326896 306524
rect 325844 306484 325850 306496
rect 326890 306484 326896 306496
rect 326948 306484 326954 306536
rect 327350 306484 327356 306536
rect 327408 306524 327414 306536
rect 327902 306524 327908 306536
rect 327408 306496 327908 306524
rect 327408 306484 327414 306496
rect 327902 306484 327908 306496
rect 327960 306484 327966 306536
rect 328362 306484 328368 306536
rect 328420 306524 328426 306536
rect 328914 306524 328920 306536
rect 328420 306496 328920 306524
rect 328420 306484 328426 306496
rect 328914 306484 328920 306496
rect 328972 306484 328978 306536
rect 325694 306416 325700 306468
rect 325752 306456 325758 306468
rect 326430 306456 326436 306468
rect 325752 306428 326436 306456
rect 325752 306416 325758 306428
rect 326430 306416 326436 306428
rect 326488 306416 326494 306468
rect 327074 306416 327080 306468
rect 327132 306456 327138 306468
rect 328178 306456 328184 306468
rect 327132 306428 328184 306456
rect 327132 306416 327138 306428
rect 328178 306416 328184 306428
rect 328236 306416 328242 306468
rect 331306 306416 331312 306468
rect 331364 306456 331370 306468
rect 331674 306456 331680 306468
rect 331364 306428 331680 306456
rect 331364 306416 331370 306428
rect 331674 306416 331680 306428
rect 331732 306416 331738 306468
rect 334066 306416 334072 306468
rect 334124 306456 334130 306468
rect 334342 306456 334348 306468
rect 334124 306428 334348 306456
rect 334124 306416 334130 306428
rect 334342 306416 334348 306428
rect 334400 306416 334406 306468
rect 323176 306360 323256 306388
rect 323176 306348 323182 306360
rect 323302 306348 323308 306400
rect 323360 306388 323366 306400
rect 324038 306388 324044 306400
rect 323360 306360 324044 306388
rect 323360 306348 323366 306360
rect 324038 306348 324044 306360
rect 324096 306348 324102 306400
rect 324314 306348 324320 306400
rect 324372 306388 324378 306400
rect 324590 306388 324596 306400
rect 324372 306360 324596 306388
rect 324372 306348 324378 306360
rect 324590 306348 324596 306360
rect 324648 306348 324654 306400
rect 325878 306348 325884 306400
rect 325936 306388 325942 306400
rect 326246 306388 326252 306400
rect 325936 306360 326252 306388
rect 325936 306348 325942 306360
rect 326246 306348 326252 306360
rect 326304 306348 326310 306400
rect 327258 306348 327264 306400
rect 327316 306388 327322 306400
rect 327718 306388 327724 306400
rect 327316 306360 327724 306388
rect 327316 306348 327322 306360
rect 327718 306348 327724 306360
rect 327776 306348 327782 306400
rect 328426 306360 331352 306388
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 221458 306320 221464 306332
rect 3384 306292 221464 306320
rect 3384 306280 3390 306292
rect 221458 306280 221464 306292
rect 221516 306280 221522 306332
rect 230658 306280 230664 306332
rect 230716 306320 230722 306332
rect 231578 306320 231584 306332
rect 230716 306292 231584 306320
rect 230716 306280 230722 306292
rect 231578 306280 231584 306292
rect 231636 306280 231642 306332
rect 231946 306280 231952 306332
rect 232004 306320 232010 306332
rect 232498 306320 232504 306332
rect 232004 306292 232504 306320
rect 232004 306280 232010 306292
rect 232498 306280 232504 306292
rect 232556 306280 232562 306332
rect 244458 306280 244464 306332
rect 244516 306320 244522 306332
rect 245470 306320 245476 306332
rect 244516 306292 245476 306320
rect 244516 306280 244522 306292
rect 245470 306280 245476 306292
rect 245528 306280 245534 306332
rect 247034 306280 247040 306332
rect 247092 306320 247098 306332
rect 247586 306320 247592 306332
rect 247092 306292 247592 306320
rect 247092 306280 247098 306292
rect 247586 306280 247592 306292
rect 247644 306280 247650 306332
rect 248598 306280 248604 306332
rect 248656 306320 248662 306332
rect 249610 306320 249616 306332
rect 248656 306292 249616 306320
rect 248656 306280 248662 306292
rect 249610 306280 249616 306292
rect 249668 306280 249674 306332
rect 252830 306280 252836 306332
rect 252888 306320 252894 306332
rect 253014 306320 253020 306332
rect 252888 306292 253020 306320
rect 252888 306280 252894 306292
rect 253014 306280 253020 306292
rect 253072 306280 253078 306332
rect 253934 306280 253940 306332
rect 253992 306320 253998 306332
rect 254210 306320 254216 306332
rect 253992 306292 254216 306320
rect 253992 306280 253998 306292
rect 254210 306280 254216 306292
rect 254268 306280 254274 306332
rect 254302 306280 254308 306332
rect 254360 306320 254366 306332
rect 255038 306320 255044 306332
rect 254360 306292 255044 306320
rect 254360 306280 254366 306292
rect 255038 306280 255044 306292
rect 255096 306280 255102 306332
rect 255314 306280 255320 306332
rect 255372 306320 255378 306332
rect 255958 306320 255964 306332
rect 255372 306292 255964 306320
rect 255372 306280 255378 306292
rect 255958 306280 255964 306292
rect 256016 306280 256022 306332
rect 256786 306280 256792 306332
rect 256844 306320 256850 306332
rect 257246 306320 257252 306332
rect 256844 306292 257252 306320
rect 256844 306280 256850 306292
rect 257246 306280 257252 306292
rect 257304 306280 257310 306332
rect 258166 306280 258172 306332
rect 258224 306320 258230 306332
rect 258718 306320 258724 306332
rect 258224 306292 258724 306320
rect 258224 306280 258230 306292
rect 258718 306280 258724 306292
rect 258776 306280 258782 306332
rect 259454 306280 259460 306332
rect 259512 306320 259518 306332
rect 260098 306320 260104 306332
rect 259512 306292 260104 306320
rect 259512 306280 259518 306292
rect 260098 306280 260104 306292
rect 260156 306280 260162 306332
rect 261018 306280 261024 306332
rect 261076 306320 261082 306332
rect 261754 306320 261760 306332
rect 261076 306292 261760 306320
rect 261076 306280 261082 306292
rect 261754 306280 261760 306292
rect 261812 306280 261818 306332
rect 262490 306280 262496 306332
rect 262548 306320 262554 306332
rect 263502 306320 263508 306332
rect 262548 306292 263508 306320
rect 262548 306280 262554 306292
rect 263502 306280 263508 306292
rect 263560 306280 263566 306332
rect 263594 306280 263600 306332
rect 263652 306320 263658 306332
rect 264422 306320 264428 306332
rect 263652 306292 264428 306320
rect 263652 306280 263658 306292
rect 264422 306280 264428 306292
rect 264480 306280 264486 306332
rect 265250 306280 265256 306332
rect 265308 306320 265314 306332
rect 265526 306320 265532 306332
rect 265308 306292 265532 306320
rect 265308 306280 265314 306292
rect 265526 306280 265532 306292
rect 265584 306280 265590 306332
rect 268010 306280 268016 306332
rect 268068 306320 268074 306332
rect 268286 306320 268292 306332
rect 268068 306292 268292 306320
rect 268068 306280 268074 306292
rect 268286 306280 268292 306292
rect 268344 306280 268350 306332
rect 269206 306280 269212 306332
rect 269264 306320 269270 306332
rect 270402 306320 270408 306332
rect 269264 306292 270408 306320
rect 269264 306280 269270 306292
rect 270402 306280 270408 306292
rect 270460 306280 270466 306332
rect 270586 306280 270592 306332
rect 270644 306320 270650 306332
rect 271506 306320 271512 306332
rect 270644 306292 271512 306320
rect 270644 306280 270650 306292
rect 271506 306280 271512 306292
rect 271564 306280 271570 306332
rect 273530 306280 273536 306332
rect 273588 306320 273594 306332
rect 274542 306320 274548 306332
rect 273588 306292 274548 306320
rect 273588 306280 273594 306292
rect 274542 306280 274548 306292
rect 274600 306280 274606 306332
rect 274910 306280 274916 306332
rect 274968 306320 274974 306332
rect 275830 306320 275836 306332
rect 274968 306292 275836 306320
rect 274968 306280 274974 306292
rect 275830 306280 275836 306292
rect 275888 306280 275894 306332
rect 277762 306280 277768 306332
rect 277820 306320 277826 306332
rect 278314 306320 278320 306332
rect 277820 306292 278320 306320
rect 277820 306280 277826 306292
rect 278314 306280 278320 306292
rect 278372 306280 278378 306332
rect 278866 306280 278872 306332
rect 278924 306320 278930 306332
rect 279970 306320 279976 306332
rect 278924 306292 279976 306320
rect 278924 306280 278930 306292
rect 279970 306280 279976 306292
rect 280028 306280 280034 306332
rect 283006 306280 283012 306332
rect 283064 306280 283070 306332
rect 283650 306320 283656 306332
rect 283116 306292 283656 306320
rect 283116 306264 283144 306292
rect 283650 306280 283656 306292
rect 283708 306280 283714 306332
rect 284294 306280 284300 306332
rect 284352 306320 284358 306332
rect 284754 306320 284760 306332
rect 284352 306292 284760 306320
rect 284352 306280 284358 306292
rect 284754 306280 284760 306292
rect 284812 306280 284818 306332
rect 287146 306280 287152 306332
rect 287204 306320 287210 306332
rect 287422 306320 287428 306332
rect 287204 306292 287428 306320
rect 287204 306280 287210 306292
rect 287422 306280 287428 306292
rect 287480 306280 287486 306332
rect 288434 306280 288440 306332
rect 288492 306320 288498 306332
rect 288802 306320 288808 306332
rect 288492 306292 288808 306320
rect 288492 306280 288498 306292
rect 288802 306280 288808 306292
rect 288860 306280 288866 306332
rect 289998 306280 290004 306332
rect 290056 306320 290062 306332
rect 290918 306320 290924 306332
rect 290056 306292 290924 306320
rect 290056 306280 290062 306292
rect 290918 306280 290924 306292
rect 290976 306280 290982 306332
rect 291654 306280 291660 306332
rect 291712 306280 291718 306332
rect 292666 306280 292672 306332
rect 292724 306320 292730 306332
rect 293678 306320 293684 306332
rect 292724 306292 293684 306320
rect 292724 306280 292730 306292
rect 293678 306280 293684 306292
rect 293736 306280 293742 306332
rect 293954 306280 293960 306332
rect 294012 306320 294018 306332
rect 294598 306320 294604 306332
rect 294012 306292 294604 306320
rect 294012 306280 294018 306292
rect 294598 306280 294604 306292
rect 294656 306280 294662 306332
rect 295518 306280 295524 306332
rect 295576 306320 295582 306332
rect 295886 306320 295892 306332
rect 295576 306292 295892 306320
rect 295576 306280 295582 306292
rect 295886 306280 295892 306292
rect 295944 306280 295950 306332
rect 298186 306280 298192 306332
rect 298244 306320 298250 306332
rect 298646 306320 298652 306332
rect 298244 306292 298652 306320
rect 298244 306280 298250 306292
rect 298646 306280 298652 306292
rect 298704 306280 298710 306332
rect 299842 306280 299848 306332
rect 299900 306320 299906 306332
rect 300394 306320 300400 306332
rect 299900 306292 300400 306320
rect 299900 306280 299906 306292
rect 300394 306280 300400 306292
rect 300452 306280 300458 306332
rect 300946 306280 300952 306332
rect 301004 306320 301010 306332
rect 301498 306320 301504 306332
rect 301004 306292 301504 306320
rect 301004 306280 301010 306292
rect 301498 306280 301504 306292
rect 301556 306280 301562 306332
rect 301590 306280 301596 306332
rect 301648 306320 301654 306332
rect 328426 306320 328454 306360
rect 301648 306292 328454 306320
rect 331324 306320 331352 306360
rect 331582 306348 331588 306400
rect 331640 306388 331646 306400
rect 332502 306388 332508 306400
rect 331640 306360 332508 306388
rect 331640 306348 331646 306360
rect 332502 306348 332508 306360
rect 332560 306348 332566 306400
rect 333974 306348 333980 306400
rect 334032 306388 334038 306400
rect 334894 306388 334900 306400
rect 334032 306360 334900 306388
rect 334032 306348 334038 306360
rect 334894 306348 334900 306360
rect 334952 306348 334958 306400
rect 338298 306348 338304 306400
rect 338356 306388 338362 306400
rect 339126 306388 339132 306400
rect 338356 306360 339132 306388
rect 338356 306348 338362 306360
rect 339126 306348 339132 306360
rect 339184 306348 339190 306400
rect 341150 306348 341156 306400
rect 341208 306388 341214 306400
rect 341610 306388 341616 306400
rect 341208 306360 341616 306388
rect 341208 306348 341214 306360
rect 341610 306348 341616 306360
rect 341668 306348 341674 306400
rect 345198 306348 345204 306400
rect 345256 306388 345262 306400
rect 345750 306388 345756 306400
rect 345256 306360 345756 306388
rect 345256 306348 345262 306360
rect 345750 306348 345756 306360
rect 345808 306348 345814 306400
rect 331324 306292 340874 306320
rect 301648 306280 301654 306292
rect 230750 306212 230756 306264
rect 230808 306252 230814 306264
rect 231026 306252 231032 306264
rect 230808 306224 231032 306252
rect 230808 306212 230814 306224
rect 231026 306212 231032 306224
rect 231084 306212 231090 306264
rect 246114 306212 246120 306264
rect 246172 306252 246178 306264
rect 246758 306252 246764 306264
rect 246172 306224 246764 306252
rect 246172 306212 246178 306224
rect 246758 306212 246764 306224
rect 246816 306212 246822 306264
rect 247218 306212 247224 306264
rect 247276 306252 247282 306264
rect 247862 306252 247868 306264
rect 247276 306224 247868 306252
rect 247276 306212 247282 306224
rect 247862 306212 247868 306224
rect 247920 306212 247926 306264
rect 259546 306212 259552 306264
rect 259604 306252 259610 306264
rect 259914 306252 259920 306264
rect 259604 306224 259920 306252
rect 259604 306212 259610 306224
rect 259914 306212 259920 306224
rect 259972 306212 259978 306264
rect 263778 306212 263784 306264
rect 263836 306252 263842 306264
rect 264330 306252 264336 306264
rect 263836 306224 264336 306252
rect 263836 306212 263842 306224
rect 264330 306212 264336 306224
rect 264388 306212 264394 306264
rect 264974 306212 264980 306264
rect 265032 306252 265038 306264
rect 265894 306252 265900 306264
rect 265032 306224 265900 306252
rect 265032 306212 265038 306224
rect 265894 306212 265900 306224
rect 265952 306212 265958 306264
rect 266814 306212 266820 306264
rect 266872 306252 266878 306264
rect 267366 306252 267372 306264
rect 266872 306224 267372 306252
rect 266872 306212 266878 306224
rect 267366 306212 267372 306224
rect 267424 306212 267430 306264
rect 267734 306212 267740 306264
rect 267792 306252 267798 306264
rect 268470 306252 268476 306264
rect 267792 306224 268476 306252
rect 267792 306212 267798 306224
rect 268470 306212 268476 306224
rect 268528 306212 268534 306264
rect 270770 306212 270776 306264
rect 270828 306252 270834 306264
rect 271046 306252 271052 306264
rect 270828 306224 271052 306252
rect 270828 306212 270834 306224
rect 271046 306212 271052 306224
rect 271104 306212 271110 306264
rect 272150 306212 272156 306264
rect 272208 306252 272214 306264
rect 272794 306252 272800 306264
rect 272208 306224 272800 306252
rect 272208 306212 272214 306224
rect 272794 306212 272800 306224
rect 272852 306212 272858 306264
rect 273622 306212 273628 306264
rect 273680 306252 273686 306264
rect 273898 306252 273904 306264
rect 273680 306224 273904 306252
rect 273680 306212 273686 306224
rect 273898 306212 273904 306224
rect 273956 306212 273962 306264
rect 275922 306212 275928 306264
rect 275980 306252 275986 306264
rect 275980 306224 282914 306252
rect 275980 306212 275986 306224
rect 255498 306144 255504 306196
rect 255556 306184 255562 306196
rect 255866 306184 255872 306196
rect 255556 306156 255872 306184
rect 255556 306144 255562 306156
rect 255866 306144 255872 306156
rect 255924 306144 255930 306196
rect 260926 306144 260932 306196
rect 260984 306184 260990 306196
rect 261386 306184 261392 306196
rect 260984 306156 261392 306184
rect 260984 306144 260990 306156
rect 261386 306144 261392 306156
rect 261444 306144 261450 306196
rect 263962 306144 263968 306196
rect 264020 306184 264026 306196
rect 264790 306184 264796 306196
rect 264020 306156 264796 306184
rect 264020 306144 264026 306156
rect 264790 306144 264796 306156
rect 264848 306144 264854 306196
rect 266538 306144 266544 306196
rect 266596 306184 266602 306196
rect 267458 306184 267464 306196
rect 266596 306156 267464 306184
rect 266596 306144 266602 306156
rect 267458 306144 267464 306156
rect 267516 306144 267522 306196
rect 267826 306144 267832 306196
rect 267884 306184 267890 306196
rect 268930 306184 268936 306196
rect 267884 306156 268936 306184
rect 267884 306144 267890 306156
rect 268930 306144 268936 306156
rect 268988 306144 268994 306196
rect 270862 306144 270868 306196
rect 270920 306184 270926 306196
rect 271322 306184 271328 306196
rect 270920 306156 271328 306184
rect 270920 306144 270926 306156
rect 271322 306144 271328 306156
rect 271380 306144 271386 306196
rect 273254 306144 273260 306196
rect 273312 306184 273318 306196
rect 273806 306184 273812 306196
rect 273312 306156 273812 306184
rect 273312 306144 273318 306156
rect 273806 306144 273812 306156
rect 273864 306144 273870 306196
rect 274726 306144 274732 306196
rect 274784 306184 274790 306196
rect 275186 306184 275192 306196
rect 274784 306156 275192 306184
rect 274784 306144 274790 306156
rect 275186 306144 275192 306156
rect 275244 306144 275250 306196
rect 276290 306144 276296 306196
rect 276348 306184 276354 306196
rect 277026 306184 277032 306196
rect 276348 306156 277032 306184
rect 276348 306144 276354 306156
rect 277026 306144 277032 306156
rect 277084 306144 277090 306196
rect 277670 306144 277676 306196
rect 277728 306184 277734 306196
rect 278682 306184 278688 306196
rect 277728 306156 278688 306184
rect 277728 306144 277734 306156
rect 278682 306144 278688 306156
rect 278740 306144 278746 306196
rect 280246 306144 280252 306196
rect 280304 306184 280310 306196
rect 280706 306184 280712 306196
rect 280304 306156 280712 306184
rect 280304 306144 280310 306156
rect 280706 306144 280712 306156
rect 280764 306144 280770 306196
rect 281626 306144 281632 306196
rect 281684 306184 281690 306196
rect 282178 306184 282184 306196
rect 281684 306156 282184 306184
rect 281684 306144 281690 306156
rect 282178 306144 282184 306156
rect 282236 306144 282242 306196
rect 282886 306184 282914 306224
rect 283098 306212 283104 306264
rect 283156 306212 283162 306264
rect 283282 306212 283288 306264
rect 283340 306252 283346 306264
rect 283742 306252 283748 306264
rect 283340 306224 283748 306252
rect 283340 306212 283346 306224
rect 283742 306212 283748 306224
rect 283800 306212 283806 306264
rect 285766 306212 285772 306264
rect 285824 306252 285830 306264
rect 286502 306252 286508 306264
rect 285824 306224 286508 306252
rect 285824 306212 285830 306224
rect 286502 306212 286508 306224
rect 286560 306212 286566 306264
rect 288894 306212 288900 306264
rect 288952 306252 288958 306264
rect 289538 306252 289544 306264
rect 288952 306224 289544 306252
rect 288952 306212 288958 306224
rect 289538 306212 289544 306224
rect 289596 306212 289602 306264
rect 291562 306212 291568 306264
rect 291620 306252 291626 306264
rect 292114 306252 292120 306264
rect 291620 306224 292120 306252
rect 291620 306212 291626 306224
rect 292114 306212 292120 306224
rect 292172 306212 292178 306264
rect 292390 306212 292396 306264
rect 292448 306252 292454 306264
rect 331122 306252 331128 306264
rect 292448 306224 331128 306252
rect 292448 306212 292454 306224
rect 331122 306212 331128 306224
rect 331180 306212 331186 306264
rect 331398 306212 331404 306264
rect 331456 306252 331462 306264
rect 331950 306252 331956 306264
rect 331456 306224 331956 306252
rect 331456 306212 331462 306224
rect 331950 306212 331956 306224
rect 332008 306212 332014 306264
rect 332594 306212 332600 306264
rect 332652 306252 332658 306264
rect 332962 306252 332968 306264
rect 332652 306224 332968 306252
rect 332652 306212 332658 306224
rect 332962 306212 332968 306224
rect 333020 306212 333026 306264
rect 334158 306212 334164 306264
rect 334216 306252 334222 306264
rect 334710 306252 334716 306264
rect 334216 306224 334716 306252
rect 334216 306212 334222 306224
rect 334710 306212 334716 306224
rect 334768 306212 334774 306264
rect 335354 306212 335360 306264
rect 335412 306252 335418 306264
rect 335722 306252 335728 306264
rect 335412 306224 335728 306252
rect 335412 306212 335418 306224
rect 335722 306212 335728 306224
rect 335780 306212 335786 306264
rect 339678 306212 339684 306264
rect 339736 306252 339742 306264
rect 340322 306252 340328 306264
rect 339736 306224 340328 306252
rect 339736 306212 339742 306224
rect 340322 306212 340328 306224
rect 340380 306212 340386 306264
rect 340846 306252 340874 306292
rect 341058 306280 341064 306332
rect 341116 306320 341122 306332
rect 341426 306320 341432 306332
rect 341116 306292 341432 306320
rect 341116 306280 341122 306292
rect 341426 306280 341432 306292
rect 341484 306280 341490 306332
rect 342714 306320 342720 306332
rect 341536 306292 342720 306320
rect 341536 306252 341564 306292
rect 342714 306280 342720 306292
rect 342772 306280 342778 306332
rect 344094 306280 344100 306332
rect 344152 306320 344158 306332
rect 344922 306320 344928 306332
rect 344152 306292 344928 306320
rect 344152 306280 344158 306292
rect 344922 306280 344928 306292
rect 344980 306280 344986 306332
rect 345290 306280 345296 306332
rect 345348 306320 345354 306332
rect 345474 306320 345480 306332
rect 345348 306292 345480 306320
rect 345348 306280 345354 306292
rect 345474 306280 345480 306292
rect 345532 306280 345538 306332
rect 340846 306224 341564 306252
rect 342530 306212 342536 306264
rect 342588 306252 342594 306264
rect 343358 306252 343364 306264
rect 342588 306224 343364 306252
rect 342588 306212 342594 306224
rect 343358 306212 343364 306224
rect 343416 306212 343422 306264
rect 345014 306212 345020 306264
rect 345072 306252 345078 306264
rect 345842 306252 345848 306264
rect 345072 306224 345848 306252
rect 345072 306212 345078 306224
rect 345842 306212 345848 306224
rect 345900 306212 345906 306264
rect 347958 306212 347964 306264
rect 348016 306252 348022 306264
rect 348234 306252 348240 306264
rect 348016 306224 348240 306252
rect 348016 306212 348022 306224
rect 348234 306212 348240 306224
rect 348292 306212 348298 306264
rect 349338 306212 349344 306264
rect 349396 306252 349402 306264
rect 349890 306252 349896 306264
rect 349396 306224 349896 306252
rect 349396 306212 349402 306224
rect 349890 306212 349896 306224
rect 349948 306212 349954 306264
rect 341886 306184 341892 306196
rect 282886 306156 341892 306184
rect 341886 306144 341892 306156
rect 341944 306144 341950 306196
rect 345290 306144 345296 306196
rect 345348 306184 345354 306196
rect 346210 306184 346216 306196
rect 345348 306156 346216 306184
rect 345348 306144 345354 306156
rect 346210 306144 346216 306156
rect 346268 306144 346274 306196
rect 349246 306144 349252 306196
rect 349304 306184 349310 306196
rect 349614 306184 349620 306196
rect 349304 306156 349620 306184
rect 349304 306144 349310 306156
rect 349614 306144 349620 306156
rect 349672 306144 349678 306196
rect 230750 306076 230756 306128
rect 230808 306116 230814 306128
rect 231762 306116 231768 306128
rect 230808 306088 231768 306116
rect 230808 306076 230814 306088
rect 231762 306076 231768 306088
rect 231820 306076 231826 306128
rect 255682 306076 255688 306128
rect 255740 306116 255746 306128
rect 256326 306116 256332 306128
rect 255740 306088 256332 306116
rect 255740 306076 255746 306088
rect 256326 306076 256332 306088
rect 256384 306076 256390 306128
rect 257062 306076 257068 306128
rect 257120 306116 257126 306128
rect 257614 306116 257620 306128
rect 257120 306088 257620 306116
rect 257120 306076 257126 306088
rect 257614 306076 257620 306088
rect 257672 306076 257678 306128
rect 259546 306076 259552 306128
rect 259604 306116 259610 306128
rect 260650 306116 260656 306128
rect 259604 306088 260656 306116
rect 259604 306076 259610 306088
rect 260650 306076 260656 306088
rect 260708 306076 260714 306128
rect 279050 306076 279056 306128
rect 279108 306116 279114 306128
rect 279326 306116 279332 306128
rect 279108 306088 279332 306116
rect 279108 306076 279114 306088
rect 279326 306076 279332 306088
rect 279384 306076 279390 306128
rect 281718 306076 281724 306128
rect 281776 306116 281782 306128
rect 282362 306116 282368 306128
rect 281776 306088 282368 306116
rect 281776 306076 281782 306088
rect 282362 306076 282368 306088
rect 282420 306076 282426 306128
rect 344462 306116 344468 306128
rect 282886 306088 344468 306116
rect 254118 306008 254124 306060
rect 254176 306048 254182 306060
rect 255222 306048 255228 306060
rect 254176 306020 255228 306048
rect 254176 306008 254182 306020
rect 255222 306008 255228 306020
rect 255280 306008 255286 306060
rect 259730 306008 259736 306060
rect 259788 306048 259794 306060
rect 260466 306048 260472 306060
rect 259788 306020 260472 306048
rect 259788 306008 259794 306020
rect 260466 306008 260472 306020
rect 260524 306008 260530 306060
rect 260926 306008 260932 306060
rect 260984 306048 260990 306060
rect 261938 306048 261944 306060
rect 260984 306020 261944 306048
rect 260984 306008 260990 306020
rect 261938 306008 261944 306020
rect 261996 306008 262002 306060
rect 273254 306008 273260 306060
rect 273312 306048 273318 306060
rect 273990 306048 273996 306060
rect 273312 306020 273996 306048
rect 273312 306008 273318 306020
rect 273990 306008 273996 306020
rect 274048 306008 274054 306060
rect 274726 306008 274732 306060
rect 274784 306048 274790 306060
rect 275278 306048 275284 306060
rect 274784 306020 275284 306048
rect 274784 306008 274790 306020
rect 275278 306008 275284 306020
rect 275336 306008 275342 306060
rect 277302 306008 277308 306060
rect 277360 306048 277366 306060
rect 282886 306048 282914 306088
rect 344462 306076 344468 306088
rect 344520 306076 344526 306128
rect 349430 306076 349436 306128
rect 349488 306116 349494 306128
rect 350350 306116 350356 306128
rect 349488 306088 350356 306116
rect 349488 306076 349494 306088
rect 350350 306076 350356 306088
rect 350408 306076 350414 306128
rect 277360 306020 282914 306048
rect 277360 306008 277366 306020
rect 287422 306008 287428 306060
rect 287480 306048 287486 306060
rect 288250 306048 288256 306060
rect 287480 306020 288256 306048
rect 287480 306008 287486 306020
rect 288250 306008 288256 306020
rect 288308 306008 288314 306060
rect 288434 306008 288440 306060
rect 288492 306048 288498 306060
rect 289170 306048 289176 306060
rect 288492 306020 289176 306048
rect 288492 306008 288498 306020
rect 289170 306008 289176 306020
rect 289228 306008 289234 306060
rect 291470 306008 291476 306060
rect 291528 306048 291534 306060
rect 291930 306048 291936 306060
rect 291528 306020 291936 306048
rect 291528 306008 291534 306020
rect 291930 306008 291936 306020
rect 291988 306008 291994 306060
rect 292022 306008 292028 306060
rect 292080 306048 292086 306060
rect 351178 306048 351184 306060
rect 292080 306020 351184 306048
rect 292080 306008 292086 306020
rect 351178 306008 351184 306020
rect 351236 306008 351242 306060
rect 281074 305940 281080 305992
rect 281132 305980 281138 305992
rect 350626 305980 350632 305992
rect 281132 305952 350632 305980
rect 281132 305940 281138 305952
rect 350626 305940 350632 305952
rect 350684 305940 350690 305992
rect 282362 305872 282368 305924
rect 282420 305912 282426 305924
rect 352006 305912 352012 305924
rect 282420 305884 352012 305912
rect 282420 305872 282426 305884
rect 352006 305872 352012 305884
rect 352064 305872 352070 305924
rect 282270 305804 282276 305856
rect 282328 305844 282334 305856
rect 353754 305844 353760 305856
rect 282328 305816 353760 305844
rect 282328 305804 282334 305816
rect 353754 305804 353760 305816
rect 353812 305804 353818 305856
rect 282178 305736 282184 305788
rect 282236 305776 282242 305788
rect 353386 305776 353392 305788
rect 282236 305748 353392 305776
rect 282236 305736 282242 305748
rect 353386 305736 353392 305748
rect 353444 305736 353450 305788
rect 281166 305668 281172 305720
rect 281224 305708 281230 305720
rect 353662 305708 353668 305720
rect 281224 305680 353668 305708
rect 281224 305668 281230 305680
rect 353662 305668 353668 305680
rect 353720 305668 353726 305720
rect 82170 305600 82176 305652
rect 82228 305640 82234 305652
rect 241974 305640 241980 305652
rect 82228 305612 241980 305640
rect 82228 305600 82234 305612
rect 241974 305600 241980 305612
rect 242032 305600 242038 305652
rect 278682 305600 278688 305652
rect 278740 305640 278746 305652
rect 358814 305640 358820 305652
rect 278740 305612 358820 305640
rect 278740 305600 278746 305612
rect 358814 305600 358820 305612
rect 358872 305600 358878 305652
rect 291286 305532 291292 305584
rect 291344 305572 291350 305584
rect 292206 305572 292212 305584
rect 291344 305544 292212 305572
rect 291344 305532 291350 305544
rect 292206 305532 292212 305544
rect 292264 305532 292270 305584
rect 292850 305532 292856 305584
rect 292908 305572 292914 305584
rect 293310 305572 293316 305584
rect 292908 305544 293316 305572
rect 292908 305532 292914 305544
rect 293310 305532 293316 305544
rect 293368 305532 293374 305584
rect 294230 305532 294236 305584
rect 294288 305572 294294 305584
rect 294966 305572 294972 305584
rect 294288 305544 294972 305572
rect 294288 305532 294294 305544
rect 294966 305532 294972 305544
rect 295024 305532 295030 305584
rect 298370 305532 298376 305584
rect 298428 305572 298434 305584
rect 299106 305572 299112 305584
rect 298428 305544 299112 305572
rect 298428 305532 298434 305544
rect 299106 305532 299112 305544
rect 299164 305532 299170 305584
rect 300118 305532 300124 305584
rect 300176 305572 300182 305584
rect 300176 305544 331996 305572
rect 300176 305532 300182 305544
rect 284018 305464 284024 305516
rect 284076 305504 284082 305516
rect 292022 305504 292028 305516
rect 284076 305476 292028 305504
rect 284076 305464 284082 305476
rect 292022 305464 292028 305476
rect 292080 305464 292086 305516
rect 299566 305464 299572 305516
rect 299624 305504 299630 305516
rect 300578 305504 300584 305516
rect 299624 305476 300584 305504
rect 299624 305464 299630 305476
rect 300578 305464 300584 305476
rect 300636 305464 300642 305516
rect 331858 305504 331864 305516
rect 300780 305476 331864 305504
rect 296622 305328 296628 305380
rect 296680 305368 296686 305380
rect 296806 305368 296812 305380
rect 296680 305340 296812 305368
rect 296680 305328 296686 305340
rect 296806 305328 296812 305340
rect 296864 305328 296870 305380
rect 299198 305328 299204 305380
rect 299256 305368 299262 305380
rect 300780 305368 300808 305476
rect 331858 305464 331864 305476
rect 331916 305464 331922 305516
rect 299256 305340 300808 305368
rect 302206 305408 331904 305436
rect 299256 305328 299262 305340
rect 294966 305260 294972 305312
rect 295024 305300 295030 305312
rect 300118 305300 300124 305312
rect 295024 305272 300124 305300
rect 295024 305260 295030 305272
rect 300118 305260 300124 305272
rect 300176 305260 300182 305312
rect 285674 305192 285680 305244
rect 285732 305232 285738 305244
rect 286686 305232 286692 305244
rect 285732 305204 286692 305232
rect 285732 305192 285738 305204
rect 286686 305192 286692 305204
rect 286744 305192 286750 305244
rect 296622 305192 296628 305244
rect 296680 305232 296686 305244
rect 301590 305232 301596 305244
rect 296680 305204 301596 305232
rect 296680 305192 296686 305204
rect 301590 305192 301596 305204
rect 301648 305192 301654 305244
rect 283926 305124 283932 305176
rect 283984 305164 283990 305176
rect 284202 305164 284208 305176
rect 283984 305136 284208 305164
rect 283984 305124 283990 305136
rect 284202 305124 284208 305136
rect 284260 305124 284266 305176
rect 299474 305124 299480 305176
rect 299532 305164 299538 305176
rect 300210 305164 300216 305176
rect 299532 305136 300216 305164
rect 299532 305124 299538 305136
rect 300210 305124 300216 305136
rect 300268 305124 300274 305176
rect 299290 305056 299296 305108
rect 299348 305096 299354 305108
rect 302206 305096 302234 305408
rect 302326 305328 302332 305380
rect 302384 305368 302390 305380
rect 302786 305368 302792 305380
rect 302384 305340 302792 305368
rect 302384 305328 302390 305340
rect 302786 305328 302792 305340
rect 302844 305328 302850 305380
rect 306374 305328 306380 305380
rect 306432 305368 306438 305380
rect 306834 305368 306840 305380
rect 306432 305340 306840 305368
rect 306432 305328 306438 305340
rect 306834 305328 306840 305340
rect 306892 305328 306898 305380
rect 307938 305328 307944 305380
rect 307996 305368 308002 305380
rect 309042 305368 309048 305380
rect 307996 305340 309048 305368
rect 307996 305328 308002 305340
rect 309042 305328 309048 305340
rect 309100 305328 309106 305380
rect 310606 305328 310612 305380
rect 310664 305368 310670 305380
rect 310882 305368 310888 305380
rect 310664 305340 310888 305368
rect 310664 305328 310670 305340
rect 310882 305328 310888 305340
rect 310940 305328 310946 305380
rect 321646 305328 321652 305380
rect 321704 305368 321710 305380
rect 322290 305368 322296 305380
rect 321704 305340 322296 305368
rect 321704 305328 321710 305340
rect 322290 305328 322296 305340
rect 322348 305328 322354 305380
rect 323118 305328 323124 305380
rect 323176 305368 323182 305380
rect 323854 305368 323860 305380
rect 323176 305340 323860 305368
rect 323176 305328 323182 305340
rect 323854 305328 323860 305340
rect 323912 305328 323918 305380
rect 324498 305328 324504 305380
rect 324556 305368 324562 305380
rect 325142 305368 325148 305380
rect 324556 305340 325148 305368
rect 324556 305328 324562 305340
rect 325142 305328 325148 305340
rect 325200 305328 325206 305380
rect 328638 305328 328644 305380
rect 328696 305368 328702 305380
rect 329466 305368 329472 305380
rect 328696 305340 329472 305368
rect 328696 305328 328702 305340
rect 329466 305328 329472 305340
rect 329524 305328 329530 305380
rect 330018 305328 330024 305380
rect 330076 305368 330082 305380
rect 330570 305368 330576 305380
rect 330076 305340 330576 305368
rect 330076 305328 330082 305340
rect 330570 305328 330576 305340
rect 330628 305328 330634 305380
rect 331214 305328 331220 305380
rect 331272 305368 331278 305380
rect 331766 305368 331772 305380
rect 331272 305340 331772 305368
rect 331272 305328 331278 305340
rect 331766 305328 331772 305340
rect 331824 305328 331830 305380
rect 302602 305260 302608 305312
rect 302660 305300 302666 305312
rect 303430 305300 303436 305312
rect 302660 305272 303436 305300
rect 302660 305260 302666 305272
rect 303430 305260 303436 305272
rect 303488 305260 303494 305312
rect 306558 305260 306564 305312
rect 306616 305300 306622 305312
rect 307570 305300 307576 305312
rect 306616 305272 307576 305300
rect 306616 305260 306622 305272
rect 307570 305260 307576 305272
rect 307628 305260 307634 305312
rect 324314 305260 324320 305312
rect 324372 305300 324378 305312
rect 325418 305300 325424 305312
rect 324372 305272 325424 305300
rect 324372 305260 324378 305272
rect 325418 305260 325424 305272
rect 325476 305260 325482 305312
rect 328546 305260 328552 305312
rect 328604 305300 328610 305312
rect 329558 305300 329564 305312
rect 328604 305272 329564 305300
rect 328604 305260 328610 305272
rect 329558 305260 329564 305272
rect 329616 305260 329622 305312
rect 330110 305260 330116 305312
rect 330168 305300 330174 305312
rect 330846 305300 330852 305312
rect 330168 305272 330852 305300
rect 330168 305260 330174 305272
rect 330846 305260 330852 305272
rect 330904 305260 330910 305312
rect 302418 305192 302424 305244
rect 302476 305232 302482 305244
rect 303062 305232 303068 305244
rect 302476 305204 303068 305232
rect 302476 305192 302482 305204
rect 303062 305192 303068 305204
rect 303120 305192 303126 305244
rect 306374 305192 306380 305244
rect 306432 305232 306438 305244
rect 307202 305232 307208 305244
rect 306432 305204 307208 305232
rect 306432 305192 306438 305204
rect 307202 305192 307208 305204
rect 307260 305192 307266 305244
rect 310606 305192 310612 305244
rect 310664 305232 310670 305244
rect 311526 305232 311532 305244
rect 310664 305204 311532 305232
rect 310664 305192 310670 305204
rect 311526 305192 311532 305204
rect 311584 305192 311590 305244
rect 321554 305192 321560 305244
rect 321612 305232 321618 305244
rect 322382 305232 322388 305244
rect 321612 305204 322388 305232
rect 321612 305192 321618 305204
rect 322382 305192 322388 305204
rect 322440 305192 322446 305244
rect 329926 305192 329932 305244
rect 329984 305232 329990 305244
rect 330754 305232 330760 305244
rect 329984 305204 330760 305232
rect 329984 305192 329990 305204
rect 330754 305192 330760 305204
rect 330812 305192 330818 305244
rect 331876 305164 331904 305408
rect 331968 305300 331996 305544
rect 332962 305532 332968 305584
rect 333020 305572 333026 305584
rect 333698 305572 333704 305584
rect 333020 305544 333704 305572
rect 333020 305532 333026 305544
rect 333698 305532 333704 305544
rect 333756 305532 333762 305584
rect 334250 305532 334256 305584
rect 334308 305572 334314 305584
rect 334986 305572 334992 305584
rect 334308 305544 334992 305572
rect 334308 305532 334314 305544
rect 334986 305532 334992 305544
rect 335044 305532 335050 305584
rect 335538 305532 335544 305584
rect 335596 305572 335602 305584
rect 336642 305572 336648 305584
rect 335596 305544 336648 305572
rect 335596 305532 335602 305544
rect 336642 305532 336648 305544
rect 336700 305532 336706 305584
rect 339586 305532 339592 305584
rect 339644 305572 339650 305584
rect 340414 305572 340420 305584
rect 339644 305544 340420 305572
rect 339644 305532 339650 305544
rect 340414 305532 340420 305544
rect 340472 305532 340478 305584
rect 332778 305464 332784 305516
rect 332836 305504 332842 305516
rect 333238 305504 333244 305516
rect 332836 305476 333244 305504
rect 332836 305464 332842 305476
rect 333238 305464 333244 305476
rect 333296 305464 333302 305516
rect 335354 305464 335360 305516
rect 335412 305504 335418 305516
rect 336274 305504 336280 305516
rect 335412 305476 336280 305504
rect 335412 305464 335418 305476
rect 336274 305464 336280 305476
rect 336332 305464 336338 305516
rect 332686 305396 332692 305448
rect 332744 305436 332750 305448
rect 333606 305436 333612 305448
rect 332744 305408 333612 305436
rect 332744 305396 332750 305408
rect 333606 305396 333612 305408
rect 333664 305396 333670 305448
rect 332226 305328 332232 305380
rect 332284 305368 332290 305380
rect 338574 305368 338580 305380
rect 332284 305340 338580 305368
rect 332284 305328 332290 305340
rect 338574 305328 338580 305340
rect 338632 305328 338638 305380
rect 337930 305300 337936 305312
rect 331968 305272 337936 305300
rect 337930 305260 337936 305272
rect 337988 305260 337994 305312
rect 339954 305164 339960 305176
rect 331876 305136 339960 305164
rect 339954 305124 339960 305136
rect 340012 305124 340018 305176
rect 299348 305068 302234 305096
rect 299348 305056 299354 305068
rect 305086 305056 305092 305108
rect 305144 305096 305150 305108
rect 305822 305096 305828 305108
rect 305144 305068 305828 305096
rect 305144 305056 305150 305068
rect 305822 305056 305828 305068
rect 305880 305056 305886 305108
rect 331858 305056 331864 305108
rect 331916 305096 331922 305108
rect 340782 305096 340788 305108
rect 331916 305068 340788 305096
rect 331916 305056 331922 305068
rect 340782 305056 340788 305068
rect 340840 305056 340846 305108
rect 269298 304988 269304 305040
rect 269356 305028 269362 305040
rect 269666 305028 269672 305040
rect 269356 305000 269672 305028
rect 269356 304988 269362 305000
rect 269666 304988 269672 305000
rect 269724 304988 269730 305040
rect 331214 304988 331220 305040
rect 331272 305028 331278 305040
rect 332318 305028 332324 305040
rect 331272 305000 332324 305028
rect 331272 304988 331278 305000
rect 332318 304988 332324 305000
rect 332376 304988 332382 305040
rect 304534 304512 304540 304564
rect 304592 304512 304598 304564
rect 88978 304308 88984 304360
rect 89036 304348 89042 304360
rect 242986 304348 242992 304360
rect 89036 304320 242992 304348
rect 89036 304308 89042 304320
rect 242986 304308 242992 304320
rect 243044 304308 243050 304360
rect 303614 304308 303620 304360
rect 303672 304348 303678 304360
rect 304074 304348 304080 304360
rect 303672 304320 304080 304348
rect 303672 304308 303678 304320
rect 304074 304308 304080 304320
rect 304132 304308 304138 304360
rect 7558 304240 7564 304292
rect 7616 304280 7622 304292
rect 230474 304280 230480 304292
rect 7616 304252 230480 304280
rect 7616 304240 7622 304252
rect 230474 304240 230480 304252
rect 230532 304240 230538 304292
rect 251450 304240 251456 304292
rect 251508 304280 251514 304292
rect 251726 304280 251732 304292
rect 251508 304252 251732 304280
rect 251508 304240 251514 304252
rect 251726 304240 251732 304252
rect 251784 304240 251790 304292
rect 271966 304240 271972 304292
rect 272024 304280 272030 304292
rect 272242 304280 272248 304292
rect 272024 304252 272248 304280
rect 272024 304240 272030 304252
rect 272242 304240 272248 304252
rect 272300 304240 272306 304292
rect 287054 304240 287060 304292
rect 287112 304280 287118 304292
rect 287882 304280 287888 304292
rect 287112 304252 287888 304280
rect 287112 304240 287118 304252
rect 287882 304240 287888 304252
rect 287940 304240 287946 304292
rect 303614 304172 303620 304224
rect 303672 304212 303678 304224
rect 304552 304212 304580 304512
rect 315390 304444 315396 304496
rect 315448 304484 315454 304496
rect 458818 304484 458824 304496
rect 315448 304456 458824 304484
rect 315448 304444 315454 304456
rect 458818 304444 458824 304456
rect 458876 304444 458882 304496
rect 319254 304376 319260 304428
rect 319312 304416 319318 304428
rect 478138 304416 478144 304428
rect 319312 304388 478144 304416
rect 319312 304376 319318 304388
rect 478138 304376 478144 304388
rect 478196 304376 478202 304428
rect 324682 304308 324688 304360
rect 324740 304348 324746 304360
rect 514018 304348 514024 304360
rect 324740 304320 514024 304348
rect 324740 304308 324746 304320
rect 514018 304308 514024 304320
rect 514076 304308 514082 304360
rect 305178 304240 305184 304292
rect 305236 304280 305242 304292
rect 305454 304280 305460 304292
rect 305236 304252 305460 304280
rect 305236 304240 305242 304252
rect 305454 304240 305460 304252
rect 305512 304240 305518 304292
rect 309226 304240 309232 304292
rect 309284 304280 309290 304292
rect 309594 304280 309600 304292
rect 309284 304252 309600 304280
rect 309284 304240 309290 304252
rect 309594 304240 309600 304252
rect 309652 304240 309658 304292
rect 310790 304240 310796 304292
rect 310848 304280 310854 304292
rect 311066 304280 311072 304292
rect 310848 304252 311072 304280
rect 310848 304240 310854 304252
rect 311066 304240 311072 304252
rect 311124 304240 311130 304292
rect 334526 304240 334532 304292
rect 334584 304280 334590 304292
rect 566458 304280 566464 304292
rect 334584 304252 566464 304280
rect 334584 304240 334590 304252
rect 566458 304240 566464 304252
rect 566516 304240 566522 304292
rect 303672 304184 304580 304212
rect 303672 304172 303678 304184
rect 250162 303696 250168 303748
rect 250220 303736 250226 303748
rect 251082 303736 251088 303748
rect 250220 303708 251088 303736
rect 250220 303696 250226 303708
rect 251082 303696 251088 303708
rect 251140 303696 251146 303748
rect 280982 303560 280988 303612
rect 281040 303600 281046 303612
rect 354674 303600 354680 303612
rect 281040 303572 354680 303600
rect 281040 303560 281046 303572
rect 354674 303560 354680 303572
rect 354732 303560 354738 303612
rect 268470 303492 268476 303544
rect 268528 303532 268534 303544
rect 344738 303532 344744 303544
rect 268528 303504 344744 303532
rect 268528 303492 268534 303504
rect 344738 303492 344744 303504
rect 344796 303492 344802 303544
rect 268562 303424 268568 303476
rect 268620 303464 268626 303476
rect 343818 303464 343824 303476
rect 268620 303436 343824 303464
rect 268620 303424 268626 303436
rect 343818 303424 343824 303436
rect 343876 303424 343882 303476
rect 279602 303356 279608 303408
rect 279660 303396 279666 303408
rect 356054 303396 356060 303408
rect 279660 303368 356060 303396
rect 279660 303356 279666 303368
rect 356054 303356 356060 303368
rect 356112 303356 356118 303408
rect 279510 303288 279516 303340
rect 279568 303328 279574 303340
rect 356146 303328 356152 303340
rect 279568 303300 356152 303328
rect 279568 303288 279574 303300
rect 356146 303288 356152 303300
rect 356204 303288 356210 303340
rect 268378 303220 268384 303272
rect 268436 303260 268442 303272
rect 345566 303260 345572 303272
rect 268436 303232 345572 303260
rect 268436 303220 268442 303232
rect 345566 303220 345572 303232
rect 345624 303220 345630 303272
rect 276934 303152 276940 303204
rect 276992 303192 276998 303204
rect 357526 303192 357532 303204
rect 276992 303164 357532 303192
rect 276992 303152 276998 303164
rect 357526 303152 357532 303164
rect 357584 303152 357590 303204
rect 245654 303124 245660 303136
rect 244246 303096 245660 303124
rect 85574 303016 85580 303068
rect 85632 303056 85638 303068
rect 244246 303056 244274 303096
rect 245654 303084 245660 303096
rect 245712 303084 245718 303136
rect 251358 303084 251364 303136
rect 251416 303124 251422 303136
rect 252278 303124 252284 303136
rect 251416 303096 252284 303124
rect 251416 303084 251422 303096
rect 252278 303084 252284 303096
rect 252336 303084 252342 303136
rect 276842 303084 276848 303136
rect 276900 303124 276906 303136
rect 357434 303124 357440 303136
rect 276900 303096 357440 303124
rect 276900 303084 276906 303096
rect 357434 303084 357440 303096
rect 357492 303084 357498 303136
rect 85632 303028 244274 303056
rect 85632 303016 85638 303028
rect 244366 303016 244372 303068
rect 244424 303016 244430 303068
rect 276750 303016 276756 303068
rect 276808 303056 276814 303068
rect 359366 303056 359372 303068
rect 276808 303028 359372 303056
rect 276808 303016 276814 303028
rect 359366 303016 359372 303028
rect 359424 303016 359430 303068
rect 77294 302948 77300 303000
rect 77352 302988 77358 303000
rect 244384 302988 244412 303016
rect 77352 302960 244412 302988
rect 77352 302948 77358 302960
rect 274082 302948 274088 303000
rect 274140 302988 274146 303000
rect 358906 302988 358912 303000
rect 274140 302960 358912 302988
rect 274140 302948 274146 302960
rect 358906 302948 358912 302960
rect 358964 302948 358970 303000
rect 8938 302880 8944 302932
rect 8996 302920 9002 302932
rect 231394 302920 231400 302932
rect 8996 302892 231400 302920
rect 8996 302880 9002 302892
rect 231394 302880 231400 302892
rect 231452 302880 231458 302932
rect 244366 302880 244372 302932
rect 244424 302920 244430 302932
rect 245102 302920 245108 302932
rect 244424 302892 245108 302920
rect 244424 302880 244430 302892
rect 245102 302880 245108 302892
rect 245160 302880 245166 302932
rect 273898 302880 273904 302932
rect 273956 302920 273962 302932
rect 360562 302920 360568 302932
rect 273956 302892 360568 302920
rect 273956 302880 273962 302892
rect 360562 302880 360568 302892
rect 360620 302880 360626 302932
rect 271230 302812 271236 302864
rect 271288 302852 271294 302864
rect 342990 302852 342996 302864
rect 271288 302824 342996 302852
rect 271288 302812 271294 302824
rect 342990 302812 342996 302824
rect 343048 302812 343054 302864
rect 271414 302744 271420 302796
rect 271472 302784 271478 302796
rect 342070 302784 342076 302796
rect 271472 302756 342076 302784
rect 271472 302744 271478 302756
rect 342070 302744 342076 302756
rect 342128 302744 342134 302796
rect 251266 302676 251272 302728
rect 251324 302716 251330 302728
rect 251818 302716 251824 302728
rect 251324 302688 251824 302716
rect 251324 302676 251330 302688
rect 251818 302676 251824 302688
rect 251876 302676 251882 302728
rect 271322 302676 271328 302728
rect 271380 302716 271386 302728
rect 340966 302716 340972 302728
rect 271380 302688 340972 302716
rect 271380 302676 271386 302688
rect 340966 302676 340972 302688
rect 341024 302676 341030 302728
rect 269298 302336 269304 302388
rect 269356 302376 269362 302388
rect 270218 302376 270224 302388
rect 269356 302348 270224 302376
rect 269356 302336 269362 302348
rect 270218 302336 270224 302348
rect 270276 302336 270282 302388
rect 343818 302200 343824 302252
rect 343876 302240 343882 302252
rect 344278 302240 344284 302252
rect 343876 302212 344284 302240
rect 343876 302200 343882 302212
rect 344278 302200 344284 302212
rect 344336 302200 344342 302252
rect 292758 301996 292764 302048
rect 292816 302036 292822 302048
rect 293034 302036 293040 302048
rect 292816 302008 293040 302036
rect 292816 301996 292822 302008
rect 293034 301996 293040 302008
rect 293092 301996 293098 302048
rect 95878 301588 95884 301640
rect 95936 301628 95942 301640
rect 247586 301628 247592 301640
rect 95936 301600 247592 301628
rect 95936 301588 95942 301600
rect 247586 301588 247592 301600
rect 247644 301588 247650 301640
rect 316586 301588 316592 301640
rect 316644 301628 316650 301640
rect 468478 301628 468484 301640
rect 316644 301600 468484 301628
rect 316644 301588 316650 301600
rect 468478 301588 468484 301600
rect 468536 301588 468542 301640
rect 93854 301520 93860 301572
rect 93912 301560 93918 301572
rect 247126 301560 247132 301572
rect 93912 301532 247132 301560
rect 93912 301520 93918 301532
rect 247126 301520 247132 301532
rect 247184 301520 247190 301572
rect 320634 301520 320640 301572
rect 320692 301560 320698 301572
rect 494054 301560 494060 301572
rect 320692 301532 494060 301560
rect 320692 301520 320698 301532
rect 494054 301520 494060 301532
rect 494112 301520 494118 301572
rect 48958 301452 48964 301504
rect 49016 301492 49022 301504
rect 239122 301492 239128 301504
rect 49016 301464 239128 301492
rect 49016 301452 49022 301464
rect 239122 301452 239128 301464
rect 239180 301452 239186 301504
rect 329374 301452 329380 301504
rect 329432 301492 329438 301504
rect 534718 301492 534724 301504
rect 329432 301464 534724 301492
rect 329432 301452 329438 301464
rect 534718 301452 534724 301464
rect 534776 301452 534782 301504
rect 288710 301248 288716 301300
rect 288768 301288 288774 301300
rect 289078 301288 289084 301300
rect 288768 301260 289084 301288
rect 288768 301248 288774 301260
rect 289078 301248 289084 301260
rect 289136 301248 289142 301300
rect 290918 300772 290924 300824
rect 290976 300812 290982 300824
rect 342438 300812 342444 300824
rect 290976 300784 342444 300812
rect 290976 300772 290982 300784
rect 342438 300772 342444 300784
rect 342496 300772 342502 300824
rect 289538 300704 289544 300756
rect 289596 300744 289602 300756
rect 341058 300744 341064 300756
rect 289596 300716 341064 300744
rect 289596 300704 289602 300716
rect 341058 300704 341064 300716
rect 341116 300704 341122 300756
rect 286778 300636 286784 300688
rect 286836 300676 286842 300688
rect 338298 300676 338304 300688
rect 286836 300648 338304 300676
rect 286836 300636 286842 300648
rect 338298 300636 338304 300648
rect 338356 300636 338362 300688
rect 289446 300568 289452 300620
rect 289504 300608 289510 300620
rect 344186 300608 344192 300620
rect 289504 300580 344192 300608
rect 289504 300568 289510 300580
rect 344186 300568 344192 300580
rect 344244 300568 344250 300620
rect 283926 300500 283932 300552
rect 283984 300540 283990 300552
rect 338206 300540 338212 300552
rect 283984 300512 338212 300540
rect 283984 300500 283990 300512
rect 338206 300500 338212 300512
rect 338264 300500 338270 300552
rect 286594 300432 286600 300484
rect 286652 300472 286658 300484
rect 343174 300472 343180 300484
rect 286652 300444 343180 300472
rect 286652 300432 286658 300444
rect 343174 300432 343180 300444
rect 343232 300432 343238 300484
rect 286870 300364 286876 300416
rect 286928 300404 286934 300416
rect 346578 300404 346584 300416
rect 286928 300376 346584 300404
rect 286928 300364 286934 300376
rect 346578 300364 346584 300376
rect 346636 300364 346642 300416
rect 285306 300296 285312 300348
rect 285364 300336 285370 300348
rect 345014 300336 345020 300348
rect 285364 300308 345020 300336
rect 285364 300296 285370 300308
rect 345014 300296 345020 300308
rect 345072 300296 345078 300348
rect 282730 300228 282736 300280
rect 282788 300268 282794 300280
rect 352466 300268 352472 300280
rect 282788 300240 352472 300268
rect 282788 300228 282794 300240
rect 352466 300228 352472 300240
rect 352524 300228 352530 300280
rect 53098 300160 53104 300212
rect 53156 300200 53162 300212
rect 238846 300200 238852 300212
rect 53156 300172 238852 300200
rect 53156 300160 53162 300172
rect 238846 300160 238852 300172
rect 238904 300160 238910 300212
rect 278406 300160 278412 300212
rect 278464 300200 278470 300212
rect 349522 300200 349528 300212
rect 278464 300172 349528 300200
rect 278464 300160 278470 300172
rect 349522 300160 349528 300172
rect 349580 300160 349586 300212
rect 40034 300092 40040 300144
rect 40092 300132 40098 300144
rect 237374 300132 237380 300144
rect 40092 300104 237380 300132
rect 40092 300092 40098 300104
rect 237374 300092 237380 300104
rect 237432 300092 237438 300144
rect 278498 300092 278504 300144
rect 278556 300132 278562 300144
rect 349338 300132 349344 300144
rect 278556 300104 349344 300132
rect 278556 300092 278562 300104
rect 349338 300092 349344 300104
rect 349396 300092 349402 300144
rect 288250 300024 288256 300076
rect 288308 300064 288314 300076
rect 339678 300064 339684 300076
rect 288308 300036 339684 300064
rect 288308 300024 288314 300036
rect 339678 300024 339684 300036
rect 339736 300024 339742 300076
rect 285122 299956 285128 300008
rect 285180 299996 285186 300008
rect 337102 299996 337108 300008
rect 285180 299968 337108 299996
rect 285180 299956 285186 299968
rect 337102 299956 337108 299968
rect 337160 299956 337166 300008
rect 292206 299888 292212 299940
rect 292264 299928 292270 299940
rect 340138 299928 340144 299940
rect 292264 299900 340144 299928
rect 292264 299888 292270 299900
rect 340138 299888 340144 299900
rect 340196 299888 340202 299940
rect 322750 298868 322756 298920
rect 322808 298908 322814 298920
rect 502978 298908 502984 298920
rect 322808 298880 502984 298908
rect 322808 298868 322814 298880
rect 502978 298868 502984 298880
rect 503036 298868 503042 298920
rect 53834 298800 53840 298852
rect 53892 298840 53898 298852
rect 238754 298840 238760 298852
rect 53892 298812 238760 298840
rect 53892 298800 53898 298812
rect 238754 298800 238760 298812
rect 238812 298800 238818 298852
rect 331766 298800 331772 298852
rect 331824 298840 331830 298852
rect 549898 298840 549904 298852
rect 331824 298812 549904 298840
rect 331824 298800 331830 298812
rect 549898 298800 549904 298812
rect 549956 298800 549962 298852
rect 10318 298732 10324 298784
rect 10376 298772 10382 298784
rect 231026 298772 231032 298784
rect 10376 298744 231032 298772
rect 10376 298732 10382 298744
rect 231026 298732 231032 298744
rect 231084 298732 231090 298784
rect 239398 298732 239404 298784
rect 239456 298772 239462 298784
rect 251542 298772 251548 298784
rect 239456 298744 251548 298772
rect 239456 298732 239462 298744
rect 251542 298732 251548 298744
rect 251600 298732 251606 298784
rect 334342 298732 334348 298784
rect 334400 298772 334406 298784
rect 563698 298772 563704 298784
rect 334400 298744 563704 298772
rect 334400 298732 334406 298744
rect 563698 298732 563704 298744
rect 563756 298732 563762 298784
rect 298002 297984 298008 298036
rect 298060 298024 298066 298036
rect 356330 298024 356336 298036
rect 298060 297996 356336 298024
rect 298060 297984 298066 297996
rect 356330 297984 356336 297996
rect 356388 297984 356394 298036
rect 297910 297916 297916 297968
rect 297968 297956 297974 297968
rect 356238 297956 356244 297968
rect 297968 297928 356244 297956
rect 297968 297916 297974 297928
rect 356238 297916 356244 297928
rect 356296 297916 356302 297968
rect 277210 297848 277216 297900
rect 277268 297888 277274 297900
rect 338390 297888 338396 297900
rect 277268 297860 338396 297888
rect 277268 297848 277274 297860
rect 338390 297848 338396 297860
rect 338448 297848 338454 297900
rect 278314 297780 278320 297832
rect 278372 297820 278378 297832
rect 341518 297820 341524 297832
rect 278372 297792 341524 297820
rect 278372 297780 278378 297792
rect 341518 297780 341524 297792
rect 341576 297780 341582 297832
rect 284846 297712 284852 297764
rect 284904 297752 284910 297764
rect 360286 297752 360292 297764
rect 284904 297724 360292 297752
rect 284904 297712 284910 297724
rect 360286 297712 360292 297724
rect 360344 297712 360350 297764
rect 279970 297644 279976 297696
rect 280028 297684 280034 297696
rect 359090 297684 359096 297696
rect 280028 297656 359096 297684
rect 280028 297644 280034 297656
rect 359090 297644 359096 297656
rect 359148 297644 359154 297696
rect 317966 297576 317972 297628
rect 318024 297616 318030 297628
rect 462958 297616 462964 297628
rect 318024 297588 462964 297616
rect 318024 297576 318030 297588
rect 462958 297576 462964 297588
rect 463016 297576 463022 297628
rect 316218 297508 316224 297560
rect 316276 297548 316282 297560
rect 473446 297548 473452 297560
rect 316276 297520 473452 297548
rect 316276 297508 316282 297520
rect 473446 297508 473452 297520
rect 473504 297508 473510 297560
rect 60734 297440 60740 297492
rect 60792 297480 60798 297492
rect 241330 297480 241336 297492
rect 60792 297452 241336 297480
rect 60792 297440 60798 297452
rect 241330 297440 241336 297452
rect 241388 297440 241394 297492
rect 285858 297440 285864 297492
rect 285916 297440 285922 297492
rect 323394 297440 323400 297492
rect 323452 297480 323458 297492
rect 507854 297480 507860 297492
rect 323452 297452 507860 297480
rect 323452 297440 323458 297452
rect 507854 297440 507860 297452
rect 507912 297440 507918 297492
rect 62114 297372 62120 297424
rect 62172 297412 62178 297424
rect 241790 297412 241796 297424
rect 62172 297384 241796 297412
rect 62172 297372 62178 297384
rect 241790 297372 241796 297384
rect 241848 297372 241854 297424
rect 285876 297276 285904 297440
rect 333146 297372 333152 297424
rect 333204 297412 333210 297424
rect 561674 297412 561680 297424
rect 333204 297384 561680 297412
rect 333204 297372 333210 297384
rect 561674 297372 561680 297384
rect 561732 297372 561738 297424
rect 285950 297276 285956 297288
rect 285876 297248 285956 297276
rect 285950 297236 285956 297248
rect 286008 297236 286014 297288
rect 323302 296080 323308 296132
rect 323360 296120 323366 296132
rect 511994 296120 512000 296132
rect 323360 296092 512000 296120
rect 323360 296080 323366 296092
rect 511994 296080 512000 296092
rect 512052 296080 512058 296132
rect 71038 296012 71044 296064
rect 71096 296052 71102 296064
rect 243446 296052 243452 296064
rect 71096 296024 243452 296052
rect 71096 296012 71102 296024
rect 243446 296012 243452 296024
rect 243504 296012 243510 296064
rect 330110 296012 330116 296064
rect 330168 296052 330174 296064
rect 548518 296052 548524 296064
rect 330168 296024 548524 296052
rect 330168 296012 330174 296024
rect 548518 296012 548524 296024
rect 548576 296012 548582 296064
rect 66898 295944 66904 295996
rect 66956 295984 66962 295996
rect 241698 295984 241704 295996
rect 66956 295956 241704 295984
rect 66956 295944 66962 295956
rect 241698 295944 241704 295956
rect 241756 295944 241762 295996
rect 334250 295944 334256 295996
rect 334308 295984 334314 295996
rect 570598 295984 570604 295996
rect 334308 295956 570604 295984
rect 334308 295944 334314 295956
rect 570598 295944 570604 295956
rect 570656 295944 570662 295996
rect 321830 294720 321836 294772
rect 321888 294760 321894 294772
rect 493318 294760 493324 294772
rect 321888 294732 493324 294760
rect 321888 294720 321894 294732
rect 493318 294720 493324 294732
rect 493376 294720 493382 294772
rect 325970 294652 325976 294704
rect 326028 294692 326034 294704
rect 521654 294692 521660 294704
rect 326028 294664 521660 294692
rect 326028 294652 326034 294664
rect 521654 294652 521660 294664
rect 521712 294652 521718 294704
rect 69014 294584 69020 294636
rect 69072 294624 69078 294636
rect 241606 294624 241612 294636
rect 69072 294596 241612 294624
rect 69072 294584 69078 294596
rect 241606 294584 241612 294596
rect 241664 294584 241670 294636
rect 327534 294584 327540 294636
rect 327592 294624 327598 294636
rect 529934 294624 529940 294636
rect 327592 294596 529940 294624
rect 327592 294584 327598 294596
rect 529934 294584 529940 294596
rect 529992 294584 529998 294636
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 228450 293944 228456 293956
rect 3384 293916 228456 293944
rect 3384 293904 3390 293916
rect 228450 293904 228456 293916
rect 228508 293904 228514 293956
rect 325878 293360 325884 293412
rect 325936 293400 325942 293412
rect 522298 293400 522304 293412
rect 325936 293372 522304 293400
rect 325936 293360 325942 293372
rect 522298 293360 522304 293372
rect 522356 293360 522362 293412
rect 327442 293292 327448 293344
rect 327500 293332 327506 293344
rect 527818 293332 527824 293344
rect 327500 293304 527824 293332
rect 327500 293292 327506 293304
rect 527818 293292 527824 293304
rect 527876 293292 527882 293344
rect 86954 293224 86960 293276
rect 87012 293264 87018 293276
rect 246022 293264 246028 293276
rect 87012 293236 246028 293264
rect 87012 293224 87018 293236
rect 246022 293224 246028 293236
rect 246080 293224 246086 293276
rect 335814 293224 335820 293276
rect 335872 293264 335878 293276
rect 578234 293264 578240 293276
rect 335872 293236 578240 293264
rect 335872 293224 335878 293236
rect 578234 293224 578240 293236
rect 578292 293224 578298 293276
rect 71774 291864 71780 291916
rect 71832 291904 71838 291916
rect 243170 291904 243176 291916
rect 71832 291876 243176 291904
rect 71832 291864 71838 291876
rect 243170 291864 243176 291876
rect 243228 291864 243234 291916
rect 328822 291864 328828 291916
rect 328880 291904 328886 291916
rect 536098 291904 536104 291916
rect 328880 291876 536104 291904
rect 328880 291864 328886 291876
rect 536098 291864 536104 291876
rect 536156 291864 536162 291916
rect 30374 291796 30380 291848
rect 30432 291836 30438 291848
rect 234982 291836 234988 291848
rect 30432 291808 234988 291836
rect 30432 291796 30438 291808
rect 234982 291796 234988 291808
rect 235040 291796 235046 291848
rect 328914 291796 328920 291848
rect 328972 291836 328978 291848
rect 538858 291836 538864 291848
rect 328972 291808 538864 291836
rect 328972 291796 328978 291808
rect 538858 291796 538864 291808
rect 538916 291796 538922 291848
rect 75914 290504 75920 290556
rect 75972 290544 75978 290556
rect 243078 290544 243084 290556
rect 75972 290516 243084 290544
rect 75972 290504 75978 290516
rect 243078 290504 243084 290516
rect 243136 290504 243142 290556
rect 330018 290504 330024 290556
rect 330076 290544 330082 290556
rect 547966 290544 547972 290556
rect 330076 290516 547972 290544
rect 330076 290504 330082 290516
rect 547966 290504 547972 290516
rect 548024 290504 548030 290556
rect 41414 290436 41420 290488
rect 41472 290476 41478 290488
rect 237742 290476 237748 290488
rect 41472 290448 237748 290476
rect 41472 290436 41478 290448
rect 237742 290436 237748 290448
rect 237800 290436 237806 290488
rect 243630 290436 243636 290488
rect 243688 290476 243694 290488
rect 252922 290476 252928 290488
rect 243688 290448 252928 290476
rect 243688 290436 243694 290448
rect 252922 290436 252928 290448
rect 252980 290436 252986 290488
rect 334158 290436 334164 290488
rect 334216 290476 334222 290488
rect 567838 290476 567844 290488
rect 334216 290448 567844 290476
rect 334216 290436 334222 290448
rect 567838 290436 567844 290448
rect 567896 290436 567902 290488
rect 310974 289212 310980 289264
rect 311032 289252 311038 289264
rect 440234 289252 440240 289264
rect 311032 289224 440240 289252
rect 311032 289212 311038 289224
rect 440234 289212 440240 289224
rect 440292 289212 440298 289264
rect 56594 289144 56600 289196
rect 56652 289184 56658 289196
rect 240410 289184 240416 289196
rect 56652 289156 240416 289184
rect 56652 289144 56658 289156
rect 240410 289144 240416 289156
rect 240468 289144 240474 289196
rect 331674 289144 331680 289196
rect 331732 289184 331738 289196
rect 552658 289184 552664 289196
rect 331732 289156 552664 289184
rect 331732 289144 331738 289156
rect 552658 289144 552664 289156
rect 552716 289144 552722 289196
rect 13078 289076 13084 289128
rect 13136 289116 13142 289128
rect 232130 289116 232136 289128
rect 13136 289088 232136 289116
rect 13136 289076 13142 289088
rect 232130 289076 232136 289088
rect 232188 289076 232194 289128
rect 335722 289076 335728 289128
rect 335780 289116 335786 289128
rect 571978 289116 571984 289128
rect 335780 289088 571984 289116
rect 335780 289076 335786 289088
rect 571978 289076 571984 289088
rect 572036 289076 572042 289128
rect 313918 287716 313924 287768
rect 313976 287756 313982 287768
rect 449894 287756 449900 287768
rect 313976 287728 449900 287756
rect 313976 287716 313982 287728
rect 449894 287716 449900 287728
rect 449952 287716 449958 287768
rect 9674 287648 9680 287700
rect 9732 287688 9738 287700
rect 230750 287688 230756 287700
rect 9732 287660 230756 287688
rect 9732 287648 9738 287660
rect 230750 287648 230756 287660
rect 230808 287648 230814 287700
rect 331582 287648 331588 287700
rect 331640 287688 331646 287700
rect 557534 287688 557540 287700
rect 331640 287660 557540 287688
rect 331640 287648 331646 287660
rect 557534 287648 557540 287660
rect 557592 287648 557598 287700
rect 312262 286492 312268 286544
rect 312320 286532 312326 286544
rect 448514 286532 448520 286544
rect 312320 286504 448520 286532
rect 312320 286492 312326 286504
rect 448514 286492 448520 286504
rect 448572 286492 448578 286544
rect 318058 286424 318064 286476
rect 318116 286464 318122 286476
rect 456886 286464 456892 286476
rect 318116 286436 456892 286464
rect 318116 286424 318122 286436
rect 456886 286424 456892 286436
rect 456944 286424 456950 286476
rect 89714 286356 89720 286408
rect 89772 286396 89778 286408
rect 245930 286396 245936 286408
rect 89772 286368 245936 286396
rect 89772 286356 89778 286368
rect 245930 286356 245936 286368
rect 245988 286356 245994 286408
rect 313642 286356 313648 286408
rect 313700 286396 313706 286408
rect 456794 286396 456800 286408
rect 313700 286368 456800 286396
rect 313700 286356 313706 286368
rect 456794 286356 456800 286368
rect 456852 286356 456858 286408
rect 46290 286288 46296 286340
rect 46348 286328 46354 286340
rect 237650 286328 237656 286340
rect 46348 286300 237656 286328
rect 46348 286288 46354 286300
rect 237650 286288 237656 286300
rect 237708 286288 237714 286340
rect 332962 286288 332968 286340
rect 333020 286328 333026 286340
rect 563790 286328 563796 286340
rect 333020 286300 563796 286328
rect 333020 286288 333026 286300
rect 563790 286288 563796 286300
rect 563848 286288 563854 286340
rect 310790 285064 310796 285116
rect 310848 285104 310854 285116
rect 440326 285104 440332 285116
rect 310848 285076 440332 285104
rect 310848 285064 310854 285076
rect 440326 285064 440332 285076
rect 440384 285064 440390 285116
rect 324682 284996 324688 285048
rect 324740 285036 324746 285048
rect 516134 285036 516140 285048
rect 324740 285008 516140 285036
rect 324740 284996 324746 285008
rect 516134 284996 516140 285008
rect 516192 284996 516198 285048
rect 34514 284928 34520 284980
rect 34572 284968 34578 284980
rect 236270 284968 236276 284980
rect 34572 284940 236276 284968
rect 34572 284928 34578 284940
rect 236270 284928 236276 284940
rect 236328 284928 236334 284980
rect 328730 284928 328736 284980
rect 328788 284968 328794 284980
rect 535454 284968 535460 284980
rect 328788 284940 535460 284968
rect 328788 284928 328794 284940
rect 535454 284928 535460 284940
rect 535512 284928 535518 284980
rect 310698 283704 310704 283756
rect 310756 283744 310762 283756
rect 442994 283744 443000 283756
rect 310756 283716 443000 283744
rect 310756 283704 310762 283716
rect 442994 283704 443000 283716
rect 443052 283704 443058 283756
rect 60826 283636 60832 283688
rect 60884 283676 60890 283688
rect 240318 283676 240324 283688
rect 60884 283648 240324 283676
rect 60884 283636 60890 283648
rect 240318 283636 240324 283648
rect 240376 283636 240382 283688
rect 313550 283636 313556 283688
rect 313608 283676 313614 283688
rect 454678 283676 454684 283688
rect 313608 283648 454684 283676
rect 313608 283636 313614 283648
rect 454678 283636 454684 283648
rect 454736 283636 454742 283688
rect 16574 283568 16580 283620
rect 16632 283608 16638 283620
rect 232038 283608 232044 283620
rect 16632 283580 232044 283608
rect 16632 283568 16638 283580
rect 232038 283568 232044 283580
rect 232096 283568 232102 283620
rect 332870 283568 332876 283620
rect 332928 283608 332934 283620
rect 554038 283608 554044 283620
rect 332928 283580 554044 283608
rect 332928 283568 332934 283580
rect 554038 283568 554044 283580
rect 554096 283568 554102 283620
rect 313458 282276 313464 282328
rect 313516 282316 313522 282328
rect 450538 282316 450544 282328
rect 313516 282288 450544 282316
rect 313516 282276 313522 282288
rect 450538 282276 450544 282288
rect 450596 282276 450602 282328
rect 70394 282208 70400 282260
rect 70452 282248 70458 282260
rect 233878 282248 233884 282260
rect 70452 282220 233884 282248
rect 70452 282208 70458 282220
rect 233878 282208 233884 282220
rect 233936 282208 233942 282260
rect 317690 282208 317696 282260
rect 317748 282248 317754 282260
rect 475378 282248 475384 282260
rect 317748 282220 475384 282248
rect 317748 282208 317754 282220
rect 475378 282208 475384 282220
rect 475436 282208 475442 282260
rect 20714 282140 20720 282192
rect 20772 282180 20778 282192
rect 233418 282180 233424 282192
rect 20772 282152 233424 282180
rect 20772 282140 20778 282152
rect 233418 282140 233424 282152
rect 233476 282140 233482 282192
rect 335630 282140 335636 282192
rect 335688 282180 335694 282192
rect 574738 282180 574744 282192
rect 335688 282152 574744 282180
rect 335688 282140 335694 282152
rect 574738 282140 574744 282152
rect 574796 282140 574802 282192
rect 312170 280916 312176 280968
rect 312228 280956 312234 280968
rect 452654 280956 452660 280968
rect 312228 280928 452660 280956
rect 312228 280916 312234 280928
rect 452654 280916 452660 280928
rect 452712 280916 452718 280968
rect 93118 280848 93124 280900
rect 93176 280888 93182 280900
rect 245838 280888 245844 280900
rect 93176 280860 245844 280888
rect 93176 280848 93182 280860
rect 245838 280848 245844 280860
rect 245896 280848 245902 280900
rect 319070 280848 319076 280900
rect 319128 280888 319134 280900
rect 488534 280888 488540 280900
rect 319128 280860 488540 280888
rect 319128 280848 319134 280860
rect 488534 280848 488540 280860
rect 488592 280848 488598 280900
rect 26234 280780 26240 280832
rect 26292 280820 26298 280832
rect 234890 280820 234896 280832
rect 26292 280792 234896 280820
rect 26292 280780 26298 280792
rect 234890 280780 234896 280792
rect 234948 280780 234954 280832
rect 334066 280780 334072 280832
rect 334124 280820 334130 280832
rect 567194 280820 567200 280832
rect 334124 280792 567200 280820
rect 334124 280780 334130 280792
rect 567194 280780 567200 280792
rect 567252 280780 567258 280832
rect 314930 279556 314936 279608
rect 314988 279596 314994 279608
rect 460934 279596 460940 279608
rect 314988 279568 460940 279596
rect 314988 279556 314994 279568
rect 460934 279556 460940 279568
rect 460992 279556 460998 279608
rect 88334 279488 88340 279540
rect 88392 279528 88398 279540
rect 245746 279528 245752 279540
rect 88392 279500 245752 279528
rect 88392 279488 88398 279500
rect 245746 279488 245752 279500
rect 245804 279488 245810 279540
rect 315022 279488 315028 279540
rect 315080 279528 315086 279540
rect 463694 279528 463700 279540
rect 315080 279500 463700 279528
rect 315080 279488 315086 279500
rect 463694 279488 463700 279500
rect 463752 279488 463758 279540
rect 28994 279420 29000 279472
rect 29052 279460 29058 279472
rect 234798 279460 234804 279472
rect 29052 279432 234804 279460
rect 29052 279420 29058 279432
rect 234798 279420 234804 279432
rect 234856 279420 234862 279472
rect 320450 279420 320456 279472
rect 320508 279460 320514 279472
rect 491294 279460 491300 279472
rect 320508 279432 491300 279460
rect 320508 279420 320514 279432
rect 491294 279420 491300 279432
rect 491352 279420 491358 279472
rect 318978 278060 318984 278112
rect 319036 278100 319042 278112
rect 485774 278100 485780 278112
rect 319036 278072 485780 278100
rect 319036 278060 319042 278072
rect 485774 278060 485780 278072
rect 485832 278060 485838 278112
rect 35158 277992 35164 278044
rect 35216 278032 35222 278044
rect 236178 278032 236184 278044
rect 35216 278004 236184 278032
rect 35216 277992 35222 278004
rect 236178 277992 236184 278004
rect 236236 277992 236242 278044
rect 323210 277992 323216 278044
rect 323268 278032 323274 278044
rect 506474 278032 506480 278044
rect 323268 278004 506480 278032
rect 323268 277992 323274 278004
rect 506474 277992 506480 278004
rect 506532 277992 506538 278044
rect 317598 276700 317604 276752
rect 317656 276740 317662 276752
rect 477494 276740 477500 276752
rect 317656 276712 477500 276740
rect 317656 276700 317662 276712
rect 477494 276700 477500 276712
rect 477552 276700 477558 276752
rect 35986 276632 35992 276684
rect 36044 276672 36050 276684
rect 236086 276672 236092 276684
rect 36044 276644 236092 276672
rect 36044 276632 36050 276644
rect 236086 276632 236092 276644
rect 236144 276632 236150 276684
rect 324590 276632 324596 276684
rect 324648 276672 324654 276684
rect 509878 276672 509884 276684
rect 324648 276644 509884 276672
rect 324648 276632 324654 276644
rect 509878 276632 509884 276644
rect 509936 276632 509942 276684
rect 320358 275340 320364 275392
rect 320416 275380 320422 275392
rect 492674 275380 492680 275392
rect 320416 275352 492680 275380
rect 320416 275340 320422 275352
rect 492674 275340 492680 275352
rect 492732 275340 492738 275392
rect 44174 275272 44180 275324
rect 44232 275312 44238 275324
rect 237558 275312 237564 275324
rect 44232 275284 237564 275312
rect 44232 275272 44238 275284
rect 237558 275272 237564 275284
rect 237616 275272 237622 275324
rect 325786 275272 325792 275324
rect 325844 275312 325850 275324
rect 526530 275312 526536 275324
rect 325844 275284 526536 275312
rect 325844 275272 325850 275284
rect 526530 275272 526536 275284
rect 526588 275272 526594 275324
rect 310606 274048 310612 274100
rect 310664 274088 310670 274100
rect 444374 274088 444380 274100
rect 310664 274060 444380 274088
rect 310664 274048 310670 274060
rect 444374 274048 444380 274060
rect 444432 274048 444438 274100
rect 321738 273980 321744 274032
rect 321796 274020 321802 274032
rect 499574 274020 499580 274032
rect 321796 273992 499580 274020
rect 321796 273980 321802 273992
rect 499574 273980 499580 273992
rect 499632 273980 499638 274032
rect 14458 273912 14464 273964
rect 14516 273952 14522 273964
rect 230658 273952 230664 273964
rect 14516 273924 230664 273952
rect 14516 273912 14522 273924
rect 230658 273912 230664 273924
rect 230716 273912 230722 273964
rect 327350 273912 327356 273964
rect 327408 273952 327414 273964
rect 531314 273952 531320 273964
rect 327408 273924 531320 273952
rect 327408 273912 327414 273924
rect 531314 273912 531320 273924
rect 531372 273912 531378 273964
rect 367738 273164 367744 273216
rect 367796 273204 367802 273216
rect 579890 273204 579896 273216
rect 367796 273176 579896 273204
rect 367796 273164 367802 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 48314 272484 48320 272536
rect 48372 272524 48378 272536
rect 239030 272524 239036 272536
rect 48372 272496 239036 272524
rect 48372 272484 48378 272496
rect 239030 272484 239036 272496
rect 239088 272484 239094 272536
rect 324498 272484 324504 272536
rect 324556 272524 324562 272536
rect 517514 272524 517520 272536
rect 324556 272496 517520 272524
rect 324556 272484 324562 272496
rect 517514 272484 517520 272496
rect 517572 272484 517578 272536
rect 312078 271260 312084 271312
rect 312136 271300 312142 271312
rect 446398 271300 446404 271312
rect 312136 271272 446404 271300
rect 312136 271260 312142 271272
rect 446398 271260 446404 271272
rect 446456 271260 446462 271312
rect 323118 271192 323124 271244
rect 323176 271232 323182 271244
rect 510614 271232 510620 271244
rect 323176 271204 510620 271232
rect 323176 271192 323182 271204
rect 510614 271192 510620 271204
rect 510672 271192 510678 271244
rect 52454 271124 52460 271176
rect 52512 271164 52518 271176
rect 238938 271164 238944 271176
rect 52512 271136 238944 271164
rect 52512 271124 52518 271136
rect 238938 271124 238944 271136
rect 238996 271124 239002 271176
rect 328638 271124 328644 271176
rect 328696 271164 328702 271176
rect 540238 271164 540244 271176
rect 328696 271136 540244 271164
rect 328696 271124 328702 271136
rect 540238 271124 540244 271136
rect 540296 271124 540302 271176
rect 313366 269900 313372 269952
rect 313424 269940 313430 269952
rect 453298 269940 453304 269952
rect 313424 269912 453304 269940
rect 313424 269900 313430 269912
rect 453298 269900 453304 269912
rect 453356 269900 453362 269952
rect 325694 269832 325700 269884
rect 325752 269872 325758 269884
rect 524414 269872 524420 269884
rect 325752 269844 524420 269872
rect 325752 269832 325758 269844
rect 524414 269832 524420 269844
rect 524472 269832 524478 269884
rect 57238 269764 57244 269816
rect 57296 269804 57302 269816
rect 240226 269804 240232 269816
rect 57296 269776 240232 269804
rect 57296 269764 57302 269776
rect 240226 269764 240232 269776
rect 240284 269764 240290 269816
rect 329926 269764 329932 269816
rect 329984 269804 329990 269816
rect 542998 269804 543004 269816
rect 329984 269776 543004 269804
rect 329984 269764 329990 269776
rect 542998 269764 543004 269776
rect 543056 269764 543062 269816
rect 314838 268472 314844 268524
rect 314896 268512 314902 268524
rect 460198 268512 460204 268524
rect 314896 268484 460204 268512
rect 314896 268472 314902 268484
rect 460198 268472 460204 268484
rect 460256 268472 460262 268524
rect 327258 268404 327264 268456
rect 327316 268444 327322 268456
rect 531406 268444 531412 268456
rect 327316 268416 531412 268444
rect 327316 268404 327322 268416
rect 531406 268404 531412 268416
rect 531464 268404 531470 268456
rect 59354 268336 59360 268388
rect 59412 268376 59418 268388
rect 240502 268376 240508 268388
rect 59412 268348 240508 268376
rect 59412 268336 59418 268348
rect 240502 268336 240508 268348
rect 240560 268336 240566 268388
rect 331490 268336 331496 268388
rect 331548 268376 331554 268388
rect 552014 268376 552020 268388
rect 331548 268348 552020 268376
rect 331548 268336 331554 268348
rect 552014 268336 552020 268348
rect 552072 268336 552078 268388
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 224218 267696 224224 267708
rect 3016 267668 224224 267696
rect 3016 267656 3022 267668
rect 224218 267656 224224 267668
rect 224276 267656 224282 267708
rect 314746 267180 314752 267232
rect 314804 267220 314810 267232
rect 464338 267220 464344 267232
rect 314804 267192 464344 267220
rect 314804 267180 314810 267192
rect 464338 267180 464344 267192
rect 464396 267180 464402 267232
rect 328546 267112 328552 267164
rect 328604 267152 328610 267164
rect 542354 267152 542360 267164
rect 328604 267124 542360 267152
rect 328604 267112 328610 267124
rect 542354 267112 542360 267124
rect 542412 267112 542418 267164
rect 331398 267044 331404 267096
rect 331456 267084 331462 267096
rect 556154 267084 556160 267096
rect 331456 267056 556160 267084
rect 331456 267044 331462 267056
rect 556154 267044 556160 267056
rect 556212 267044 556218 267096
rect 99282 266976 99288 267028
rect 99340 267016 99346 267028
rect 335538 267016 335544 267028
rect 99340 266988 335544 267016
rect 99340 266976 99346 266988
rect 335538 266976 335544 266988
rect 335596 266976 335602 267028
rect 238202 265820 238208 265872
rect 238260 265860 238266 265872
rect 350994 265860 351000 265872
rect 238260 265832 351000 265860
rect 238260 265820 238266 265832
rect 350994 265820 351000 265832
rect 351052 265820 351058 265872
rect 317506 265752 317512 265804
rect 317564 265792 317570 265804
rect 481634 265792 481640 265804
rect 317564 265764 481640 265792
rect 317564 265752 317570 265764
rect 481634 265752 481640 265764
rect 481692 265752 481698 265804
rect 329834 265684 329840 265736
rect 329892 265724 329898 265736
rect 546494 265724 546500 265736
rect 329892 265696 546500 265724
rect 329892 265684 329898 265696
rect 546494 265684 546500 265696
rect 546552 265684 546558 265736
rect 66254 265616 66260 265668
rect 66312 265656 66318 265668
rect 241882 265656 241888 265668
rect 66312 265628 241888 265656
rect 66312 265616 66318 265628
rect 241882 265616 241888 265628
rect 241940 265616 241946 265668
rect 332778 265616 332784 265668
rect 332836 265656 332842 265668
rect 560938 265656 560944 265668
rect 332836 265628 560944 265656
rect 332836 265616 332842 265628
rect 560938 265616 560944 265628
rect 560996 265616 561002 265668
rect 317414 264256 317420 264308
rect 317472 264296 317478 264308
rect 481726 264296 481732 264308
rect 317472 264268 481732 264296
rect 317472 264256 317478 264268
rect 481726 264256 481732 264268
rect 481784 264256 481790 264308
rect 75178 264188 75184 264240
rect 75236 264228 75242 264240
rect 243354 264228 243360 264240
rect 75236 264200 243360 264228
rect 75236 264188 75242 264200
rect 243354 264188 243360 264200
rect 243412 264188 243418 264240
rect 318886 264188 318892 264240
rect 318944 264228 318950 264240
rect 484394 264228 484400 264240
rect 318944 264200 484400 264228
rect 318944 264188 318950 264200
rect 484394 264188 484400 264200
rect 484452 264188 484458 264240
rect 77386 262896 77392 262948
rect 77444 262936 77450 262948
rect 243262 262936 243268 262948
rect 77444 262908 243268 262936
rect 77444 262896 77450 262908
rect 243262 262896 243268 262908
rect 243320 262896 243326 262948
rect 318794 262896 318800 262948
rect 318852 262936 318858 262948
rect 490006 262936 490012 262948
rect 318852 262908 490012 262936
rect 318852 262896 318858 262908
rect 490006 262896 490012 262908
rect 490064 262896 490070 262948
rect 4154 262828 4160 262880
rect 4212 262868 4218 262880
rect 230934 262868 230940 262880
rect 4212 262840 230940 262868
rect 4212 262828 4218 262840
rect 230934 262828 230940 262840
rect 230992 262828 230998 262880
rect 320266 262828 320272 262880
rect 320324 262868 320330 262880
rect 495434 262868 495440 262880
rect 320324 262840 495440 262868
rect 320324 262828 320330 262840
rect 495434 262828 495440 262840
rect 495492 262828 495498 262880
rect 84194 261536 84200 261588
rect 84252 261576 84258 261588
rect 244458 261576 244464 261588
rect 84252 261548 244464 261576
rect 84252 261536 84258 261548
rect 244458 261536 244464 261548
rect 244516 261536 244522 261588
rect 320174 261536 320180 261588
rect 320232 261576 320238 261588
rect 496078 261576 496084 261588
rect 320232 261548 496084 261576
rect 320232 261536 320238 261548
rect 496078 261536 496084 261548
rect 496136 261536 496142 261588
rect 31754 261468 31760 261520
rect 31812 261508 31818 261520
rect 234706 261508 234712 261520
rect 31812 261480 234712 261508
rect 31812 261468 31818 261480
rect 234706 261468 234712 261480
rect 234764 261468 234770 261520
rect 321646 261468 321652 261520
rect 321704 261508 321710 261520
rect 502334 261508 502340 261520
rect 321704 261480 502340 261508
rect 321704 261468 321710 261480
rect 502334 261468 502340 261480
rect 502392 261468 502398 261520
rect 311986 260244 311992 260296
rect 312044 260284 312050 260296
rect 445754 260284 445760 260296
rect 312044 260256 445760 260284
rect 312044 260244 312050 260256
rect 445754 260244 445760 260256
rect 445812 260244 445818 260296
rect 91094 260176 91100 260228
rect 91152 260216 91158 260228
rect 246114 260216 246120 260228
rect 91152 260188 246120 260216
rect 91152 260176 91158 260188
rect 246114 260176 246120 260188
rect 246172 260176 246178 260228
rect 364978 260176 364984 260228
rect 365036 260216 365042 260228
rect 580442 260216 580448 260228
rect 365036 260188 580448 260216
rect 365036 260176 365042 260188
rect 580442 260176 580448 260188
rect 580500 260176 580506 260228
rect 13814 260108 13820 260160
rect 13872 260148 13878 260160
rect 231946 260148 231952 260160
rect 13872 260120 231952 260148
rect 13872 260108 13878 260120
rect 231946 260108 231952 260120
rect 232004 260108 232010 260160
rect 332686 260108 332692 260160
rect 332744 260148 332750 260160
rect 564526 260148 564532 260160
rect 332744 260120 564532 260148
rect 332744 260108 332750 260120
rect 564526 260108 564532 260120
rect 564584 260108 564590 260160
rect 314654 258816 314660 258868
rect 314712 258856 314718 258868
rect 466454 258856 466460 258868
rect 314712 258828 466460 258856
rect 314712 258816 314718 258828
rect 466454 258816 466460 258828
rect 466512 258816 466518 258868
rect 319438 258748 319444 258800
rect 319496 258788 319502 258800
rect 471974 258788 471980 258800
rect 319496 258760 471980 258788
rect 319496 258748 319502 258760
rect 471974 258748 471980 258760
rect 472032 258748 472038 258800
rect 63494 258680 63500 258732
rect 63552 258720 63558 258732
rect 236638 258720 236644 258732
rect 63552 258692 236644 258720
rect 63552 258680 63558 258692
rect 236638 258680 236644 258692
rect 236696 258680 236702 258732
rect 363598 258680 363604 258732
rect 363656 258720 363662 258732
rect 580350 258720 580356 258732
rect 363656 258692 580356 258720
rect 363656 258680 363662 258692
rect 580350 258680 580356 258692
rect 580408 258680 580414 258732
rect 373258 257320 373264 257372
rect 373316 257360 373322 257372
rect 581086 257360 581092 257372
rect 373316 257332 581092 257360
rect 373316 257320 373322 257332
rect 581086 257320 581092 257332
rect 581144 257320 581150 257372
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 225598 255252 225604 255264
rect 3200 255224 225604 255252
rect 3200 255212 3206 255224
rect 225598 255212 225604 255224
rect 225656 255212 225662 255264
rect 299382 254736 299388 254788
rect 299440 254776 299446 254788
rect 336918 254776 336924 254788
rect 299440 254748 336924 254776
rect 299440 254736 299446 254748
rect 336918 254736 336924 254748
rect 336976 254736 336982 254788
rect 297542 254668 297548 254720
rect 297600 254708 297606 254720
rect 342622 254708 342628 254720
rect 297600 254680 342628 254708
rect 297600 254668 297606 254680
rect 342622 254668 342628 254680
rect 342680 254668 342686 254720
rect 316034 254600 316040 254652
rect 316092 254640 316098 254652
rect 467834 254640 467840 254652
rect 316092 254612 467840 254640
rect 316092 254600 316098 254612
rect 467834 254600 467840 254612
rect 467892 254600 467898 254652
rect 316126 254532 316132 254584
rect 316184 254572 316190 254584
rect 474734 254572 474740 254584
rect 316184 254544 474740 254572
rect 316184 254532 316190 254544
rect 474734 254532 474740 254544
rect 474792 254532 474798 254584
rect 297634 253444 297640 253496
rect 297692 253484 297698 253496
rect 339586 253484 339592 253496
rect 297692 253456 339592 253484
rect 297692 253444 297698 253456
rect 339586 253444 339592 253456
rect 339644 253444 339650 253496
rect 297174 253376 297180 253428
rect 297232 253416 297238 253428
rect 343818 253416 343824 253428
rect 297232 253388 343824 253416
rect 297232 253376 297238 253388
rect 343818 253376 343824 253388
rect 343876 253376 343882 253428
rect 309502 253308 309508 253360
rect 309560 253348 309566 253360
rect 436738 253348 436744 253360
rect 309560 253320 436744 253348
rect 309560 253308 309566 253320
rect 436738 253308 436744 253320
rect 436796 253308 436802 253360
rect 333974 253240 333980 253292
rect 334032 253280 334038 253292
rect 571334 253280 571340 253292
rect 334032 253252 571340 253280
rect 334032 253240 334038 253252
rect 571334 253240 571340 253252
rect 571392 253240 571398 253292
rect 27706 253172 27712 253224
rect 27764 253212 27770 253224
rect 235074 253212 235080 253224
rect 27764 253184 235080 253212
rect 27764 253172 27770 253184
rect 235074 253172 235080 253184
rect 235132 253172 235138 253224
rect 335446 253172 335452 253224
rect 335504 253212 335510 253224
rect 574094 253212 574100 253224
rect 335504 253184 574100 253212
rect 335504 253172 335510 253184
rect 574094 253172 574100 253184
rect 574152 253172 574158 253224
rect 297450 252016 297456 252068
rect 297508 252056 297514 252068
rect 341150 252056 341156 252068
rect 297508 252028 341156 252056
rect 297508 252016 297514 252028
rect 341150 252016 341156 252028
rect 341208 252016 341214 252068
rect 321554 251948 321560 252000
rect 321612 251988 321618 252000
rect 503714 251988 503720 252000
rect 321612 251960 503720 251988
rect 321612 251948 321618 251960
rect 503714 251948 503720 251960
rect 503772 251948 503778 252000
rect 323026 251880 323032 251932
rect 323084 251920 323090 251932
rect 506566 251920 506572 251932
rect 323084 251892 506572 251920
rect 323084 251880 323090 251892
rect 506566 251880 506572 251892
rect 506624 251880 506630 251932
rect 12434 251812 12440 251864
rect 12492 251852 12498 251864
rect 232222 251852 232228 251864
rect 12492 251824 232228 251852
rect 12492 251812 12498 251824
rect 232222 251812 232228 251824
rect 232280 251812 232286 251864
rect 332594 251812 332600 251864
rect 332652 251852 332658 251864
rect 560294 251852 560300 251864
rect 332652 251824 560300 251852
rect 332652 251812 332658 251824
rect 560294 251812 560300 251824
rect 560352 251812 560358 251864
rect 238386 250588 238392 250640
rect 238444 250628 238450 250640
rect 355134 250628 355140 250640
rect 238444 250600 355140 250628
rect 238444 250588 238450 250600
rect 355134 250588 355140 250600
rect 355192 250588 355198 250640
rect 310514 250520 310520 250572
rect 310572 250560 310578 250572
rect 441614 250560 441620 250572
rect 310572 250532 441620 250560
rect 310572 250520 310578 250532
rect 441614 250520 441620 250532
rect 441672 250520 441678 250572
rect 39390 250452 39396 250504
rect 39448 250492 39454 250504
rect 236362 250492 236368 250504
rect 39448 250464 236368 250492
rect 39448 250452 39454 250464
rect 236362 250452 236368 250464
rect 236420 250452 236426 250504
rect 324406 250452 324412 250504
rect 324464 250492 324470 250504
rect 514110 250492 514116 250504
rect 324464 250464 514116 250492
rect 324464 250452 324470 250464
rect 514110 250452 514116 250464
rect 514168 250452 514174 250504
rect 313274 249092 313280 249144
rect 313332 249132 313338 249144
rect 459554 249132 459560 249144
rect 313332 249104 459560 249132
rect 313332 249092 313338 249104
rect 459554 249092 459560 249104
rect 459612 249092 459618 249144
rect 4798 249024 4804 249076
rect 4856 249064 4862 249076
rect 229186 249064 229192 249076
rect 4856 249036 229192 249064
rect 4856 249024 4862 249036
rect 229186 249024 229192 249036
rect 229244 249024 229250 249076
rect 331306 249024 331312 249076
rect 331364 249064 331370 249076
rect 553394 249064 553400 249076
rect 331364 249036 553400 249064
rect 331364 249024 331370 249036
rect 553394 249024 553400 249036
rect 553452 249024 553458 249076
rect 289354 248344 289360 248396
rect 289412 248384 289418 248396
rect 303798 248384 303804 248396
rect 289412 248356 303804 248384
rect 289412 248344 289418 248356
rect 303798 248344 303804 248356
rect 303856 248344 303862 248396
rect 298646 248276 298652 248328
rect 298704 248316 298710 248328
rect 345474 248316 345480 248328
rect 298704 248288 345480 248316
rect 298704 248276 298710 248288
rect 345474 248276 345480 248288
rect 345532 248276 345538 248328
rect 296530 248208 296536 248260
rect 296588 248248 296594 248260
rect 344094 248248 344100 248260
rect 296588 248220 344100 248248
rect 296588 248208 296594 248220
rect 344094 248208 344100 248220
rect 344152 248208 344158 248260
rect 292298 248140 292304 248192
rect 292356 248180 292362 248192
rect 345198 248180 345204 248192
rect 292356 248152 345204 248180
rect 292356 248140 292362 248152
rect 345198 248140 345204 248152
rect 345256 248140 345262 248192
rect 358998 248140 359004 248192
rect 359056 248180 359062 248192
rect 438210 248180 438216 248192
rect 359056 248152 438216 248180
rect 359056 248140 359062 248152
rect 438210 248140 438216 248152
rect 438268 248140 438274 248192
rect 293678 248072 293684 248124
rect 293736 248112 293742 248124
rect 350902 248112 350908 248124
rect 293736 248084 350908 248112
rect 293736 248072 293742 248084
rect 350902 248072 350908 248084
rect 350960 248072 350966 248124
rect 356422 248072 356428 248124
rect 356480 248112 356486 248124
rect 436922 248112 436928 248124
rect 356480 248084 436928 248112
rect 356480 248072 356486 248084
rect 436922 248072 436928 248084
rect 436980 248072 436986 248124
rect 290734 248004 290740 248056
rect 290792 248044 290798 248056
rect 347958 248044 347964 248056
rect 290792 248016 347964 248044
rect 290792 248004 290798 248016
rect 347958 248004 347964 248016
rect 348016 248004 348022 248056
rect 357710 248004 357716 248056
rect 357768 248044 357774 248056
rect 440510 248044 440516 248056
rect 357768 248016 440516 248044
rect 357768 248004 357774 248016
rect 440510 248004 440516 248016
rect 440568 248004 440574 248056
rect 288158 247936 288164 247988
rect 288216 247976 288222 247988
rect 348326 247976 348332 247988
rect 288216 247948 348332 247976
rect 288216 247936 288222 247948
rect 348326 247936 348332 247948
rect 348384 247936 348390 247988
rect 359274 247936 359280 247988
rect 359332 247976 359338 247988
rect 441706 247976 441712 247988
rect 359332 247948 441712 247976
rect 359332 247936 359338 247948
rect 441706 247936 441712 247948
rect 441764 247936 441770 247988
rect 285582 247868 285588 247920
rect 285640 247908 285646 247920
rect 304074 247908 304080 247920
rect 285640 247880 304080 247908
rect 285640 247868 285646 247880
rect 304074 247868 304080 247880
rect 304132 247868 304138 247920
rect 308214 247868 308220 247920
rect 308272 247908 308278 247920
rect 437566 247908 437572 247920
rect 308272 247880 437572 247908
rect 308272 247868 308278 247880
rect 437566 247868 437572 247880
rect 437624 247868 437630 247920
rect 287974 247800 287980 247852
rect 288032 247840 288038 247852
rect 305362 247840 305368 247852
rect 288032 247812 305368 247840
rect 288032 247800 288038 247812
rect 305362 247800 305368 247812
rect 305420 247800 305426 247852
rect 308122 247800 308128 247852
rect 308180 247840 308186 247852
rect 438854 247840 438860 247852
rect 308180 247812 438860 247840
rect 308180 247800 308186 247812
rect 438854 247800 438860 247812
rect 438912 247800 438918 247852
rect 287882 247732 287888 247784
rect 287940 247772 287946 247784
rect 303982 247772 303988 247784
rect 287940 247744 303988 247772
rect 287940 247732 287946 247744
rect 303982 247732 303988 247744
rect 304040 247732 304046 247784
rect 322934 247732 322940 247784
rect 322992 247772 322998 247784
rect 509234 247772 509240 247784
rect 322992 247744 509240 247772
rect 322992 247732 322998 247744
rect 509234 247732 509240 247744
rect 509292 247732 509298 247784
rect 3694 247664 3700 247716
rect 3752 247704 3758 247716
rect 228358 247704 228364 247716
rect 3752 247676 228364 247704
rect 3752 247664 3758 247676
rect 228358 247664 228364 247676
rect 228416 247664 228422 247716
rect 289170 247664 289176 247716
rect 289228 247704 289234 247716
rect 305270 247704 305276 247716
rect 289228 247676 305276 247704
rect 289228 247664 289234 247676
rect 305270 247664 305276 247676
rect 305328 247664 305334 247716
rect 327166 247664 327172 247716
rect 327224 247704 327230 247716
rect 528554 247704 528560 247716
rect 327224 247676 528560 247704
rect 327224 247664 327230 247676
rect 528554 247664 528560 247676
rect 528612 247664 528618 247716
rect 284754 247596 284760 247648
rect 284812 247636 284818 247648
rect 305178 247636 305184 247648
rect 284812 247608 305184 247636
rect 284812 247596 284818 247608
rect 305178 247596 305184 247608
rect 305236 247596 305242 247648
rect 286962 247528 286968 247580
rect 287020 247568 287026 247580
rect 303890 247568 303896 247580
rect 287020 247540 303896 247568
rect 287020 247528 287026 247540
rect 303890 247528 303896 247540
rect 303948 247528 303954 247580
rect 286686 247460 286692 247512
rect 286744 247500 286750 247512
rect 305454 247500 305460 247512
rect 286744 247472 305460 247500
rect 286744 247460 286750 247472
rect 305454 247460 305460 247472
rect 305512 247460 305518 247512
rect 300762 246644 300768 246696
rect 300820 246684 300826 246696
rect 346486 246684 346492 246696
rect 300820 246656 346492 246684
rect 300820 246644 300826 246656
rect 346486 246644 346492 246656
rect 346544 246644 346550 246696
rect 297266 246576 297272 246628
rect 297324 246616 297330 246628
rect 349430 246616 349436 246628
rect 297324 246588 349436 246616
rect 297324 246576 297330 246588
rect 349430 246576 349436 246588
rect 349488 246576 349494 246628
rect 289630 246508 289636 246560
rect 289688 246548 289694 246560
rect 349246 246548 349252 246560
rect 289688 246520 349252 246548
rect 289688 246508 289694 246520
rect 349246 246508 349252 246520
rect 349304 246508 349310 246560
rect 311894 246440 311900 246492
rect 311952 246480 311958 246492
rect 448606 246480 448612 246492
rect 311952 246452 448612 246480
rect 311952 246440 311958 246452
rect 448606 246440 448612 246452
rect 448664 246440 448670 246492
rect 327074 246372 327080 246424
rect 327132 246412 327138 246424
rect 534074 246412 534080 246424
rect 327132 246384 534080 246412
rect 327132 246372 327138 246384
rect 534074 246372 534080 246384
rect 534132 246372 534138 246424
rect 7650 246304 7656 246356
rect 7708 246344 7714 246356
rect 230842 246344 230848 246356
rect 7708 246316 230848 246344
rect 7708 246304 7714 246316
rect 230842 246304 230848 246316
rect 230900 246304 230906 246356
rect 331214 246304 331220 246356
rect 331272 246344 331278 246356
rect 556246 246344 556252 246356
rect 331272 246316 556252 246344
rect 331272 246304 331278 246316
rect 556246 246304 556252 246316
rect 556304 246304 556310 246356
rect 292114 245556 292120 245608
rect 292172 245596 292178 245608
rect 302326 245596 302332 245608
rect 292172 245568 302332 245596
rect 292172 245556 292178 245568
rect 302326 245556 302332 245568
rect 302384 245556 302390 245608
rect 357618 245556 357624 245608
rect 357676 245596 357682 245608
rect 440602 245596 440608 245608
rect 357676 245568 440608 245596
rect 357676 245556 357682 245568
rect 440602 245556 440608 245568
rect 440660 245556 440666 245608
rect 307938 245488 307944 245540
rect 307996 245528 308002 245540
rect 437658 245528 437664 245540
rect 307996 245500 437664 245528
rect 307996 245488 308002 245500
rect 437658 245488 437664 245500
rect 437716 245488 437722 245540
rect 291746 245420 291752 245472
rect 291804 245460 291810 245472
rect 306650 245460 306656 245472
rect 291804 245432 306656 245460
rect 291804 245420 291810 245432
rect 306650 245420 306656 245432
rect 306708 245420 306714 245472
rect 309226 245420 309232 245472
rect 309284 245460 309290 245472
rect 439038 245460 439044 245472
rect 309284 245432 439044 245460
rect 309284 245420 309290 245432
rect 439038 245420 439044 245432
rect 439096 245420 439102 245472
rect 293402 245352 293408 245404
rect 293460 245392 293466 245404
rect 304994 245392 305000 245404
rect 293460 245364 305000 245392
rect 293460 245352 293466 245364
rect 304994 245352 305000 245364
rect 305052 245352 305058 245404
rect 307846 245352 307852 245404
rect 307904 245392 307910 245404
rect 437842 245392 437848 245404
rect 307904 245364 437848 245392
rect 307904 245352 307910 245364
rect 437842 245352 437848 245364
rect 437900 245352 437906 245404
rect 295058 245284 295064 245336
rect 295116 245324 295122 245336
rect 305086 245324 305092 245336
rect 295116 245296 305092 245324
rect 295116 245284 295122 245296
rect 305086 245284 305092 245296
rect 305144 245284 305150 245336
rect 308030 245284 308036 245336
rect 308088 245324 308094 245336
rect 439130 245324 439136 245336
rect 308088 245296 439136 245324
rect 308088 245284 308094 245296
rect 439130 245284 439136 245296
rect 439188 245284 439194 245336
rect 293770 245216 293776 245268
rect 293828 245256 293834 245268
rect 302418 245256 302424 245268
rect 293828 245228 302424 245256
rect 293828 245216 293834 245228
rect 302418 245216 302424 245228
rect 302476 245216 302482 245268
rect 306742 245216 306748 245268
rect 306800 245256 306806 245268
rect 437934 245256 437940 245268
rect 306800 245228 437940 245256
rect 306800 245216 306806 245228
rect 437934 245216 437940 245228
rect 437992 245216 437998 245268
rect 295242 245148 295248 245200
rect 295300 245188 295306 245200
rect 299566 245188 299572 245200
rect 295300 245160 299572 245188
rect 295300 245148 295306 245160
rect 299566 245148 299572 245160
rect 299624 245148 299630 245200
rect 306466 245148 306472 245200
rect 306524 245188 306530 245200
rect 437750 245188 437756 245200
rect 306524 245160 437756 245188
rect 306524 245148 306530 245160
rect 437750 245148 437756 245160
rect 437808 245148 437814 245200
rect 288342 245080 288348 245132
rect 288400 245120 288406 245132
rect 296898 245120 296904 245132
rect 288400 245092 296904 245120
rect 288400 245080 288406 245092
rect 296898 245080 296904 245092
rect 296956 245080 296962 245132
rect 307754 245080 307760 245132
rect 307812 245120 307818 245132
rect 439314 245120 439320 245132
rect 307812 245092 439320 245120
rect 307812 245080 307818 245092
rect 439314 245080 439320 245092
rect 439372 245080 439378 245132
rect 295150 245012 295156 245064
rect 295208 245052 295214 245064
rect 303706 245052 303712 245064
rect 295208 245024 303712 245052
rect 295208 245012 295214 245024
rect 303706 245012 303712 245024
rect 303764 245012 303770 245064
rect 306558 245012 306564 245064
rect 306616 245052 306622 245064
rect 438946 245052 438952 245064
rect 306616 245024 438952 245052
rect 306616 245012 306622 245024
rect 438946 245012 438952 245024
rect 439004 245012 439010 245064
rect 22094 244944 22100 244996
rect 22152 244984 22158 244996
rect 233510 244984 233516 244996
rect 22152 244956 233516 244984
rect 22152 244944 22158 244956
rect 233510 244944 233516 244956
rect 233568 244944 233574 244996
rect 291102 244944 291108 244996
rect 291160 244984 291166 244996
rect 299750 244984 299756 244996
rect 291160 244956 299756 244984
rect 291160 244944 291166 244956
rect 299750 244944 299756 244956
rect 299808 244944 299814 244996
rect 306374 244944 306380 244996
rect 306432 244984 306438 244996
rect 439222 244984 439228 244996
rect 306432 244956 439228 244984
rect 306432 244944 306438 244956
rect 439222 244944 439228 244956
rect 439280 244944 439286 244996
rect 17954 244876 17960 244928
rect 18012 244916 18018 244928
rect 233326 244916 233332 244928
rect 18012 244888 233332 244916
rect 18012 244876 18018 244888
rect 233326 244876 233332 244888
rect 233384 244876 233390 244928
rect 291010 244876 291016 244928
rect 291068 244916 291074 244928
rect 300854 244916 300860 244928
rect 291068 244888 300860 244916
rect 291068 244876 291074 244888
rect 300854 244876 300860 244888
rect 300912 244876 300918 244928
rect 324314 244876 324320 244928
rect 324372 244916 324378 244928
rect 520274 244916 520280 244928
rect 324372 244888 520280 244916
rect 324372 244876 324378 244888
rect 520274 244876 520280 244888
rect 520332 244876 520338 244928
rect 298922 244808 298928 244860
rect 298980 244848 298986 244860
rect 339862 244848 339868 244860
rect 298980 244820 339868 244848
rect 298980 244808 298986 244820
rect 339862 244808 339868 244820
rect 339920 244808 339926 244860
rect 359182 244808 359188 244860
rect 359240 244848 359246 244860
rect 441798 244848 441804 244860
rect 359240 244820 441804 244848
rect 359240 244808 359246 244820
rect 441798 244808 441804 244820
rect 441856 244808 441862 244860
rect 297726 244740 297732 244792
rect 297784 244780 297790 244792
rect 335354 244780 335360 244792
rect 297784 244752 335360 244780
rect 297784 244740 297790 244752
rect 335354 244740 335360 244752
rect 335412 244740 335418 244792
rect 356514 244740 356520 244792
rect 356572 244780 356578 244792
rect 438302 244780 438308 244792
rect 356572 244752 438308 244780
rect 356572 244740 356578 244752
rect 438302 244740 438308 244752
rect 438360 244740 438366 244792
rect 290642 244672 290648 244724
rect 290700 244712 290706 244724
rect 306834 244712 306840 244724
rect 290700 244684 306840 244712
rect 290700 244672 290706 244684
rect 306834 244672 306840 244684
rect 306892 244672 306898 244724
rect 360378 244672 360384 244724
rect 360436 244712 360442 244724
rect 439682 244712 439688 244724
rect 360436 244684 439688 244712
rect 360436 244672 360442 244684
rect 439682 244672 439688 244684
rect 439740 244672 439746 244724
rect 298830 244604 298836 244656
rect 298888 244644 298894 244656
rect 342530 244644 342536 244656
rect 298888 244616 342536 244644
rect 298888 244604 298894 244616
rect 342530 244604 342536 244616
rect 342588 244604 342594 244656
rect 97902 244332 97908 244384
rect 97960 244372 97966 244384
rect 297174 244372 297180 244384
rect 97960 244344 297180 244372
rect 97960 244332 97966 244344
rect 297174 244332 297180 244344
rect 297232 244372 297238 244384
rect 297358 244372 297364 244384
rect 297232 244344 297364 244372
rect 297232 244332 297238 244344
rect 297358 244332 297364 244344
rect 297416 244332 297422 244384
rect 297818 244332 297824 244384
rect 297876 244372 297882 244384
rect 303614 244372 303620 244384
rect 297876 244344 303620 244372
rect 297876 244332 297882 244344
rect 303614 244332 303620 244344
rect 303672 244332 303678 244384
rect 3602 244264 3608 244316
rect 3660 244304 3666 244316
rect 299106 244304 299112 244316
rect 3660 244276 299112 244304
rect 3660 244264 3666 244276
rect 299106 244264 299112 244276
rect 299164 244264 299170 244316
rect 295058 243924 295064 243976
rect 295116 243964 295122 243976
rect 300762 243964 300768 243976
rect 295116 243936 300768 243964
rect 295116 243924 295122 243936
rect 300762 243924 300768 243936
rect 300820 243924 300826 243976
rect 299014 243856 299020 243908
rect 299072 243896 299078 243908
rect 344002 243896 344008 243908
rect 299072 243868 344008 243896
rect 299072 243856 299078 243868
rect 344002 243856 344008 243868
rect 344060 243856 344066 243908
rect 299106 243788 299112 243840
rect 299164 243828 299170 243840
rect 345382 243828 345388 243840
rect 299164 243800 345388 243828
rect 299164 243788 299170 243800
rect 345382 243788 345388 243800
rect 345440 243788 345446 243840
rect 293770 243720 293776 243772
rect 293828 243760 293834 243772
rect 348050 243760 348056 243772
rect 293828 243732 348056 243760
rect 293828 243720 293834 243732
rect 348050 243720 348056 243732
rect 348108 243720 348114 243772
rect 297818 243652 297824 243704
rect 297876 243692 297882 243704
rect 357894 243692 357900 243704
rect 297876 243664 357900 243692
rect 297876 243652 297882 243664
rect 357894 243652 357900 243664
rect 357952 243652 357958 243704
rect 285214 243584 285220 243636
rect 285272 243624 285278 243636
rect 346854 243624 346860 243636
rect 285272 243596 346860 243624
rect 285272 243584 285278 243596
rect 346854 243584 346860 243596
rect 346912 243584 346918 243636
rect 286686 243516 286692 243568
rect 286744 243556 286750 243568
rect 357802 243556 357808 243568
rect 286744 243528 357808 243556
rect 286744 243516 286750 243528
rect 357802 243516 357808 243528
rect 357860 243516 357866 243568
rect 97810 243380 97816 243432
rect 97868 243420 97874 243432
rect 298646 243420 298652 243432
rect 97868 243392 298652 243420
rect 97868 243380 97874 243392
rect 298646 243380 298652 243392
rect 298704 243380 298710 243432
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 98638 241448 98644 241460
rect 3292 241420 98644 241448
rect 3292 241408 3298 241420
rect 98638 241408 98644 241420
rect 98696 241408 98702 241460
rect 3142 215228 3148 215280
rect 3200 215268 3206 215280
rect 93210 215268 93216 215280
rect 3200 215240 93216 215268
rect 3200 215228 3206 215240
rect 93210 215228 93216 215240
rect 93268 215228 93274 215280
rect 293678 197276 293684 197328
rect 293736 197316 293742 197328
rect 297174 197316 297180 197328
rect 293736 197288 297180 197316
rect 293736 197276 293742 197288
rect 297174 197276 297180 197288
rect 297232 197276 297238 197328
rect 297266 196392 297272 196444
rect 297324 196432 297330 196444
rect 298554 196432 298560 196444
rect 297324 196404 298560 196432
rect 297324 196392 297330 196404
rect 298554 196392 298560 196404
rect 298612 196392 298618 196444
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 95970 189020 95976 189032
rect 3200 188992 95976 189020
rect 3200 188980 3206 188992
rect 95970 188980 95976 188992
rect 96028 188980 96034 189032
rect 285122 171028 285128 171080
rect 285180 171068 285186 171080
rect 298002 171068 298008 171080
rect 285180 171040 298008 171068
rect 285180 171028 285186 171040
rect 298002 171028 298008 171040
rect 298060 171028 298066 171080
rect 238294 170348 238300 170400
rect 238352 170388 238358 170400
rect 285122 170388 285128 170400
rect 238352 170360 285128 170388
rect 238352 170348 238358 170360
rect 285122 170348 285128 170360
rect 285180 170348 285186 170400
rect 295058 169260 295064 169312
rect 295116 169300 295122 169312
rect 297266 169300 297272 169312
rect 295116 169272 297272 169300
rect 295116 169260 295122 169272
rect 297266 169260 297272 169272
rect 297324 169260 297330 169312
rect 238478 167628 238484 167680
rect 238536 167668 238542 167680
rect 297726 167668 297732 167680
rect 238536 167640 297732 167668
rect 238536 167628 238542 167640
rect 297726 167628 297732 167640
rect 297784 167628 297790 167680
rect 3510 164160 3516 164212
rect 3568 164200 3574 164212
rect 86218 164200 86224 164212
rect 3568 164172 86224 164200
rect 3568 164160 3574 164172
rect 86218 164160 86224 164172
rect 86276 164160 86282 164212
rect 261202 162120 261208 162172
rect 261260 162160 261266 162172
rect 277026 162160 277032 162172
rect 261260 162132 277032 162160
rect 261260 162120 261266 162132
rect 277026 162120 277032 162132
rect 277084 162120 277090 162172
rect 97902 159876 97908 159928
rect 97960 159916 97966 159928
rect 298830 159916 298836 159928
rect 97960 159888 298836 159916
rect 97960 159876 97966 159888
rect 298830 159876 298836 159888
rect 298888 159876 298894 159928
rect 97534 159808 97540 159860
rect 97592 159848 97598 159860
rect 297634 159848 297640 159860
rect 97592 159820 297640 159848
rect 97592 159808 97598 159820
rect 297634 159808 297640 159820
rect 297692 159808 297698 159860
rect 97718 159740 97724 159792
rect 97776 159780 97782 159792
rect 297450 159780 297456 159792
rect 97776 159752 297456 159780
rect 97776 159740 97782 159752
rect 297450 159740 297456 159752
rect 297508 159740 297514 159792
rect 97810 159672 97816 159724
rect 97868 159712 97874 159724
rect 297358 159712 297364 159724
rect 97868 159684 297364 159712
rect 97868 159672 97874 159684
rect 297358 159672 297364 159684
rect 297416 159672 297422 159724
rect 97350 159604 97356 159656
rect 97408 159644 97414 159656
rect 238478 159644 238484 159656
rect 97408 159616 238484 159644
rect 97408 159604 97414 159616
rect 238478 159604 238484 159616
rect 238536 159604 238542 159656
rect 298922 159604 298928 159656
rect 298980 159644 298986 159656
rect 299290 159644 299296 159656
rect 298980 159616 299296 159644
rect 298980 159604 298986 159616
rect 299290 159604 299296 159616
rect 299348 159604 299354 159656
rect 97442 159536 97448 159588
rect 97500 159576 97506 159588
rect 238294 159576 238300 159588
rect 97500 159548 238300 159576
rect 97500 159536 97506 159548
rect 238294 159536 238300 159548
rect 238352 159536 238358 159588
rect 286318 159536 286324 159588
rect 286376 159576 286382 159588
rect 299474 159576 299480 159588
rect 286376 159548 299480 159576
rect 286376 159536 286382 159548
rect 299474 159536 299480 159548
rect 299532 159536 299538 159588
rect 287514 159468 287520 159520
rect 287572 159508 287578 159520
rect 313274 159508 313280 159520
rect 287572 159480 313280 159508
rect 287572 159468 287578 159480
rect 313274 159468 313280 159480
rect 313332 159468 313338 159520
rect 288986 159400 288992 159452
rect 289044 159440 289050 159452
rect 320174 159440 320180 159452
rect 289044 159412 320180 159440
rect 289044 159400 289050 159412
rect 320174 159400 320180 159412
rect 320232 159400 320238 159452
rect 234614 159332 234620 159384
rect 234672 159372 234678 159384
rect 273806 159372 273812 159384
rect 234672 159344 273812 159372
rect 234672 159332 234678 159344
rect 273806 159332 273812 159344
rect 273864 159332 273870 159384
rect 296530 159332 296536 159384
rect 296588 159372 296594 159384
rect 345934 159372 345940 159384
rect 296588 159344 345940 159372
rect 296588 159332 296594 159344
rect 345934 159332 345940 159344
rect 345992 159332 345998 159384
rect 297266 159264 297272 159316
rect 297324 159304 297330 159316
rect 350994 159304 351000 159316
rect 297324 159276 351000 159304
rect 297324 159264 297330 159276
rect 350994 159264 351000 159276
rect 351052 159264 351058 159316
rect 292298 159196 292304 159248
rect 292356 159236 292362 159248
rect 348234 159236 348240 159248
rect 292356 159208 348240 159236
rect 292356 159196 292362 159208
rect 348234 159196 348240 159208
rect 348292 159196 348298 159248
rect 163498 159128 163504 159180
rect 163556 159168 163562 159180
rect 290458 159168 290464 159180
rect 163556 159140 290464 159168
rect 163556 159128 163562 159140
rect 290458 159128 290464 159140
rect 290516 159128 290522 159180
rect 293770 159128 293776 159180
rect 293828 159168 293834 159180
rect 356054 159168 356060 159180
rect 293828 159140 356060 159168
rect 293828 159128 293834 159140
rect 356054 159128 356060 159140
rect 356112 159128 356118 159180
rect 203426 159060 203432 159112
rect 203484 159100 203490 159112
rect 274082 159100 274088 159112
rect 203484 159072 274088 159100
rect 203484 159060 203490 159072
rect 274082 159060 274088 159072
rect 274140 159060 274146 159112
rect 290734 159060 290740 159112
rect 290792 159100 290798 159112
rect 358446 159100 358452 159112
rect 290792 159072 358452 159100
rect 290792 159060 290798 159072
rect 358446 159060 358452 159072
rect 358504 159060 358510 159112
rect 165982 158992 165988 159044
rect 166040 159032 166046 159044
rect 238110 159032 238116 159044
rect 166040 159004 238116 159032
rect 166040 158992 166046 159004
rect 238110 158992 238116 159004
rect 238168 158992 238174 159044
rect 298554 158992 298560 159044
rect 298612 159032 298618 159044
rect 365898 159032 365904 159044
rect 298612 159004 365904 159032
rect 298612 158992 298618 159004
rect 365898 158992 365904 159004
rect 365956 158992 365962 159044
rect 160922 158924 160928 158976
rect 160980 158964 160986 158976
rect 251910 158964 251916 158976
rect 160980 158936 251916 158964
rect 160980 158924 160986 158936
rect 251910 158924 251916 158936
rect 251968 158924 251974 158976
rect 285214 158924 285220 158976
rect 285272 158964 285278 158976
rect 353570 158964 353576 158976
rect 285272 158936 353576 158964
rect 285272 158924 285278 158936
rect 353570 158924 353576 158936
rect 353628 158924 353634 158976
rect 158530 158856 158536 158908
rect 158588 158896 158594 158908
rect 250438 158896 250444 158908
rect 158588 158868 250444 158896
rect 158588 158856 158594 158868
rect 250438 158856 250444 158868
rect 250496 158856 250502 158908
rect 297174 158856 297180 158908
rect 297232 158896 297238 158908
rect 368198 158896 368204 158908
rect 297232 158868 368204 158896
rect 297232 158856 297238 158868
rect 368198 158856 368204 158868
rect 368256 158856 368262 158908
rect 168282 158788 168288 158840
rect 168340 158828 168346 158840
rect 287698 158828 287704 158840
rect 168340 158800 287704 158828
rect 168340 158788 168346 158800
rect 287698 158788 287704 158800
rect 287756 158788 287762 158840
rect 288158 158788 288164 158840
rect 288216 158828 288222 158840
rect 360838 158828 360844 158840
rect 288216 158800 360844 158828
rect 288216 158788 288222 158800
rect 360838 158788 360844 158800
rect 360896 158788 360902 158840
rect 289630 158720 289636 158772
rect 289688 158760 289694 158772
rect 363414 158760 363420 158772
rect 289688 158732 363420 158760
rect 289688 158720 289694 158732
rect 363414 158720 363420 158732
rect 363472 158720 363478 158772
rect 393498 158720 393504 158772
rect 393556 158760 393562 158772
rect 440510 158760 440516 158772
rect 393556 158732 440516 158760
rect 393556 158720 393562 158732
rect 440510 158720 440516 158732
rect 440568 158720 440574 158772
rect 119706 158652 119712 158704
rect 119764 158692 119770 158704
rect 286134 158692 286140 158704
rect 119764 158664 286140 158692
rect 119764 158652 119770 158664
rect 286134 158652 286140 158664
rect 286192 158652 286198 158704
rect 290918 158652 290924 158704
rect 290976 158692 290982 158704
rect 338390 158692 338396 158704
rect 290976 158664 338396 158692
rect 290976 158652 290982 158664
rect 338390 158652 338396 158664
rect 338448 158652 338454 158704
rect 371050 158652 371056 158704
rect 371108 158692 371114 158704
rect 439590 158692 439596 158704
rect 371108 158664 439596 158692
rect 371108 158652 371114 158664
rect 439590 158652 439596 158664
rect 439648 158652 439654 158704
rect 131298 158584 131304 158636
rect 131356 158624 131362 158636
rect 276014 158624 276020 158636
rect 131356 158596 276020 158624
rect 131356 158584 131362 158596
rect 276014 158584 276020 158596
rect 276072 158584 276078 158636
rect 280890 158584 280896 158636
rect 280948 158624 280954 158636
rect 281166 158624 281172 158636
rect 280948 158596 281172 158624
rect 280948 158584 280954 158596
rect 281166 158584 281172 158596
rect 281224 158584 281230 158636
rect 294966 158584 294972 158636
rect 295024 158624 295030 158636
rect 328270 158624 328276 158636
rect 295024 158596 328276 158624
rect 295024 158584 295030 158596
rect 328270 158584 328276 158596
rect 328328 158584 328334 158636
rect 373442 158584 373448 158636
rect 373500 158624 373506 158636
rect 440418 158624 440424 158636
rect 373500 158596 440424 158624
rect 373500 158584 373506 158596
rect 440418 158584 440424 158596
rect 440476 158584 440482 158636
rect 130194 158516 130200 158568
rect 130252 158556 130258 158568
rect 299014 158556 299020 158568
rect 130252 158528 299020 158556
rect 130252 158516 130258 158528
rect 299014 158516 299020 158528
rect 299072 158556 299078 158568
rect 299290 158556 299296 158568
rect 299072 158528 299296 158556
rect 299072 158516 299078 158528
rect 299290 158516 299296 158528
rect 299348 158516 299354 158568
rect 299566 158516 299572 158568
rect 299624 158556 299630 158568
rect 332226 158556 332232 158568
rect 299624 158528 332232 158556
rect 299624 158516 299630 158528
rect 332226 158516 332232 158528
rect 332284 158516 332290 158568
rect 376018 158516 376024 158568
rect 376076 158556 376082 158568
rect 438026 158556 438032 158568
rect 376076 158528 438032 158556
rect 376076 158516 376082 158528
rect 438026 158516 438032 158528
rect 438084 158516 438090 158568
rect 288250 158488 288256 158500
rect 277366 158460 288256 158488
rect 121178 158380 121184 158432
rect 121236 158420 121242 158432
rect 277366 158420 277394 158460
rect 288250 158448 288256 158460
rect 288308 158488 288314 158500
rect 320542 158488 320548 158500
rect 288308 158460 320548 158488
rect 288308 158448 288314 158460
rect 320542 158448 320548 158460
rect 320600 158448 320606 158500
rect 378594 158448 378600 158500
rect 378652 158488 378658 158500
rect 439406 158488 439412 158500
rect 378652 158460 439412 158488
rect 378652 158448 378658 158460
rect 439406 158448 439412 158460
rect 439464 158448 439470 158500
rect 121236 158392 277394 158420
rect 121236 158380 121242 158392
rect 289446 158380 289452 158432
rect 289504 158420 289510 158432
rect 343542 158420 343548 158432
rect 289504 158392 343548 158420
rect 289504 158380 289510 158392
rect 343542 158380 343548 158392
rect 343600 158380 343606 158432
rect 380986 158380 380992 158432
rect 381044 158420 381050 158432
rect 436830 158420 436836 158432
rect 381044 158392 436836 158420
rect 381044 158380 381050 158392
rect 436830 158380 436836 158392
rect 436888 158380 436894 158432
rect 286594 158312 286600 158364
rect 286652 158352 286658 158364
rect 340966 158352 340972 158364
rect 286652 158324 340972 158352
rect 286652 158312 286658 158324
rect 340966 158312 340972 158324
rect 341024 158312 341030 158364
rect 383562 158312 383568 158364
rect 383620 158352 383626 158364
rect 438118 158352 438124 158364
rect 383620 158324 438124 158352
rect 383620 158312 383626 158324
rect 438118 158312 438124 158324
rect 438176 158312 438182 158364
rect 122098 158244 122104 158296
rect 122156 158284 122162 158296
rect 289630 158284 289636 158296
rect 122156 158256 289636 158284
rect 122156 158244 122162 158256
rect 289630 158244 289636 158256
rect 289688 158244 289694 158296
rect 292206 158244 292212 158296
rect 292264 158284 292270 158296
rect 333606 158284 333612 158296
rect 292264 158256 333612 158284
rect 292264 158244 292270 158256
rect 333606 158244 333612 158256
rect 333664 158244 333670 158296
rect 385954 158244 385960 158296
rect 386012 158284 386018 158296
rect 439498 158284 439504 158296
rect 386012 158256 439504 158284
rect 386012 158244 386018 158256
rect 439498 158244 439504 158256
rect 439556 158244 439562 158296
rect 295886 158176 295892 158228
rect 295944 158216 295950 158228
rect 296622 158216 296628 158228
rect 295944 158188 296628 158216
rect 295944 158176 295950 158188
rect 296622 158176 296628 158188
rect 296680 158216 296686 158228
rect 328638 158216 328644 158228
rect 296680 158188 328644 158216
rect 296680 158176 296686 158188
rect 328638 158176 328644 158188
rect 328696 158176 328702 158228
rect 388530 158176 388536 158228
rect 388588 158216 388594 158228
rect 436922 158216 436928 158228
rect 388588 158188 436928 158216
rect 388588 158176 388594 158188
rect 436922 158176 436928 158188
rect 436980 158176 436986 158228
rect 133506 158108 133512 158160
rect 133564 158148 133570 158160
rect 284570 158148 284576 158160
rect 133564 158120 284576 158148
rect 133564 158108 133570 158120
rect 284570 158108 284576 158120
rect 284628 158108 284634 158160
rect 286134 158108 286140 158160
rect 286192 158148 286198 158160
rect 286778 158148 286784 158160
rect 286192 158120 286784 158148
rect 286192 158108 286198 158120
rect 286778 158108 286784 158120
rect 286836 158148 286842 158160
rect 319438 158148 319444 158160
rect 286836 158120 319444 158148
rect 286836 158108 286842 158120
rect 319438 158108 319444 158120
rect 319496 158108 319502 158160
rect 391474 158108 391480 158160
rect 391532 158148 391538 158160
rect 438302 158148 438308 158160
rect 391532 158120 438308 158148
rect 391532 158108 391538 158120
rect 438302 158108 438308 158120
rect 438360 158108 438366 158160
rect 127618 158040 127624 158092
rect 127676 158080 127682 158092
rect 274634 158080 274640 158092
rect 127676 158052 274640 158080
rect 127676 158040 127682 158052
rect 274634 158040 274640 158052
rect 274692 158040 274698 158092
rect 278314 158040 278320 158092
rect 278372 158080 278378 158092
rect 335998 158080 336004 158092
rect 278372 158052 336004 158080
rect 278372 158040 278378 158052
rect 335998 158040 336004 158052
rect 336056 158040 336062 158092
rect 395890 158040 395896 158092
rect 395948 158080 395954 158092
rect 440602 158080 440608 158092
rect 395948 158052 440608 158080
rect 395948 158040 395954 158052
rect 440602 158040 440608 158052
rect 440660 158040 440666 158092
rect 277210 157972 277216 158024
rect 277268 158012 277274 158024
rect 330478 158012 330484 158024
rect 277268 157984 330484 158012
rect 277268 157972 277274 157984
rect 330478 157972 330484 157984
rect 330536 157972 330542 158024
rect 398466 157972 398472 158024
rect 398524 158012 398530 158024
rect 441706 158012 441712 158024
rect 398524 157984 441712 158012
rect 398524 157972 398530 157984
rect 441706 157972 441712 157984
rect 441764 157972 441770 158024
rect 159818 157904 159824 157956
rect 159876 157944 159882 157956
rect 284662 157944 284668 157956
rect 159876 157916 284668 157944
rect 159876 157904 159882 157916
rect 284662 157904 284668 157916
rect 284720 157904 284726 157956
rect 299290 157904 299296 157956
rect 299348 157944 299354 157956
rect 329926 157944 329932 157956
rect 299348 157916 329932 157944
rect 299348 157904 299354 157916
rect 329926 157904 329932 157916
rect 329984 157904 329990 157956
rect 401410 157904 401416 157956
rect 401468 157944 401474 157956
rect 441798 157944 441804 157956
rect 401468 157916 441804 157944
rect 401468 157904 401474 157916
rect 441798 157904 441804 157916
rect 441856 157904 441862 157956
rect 158162 157836 158168 157888
rect 158220 157876 158226 157888
rect 278682 157876 278688 157888
rect 158220 157848 278688 157876
rect 158220 157836 158226 157848
rect 278682 157836 278688 157848
rect 278740 157836 278746 157888
rect 326430 157876 326436 157888
rect 306346 157848 326436 157876
rect 191098 157768 191104 157820
rect 191156 157808 191162 157820
rect 279602 157808 279608 157820
rect 191156 157780 279608 157808
rect 191156 157768 191162 157780
rect 279602 157768 279608 157780
rect 279660 157768 279666 157820
rect 128722 157700 128728 157752
rect 128780 157740 128786 157752
rect 295886 157740 295892 157752
rect 128780 157712 295892 157740
rect 128780 157700 128786 157712
rect 295886 157700 295892 157712
rect 295944 157700 295950 157752
rect 97626 157632 97632 157684
rect 97684 157672 97690 157684
rect 297542 157672 297548 157684
rect 97684 157644 297548 157672
rect 97684 157632 97690 157644
rect 297542 157632 297548 157644
rect 297600 157632 297606 157684
rect 126514 157564 126520 157616
rect 126572 157604 126578 157616
rect 299198 157604 299204 157616
rect 126572 157576 299204 157604
rect 126572 157564 126578 157576
rect 299198 157564 299204 157576
rect 299256 157604 299262 157616
rect 306346 157604 306374 157848
rect 326430 157836 326436 157848
rect 326488 157836 326494 157888
rect 403802 157836 403808 157888
rect 403860 157876 403866 157888
rect 438210 157876 438216 157888
rect 403860 157848 438216 157876
rect 403860 157836 403866 157848
rect 438210 157836 438216 157848
rect 438268 157836 438274 157888
rect 320082 157768 320088 157820
rect 320140 157808 320146 157820
rect 325142 157808 325148 157820
rect 320140 157780 325148 157808
rect 320140 157768 320146 157780
rect 325142 157768 325148 157780
rect 325200 157768 325206 157820
rect 406746 157768 406752 157820
rect 406804 157808 406810 157820
rect 439682 157808 439688 157820
rect 406804 157780 439688 157808
rect 406804 157768 406810 157780
rect 439682 157768 439688 157780
rect 439740 157768 439746 157820
rect 299256 157576 306374 157604
rect 299256 157564 299262 157576
rect 132402 157496 132408 157548
rect 132460 157536 132466 157548
rect 299106 157536 299112 157548
rect 132460 157508 299112 157536
rect 132460 157496 132466 157508
rect 299106 157496 299112 157508
rect 299164 157496 299170 157548
rect 329190 157428 329196 157480
rect 329248 157468 329254 157480
rect 355226 157468 355232 157480
rect 329248 157440 355232 157468
rect 329248 157428 329254 157440
rect 355226 157428 355232 157440
rect 355284 157428 355290 157480
rect 327350 157360 327356 157412
rect 327408 157400 327414 157412
rect 356974 157400 356980 157412
rect 327408 157372 356980 157400
rect 327408 157360 327414 157372
rect 356974 157360 356980 157372
rect 357032 157360 357038 157412
rect 280982 157292 280988 157344
rect 281040 157332 281046 157344
rect 281166 157332 281172 157344
rect 281040 157304 281172 157332
rect 281040 157292 281046 157304
rect 281166 157292 281172 157304
rect 281224 157332 281230 157344
rect 349798 157332 349804 157344
rect 281224 157304 349804 157332
rect 281224 157292 281230 157304
rect 349798 157292 349804 157304
rect 349856 157292 349862 157344
rect 125318 157224 125324 157276
rect 125376 157264 125382 157276
rect 292390 157264 292396 157276
rect 125376 157236 292396 157264
rect 125376 157224 125382 157236
rect 292390 157224 292396 157236
rect 292448 157264 292454 157276
rect 324222 157264 324228 157276
rect 292448 157236 324228 157264
rect 292448 157224 292454 157236
rect 324222 157224 324228 157236
rect 324280 157224 324286 157276
rect 123202 157156 123208 157208
rect 123260 157196 123266 157208
rect 290826 157196 290832 157208
rect 123260 157168 290832 157196
rect 123260 157156 123266 157168
rect 290826 157156 290832 157168
rect 290884 157196 290890 157208
rect 323118 157196 323124 157208
rect 290884 157168 323124 157196
rect 290884 157156 290890 157168
rect 323118 157156 323124 157168
rect 323176 157156 323182 157208
rect 278130 157088 278136 157140
rect 278188 157128 278194 157140
rect 278406 157128 278412 157140
rect 278188 157100 278412 157128
rect 278188 157088 278194 157100
rect 278406 157088 278412 157100
rect 278464 157128 278470 157140
rect 338758 157128 338764 157140
rect 278464 157100 338764 157128
rect 278464 157088 278470 157100
rect 338758 157088 338764 157100
rect 338816 157088 338822 157140
rect 134886 157020 134892 157072
rect 134944 157060 134950 157072
rect 286870 157060 286876 157072
rect 134944 157032 286876 157060
rect 134944 157020 134950 157032
rect 286870 157020 286876 157032
rect 286928 157060 286934 157072
rect 334526 157060 334532 157072
rect 286928 157032 334532 157060
rect 286928 157020 286934 157032
rect 334526 157020 334532 157032
rect 334584 157020 334590 157072
rect 135898 156952 135904 157004
rect 135956 156992 135962 157004
rect 281442 156992 281448 157004
rect 135956 156964 281448 156992
rect 135956 156952 135962 156964
rect 281442 156952 281448 156964
rect 281500 156992 281506 157004
rect 335630 156992 335636 157004
rect 281500 156964 335636 156992
rect 281500 156952 281506 156964
rect 335630 156952 335636 156964
rect 335688 156952 335694 157004
rect 137002 156884 137008 156936
rect 137060 156924 137066 156936
rect 281350 156924 281356 156936
rect 137060 156896 281356 156924
rect 137060 156884 137066 156896
rect 281350 156884 281356 156896
rect 281408 156924 281414 156936
rect 281408 156896 281948 156924
rect 281408 156884 281414 156896
rect 139210 156816 139216 156868
rect 139268 156856 139274 156868
rect 281920 156856 281948 156896
rect 284478 156884 284484 156936
rect 284536 156924 284542 156936
rect 286318 156924 286324 156936
rect 284536 156896 286324 156924
rect 284536 156884 284542 156896
rect 286318 156884 286324 156896
rect 286376 156884 286382 156936
rect 336826 156924 336832 156936
rect 286428 156896 336832 156924
rect 286428 156856 286456 156896
rect 336826 156884 336832 156896
rect 336884 156884 336890 156936
rect 338114 156856 338120 156868
rect 139268 156828 278268 156856
rect 281920 156828 286456 156856
rect 286520 156828 338120 156856
rect 139268 156816 139274 156828
rect 140682 156748 140688 156800
rect 140740 156788 140746 156800
rect 278130 156788 278136 156800
rect 140740 156760 278136 156788
rect 140740 156748 140746 156760
rect 278130 156748 278136 156760
rect 278188 156748 278194 156800
rect 278240 156788 278268 156828
rect 281258 156788 281264 156800
rect 278240 156760 281264 156788
rect 281258 156748 281264 156760
rect 281316 156788 281322 156800
rect 286520 156788 286548 156828
rect 338114 156816 338120 156828
rect 338172 156816 338178 156868
rect 281316 156760 286548 156788
rect 281316 156748 281322 156760
rect 286594 156748 286600 156800
rect 286652 156788 286658 156800
rect 316034 156788 316040 156800
rect 286652 156760 316040 156788
rect 286652 156748 286658 156760
rect 316034 156748 316040 156760
rect 316092 156748 316098 156800
rect 150250 156680 150256 156732
rect 150308 156720 150314 156732
rect 281166 156720 281172 156732
rect 150308 156692 281172 156720
rect 150308 156680 150314 156692
rect 281166 156680 281172 156692
rect 281224 156680 281230 156732
rect 285950 156680 285956 156732
rect 286008 156720 286014 156732
rect 302234 156720 302240 156732
rect 286008 156692 302240 156720
rect 286008 156680 286014 156692
rect 302234 156680 302240 156692
rect 302292 156680 302298 156732
rect 178954 156612 178960 156664
rect 179012 156652 179018 156664
rect 282270 156652 282276 156664
rect 179012 156624 282276 156652
rect 179012 156612 179018 156624
rect 282270 156612 282276 156624
rect 282328 156612 282334 156664
rect 293494 156612 293500 156664
rect 293552 156652 293558 156664
rect 327074 156652 327080 156664
rect 293552 156624 327080 156652
rect 293552 156612 293558 156624
rect 327074 156612 327080 156624
rect 327132 156612 327138 156664
rect 181714 156544 181720 156596
rect 181772 156584 181778 156596
rect 282178 156584 282184 156596
rect 181772 156556 282184 156584
rect 181772 156544 181778 156556
rect 282178 156544 282184 156556
rect 282236 156544 282242 156596
rect 287422 156544 287428 156596
rect 287480 156584 287486 156596
rect 316034 156584 316040 156596
rect 287480 156556 316040 156584
rect 287480 156544 287486 156556
rect 316034 156544 316040 156556
rect 316092 156544 316098 156596
rect 198458 156476 198464 156528
rect 198516 156516 198522 156528
rect 276934 156516 276940 156528
rect 198516 156488 276940 156516
rect 198516 156476 198522 156488
rect 276934 156476 276940 156488
rect 276992 156476 276998 156528
rect 316678 156516 316684 156528
rect 287026 156488 316684 156516
rect 231854 156408 231860 156460
rect 231912 156448 231918 156460
rect 272242 156448 272248 156460
rect 231912 156420 272248 156448
rect 231912 156408 231918 156420
rect 272242 156408 272248 156420
rect 272300 156408 272306 156460
rect 117314 156340 117320 156392
rect 117372 156380 117378 156392
rect 284110 156380 284116 156392
rect 117372 156352 284116 156380
rect 117372 156340 117378 156352
rect 284110 156340 284116 156352
rect 284168 156380 284174 156392
rect 287026 156380 287054 156488
rect 316678 156476 316684 156488
rect 316736 156476 316742 156528
rect 284168 156352 287054 156380
rect 284168 156340 284174 156352
rect 116854 156272 116860 156324
rect 116912 156312 116918 156324
rect 285490 156312 285496 156324
rect 116912 156284 285496 156312
rect 116912 156272 116918 156284
rect 285490 156272 285496 156284
rect 285548 156312 285554 156324
rect 286594 156312 286600 156324
rect 285548 156284 286600 156312
rect 285548 156272 285554 156284
rect 286594 156272 286600 156284
rect 286652 156272 286658 156324
rect 125410 155864 125416 155916
rect 125468 155904 125474 155916
rect 298922 155904 298928 155916
rect 125468 155876 298928 155904
rect 125468 155864 125474 155876
rect 298922 155864 298928 155876
rect 298980 155904 298986 155916
rect 320082 155904 320088 155916
rect 298980 155876 320088 155904
rect 298980 155864 298986 155876
rect 320082 155864 320088 155876
rect 320140 155864 320146 155916
rect 283558 155796 283564 155848
rect 283616 155836 283622 155848
rect 285950 155836 285956 155848
rect 283616 155808 285956 155836
rect 283616 155796 283622 155808
rect 285950 155796 285956 155808
rect 286008 155796 286014 155848
rect 346394 155836 346400 155848
rect 286060 155808 346400 155836
rect 141786 155728 141792 155780
rect 141844 155768 141850 155780
rect 281074 155768 281080 155780
rect 141844 155740 281080 155768
rect 141844 155728 141850 155740
rect 281074 155728 281080 155740
rect 281132 155768 281138 155780
rect 281442 155768 281448 155780
rect 281132 155740 281448 155768
rect 281132 155728 281138 155740
rect 281442 155728 281448 155740
rect 281500 155728 281506 155780
rect 282362 155728 282368 155780
rect 282420 155768 282426 155780
rect 282822 155768 282828 155780
rect 282420 155740 282828 155768
rect 282420 155728 282426 155740
rect 282822 155728 282828 155740
rect 282880 155768 282886 155780
rect 286060 155768 286088 155808
rect 346394 155796 346400 155808
rect 346452 155796 346458 155848
rect 282880 155740 286088 155768
rect 282880 155728 282886 155740
rect 286134 155728 286140 155780
rect 286192 155768 286198 155780
rect 348694 155768 348700 155780
rect 286192 155740 348700 155768
rect 286192 155728 286198 155740
rect 348694 155728 348700 155740
rect 348752 155728 348758 155780
rect 140590 155660 140596 155712
rect 140648 155700 140654 155712
rect 278498 155700 278504 155712
rect 140648 155672 278504 155700
rect 140648 155660 140654 155672
rect 278498 155660 278504 155672
rect 278556 155700 278562 155712
rect 278682 155700 278688 155712
rect 278556 155672 278688 155700
rect 278556 155660 278562 155672
rect 278682 155660 278688 155672
rect 278740 155660 278746 155712
rect 280062 155660 280068 155712
rect 280120 155700 280126 155712
rect 343910 155700 343916 155712
rect 280120 155672 343916 155700
rect 280120 155660 280126 155672
rect 343910 155660 343916 155672
rect 343968 155660 343974 155712
rect 145282 155592 145288 155644
rect 145340 155632 145346 155644
rect 282730 155632 282736 155644
rect 145340 155604 282736 155632
rect 145340 155592 145346 155604
rect 282730 155592 282736 155604
rect 282788 155632 282794 155644
rect 345106 155632 345112 155644
rect 282788 155604 345112 155632
rect 282788 155592 282794 155604
rect 345106 155592 345112 155604
rect 345164 155592 345170 155644
rect 144270 155524 144276 155576
rect 144328 155564 144334 155576
rect 280062 155564 280068 155576
rect 144328 155536 280068 155564
rect 144328 155524 144334 155536
rect 280062 155524 280068 155536
rect 280120 155524 280126 155576
rect 283374 155524 283380 155576
rect 283432 155564 283438 155576
rect 284202 155564 284208 155576
rect 283432 155536 284208 155564
rect 283432 155524 283438 155536
rect 284202 155524 284208 155536
rect 284260 155564 284266 155576
rect 346854 155564 346860 155576
rect 284260 155536 346860 155564
rect 284260 155524 284266 155536
rect 346854 155524 346860 155536
rect 346912 155524 346918 155576
rect 281442 155456 281448 155508
rect 281500 155496 281506 155508
rect 341150 155496 341156 155508
rect 281500 155468 341156 155496
rect 281500 155456 281506 155468
rect 341150 155456 341156 155468
rect 341208 155456 341214 155508
rect 146386 155388 146392 155440
rect 146444 155428 146450 155440
rect 282362 155428 282368 155440
rect 146444 155400 282368 155428
rect 146444 155388 146450 155400
rect 282362 155388 282368 155400
rect 282420 155388 282426 155440
rect 283466 155388 283472 155440
rect 283524 155428 283530 155440
rect 284018 155428 284024 155440
rect 283524 155400 284024 155428
rect 283524 155388 283530 155400
rect 284018 155388 284024 155400
rect 284076 155428 284082 155440
rect 342806 155428 342812 155440
rect 284076 155400 342812 155428
rect 284076 155388 284082 155400
rect 342806 155388 342812 155400
rect 342864 155388 342870 155440
rect 148778 155320 148784 155372
rect 148836 155360 148842 155372
rect 280890 155360 280896 155372
rect 148836 155332 280896 155360
rect 148836 155320 148842 155332
rect 280890 155320 280896 155332
rect 280948 155360 280954 155372
rect 286134 155360 286140 155372
rect 280948 155332 286140 155360
rect 280948 155320 280954 155332
rect 286134 155320 286140 155332
rect 286192 155320 286198 155372
rect 288894 155320 288900 155372
rect 288952 155360 288958 155372
rect 324314 155360 324320 155372
rect 288952 155332 324320 155360
rect 288952 155320 288958 155332
rect 324314 155320 324320 155332
rect 324372 155320 324378 155372
rect 193950 155252 193956 155304
rect 194008 155292 194014 155304
rect 279510 155292 279516 155304
rect 194008 155264 279516 155292
rect 194008 155252 194014 155264
rect 279510 155252 279516 155264
rect 279568 155252 279574 155304
rect 292942 155252 292948 155304
rect 293000 155292 293006 155304
rect 340874 155292 340880 155304
rect 293000 155264 340880 155292
rect 293000 155252 293006 155264
rect 340874 155252 340880 155264
rect 340932 155252 340938 155304
rect 195882 155184 195888 155236
rect 195940 155224 195946 155236
rect 276842 155224 276848 155236
rect 195940 155196 276848 155224
rect 195940 155184 195946 155196
rect 276842 155184 276848 155196
rect 276900 155184 276906 155236
rect 294322 155184 294328 155236
rect 294380 155224 294386 155236
rect 350534 155224 350540 155236
rect 294380 155196 350540 155224
rect 294380 155184 294386 155196
rect 350534 155184 350540 155196
rect 350592 155184 350598 155236
rect 201034 155116 201040 155168
rect 201092 155156 201098 155168
rect 276750 155156 276756 155168
rect 201092 155128 276756 155156
rect 201092 155116 201098 155128
rect 276750 155116 276756 155128
rect 276808 155116 276814 155168
rect 286042 155116 286048 155168
rect 286100 155156 286106 155168
rect 306374 155156 306380 155168
rect 286100 155128 306380 155156
rect 286100 155116 286106 155128
rect 306374 155116 306380 155128
rect 306432 155116 306438 155168
rect 206278 155048 206284 155100
rect 206336 155088 206342 155100
rect 273898 155088 273904 155100
rect 206336 155060 273904 155088
rect 206336 155048 206342 155060
rect 273898 155048 273904 155060
rect 273956 155048 273962 155100
rect 278682 155048 278688 155100
rect 278740 155088 278746 155100
rect 339494 155088 339500 155100
rect 278740 155060 339500 155088
rect 278740 155048 278746 155060
rect 339494 155048 339500 155060
rect 339552 155048 339558 155100
rect 233234 154980 233240 155032
rect 233292 155020 233298 155032
rect 272150 155020 272156 155032
rect 233292 154992 272156 155020
rect 233292 154980 233298 154992
rect 272150 154980 272156 154992
rect 272208 154980 272214 155032
rect 147766 154912 147772 154964
rect 147824 154952 147830 154964
rect 283374 154952 283380 154964
rect 147824 154924 283380 154952
rect 147824 154912 147830 154924
rect 283374 154912 283380 154924
rect 283432 154912 283438 154964
rect 143074 154844 143080 154896
rect 143132 154884 143138 154896
rect 283466 154884 283472 154896
rect 143132 154856 283472 154884
rect 143132 154844 143138 154856
rect 283466 154844 283472 154856
rect 283524 154844 283530 154896
rect 278682 154504 278688 154556
rect 278740 154544 278746 154556
rect 351086 154544 351092 154556
rect 278740 154516 351092 154544
rect 278740 154504 278746 154516
rect 351086 154504 351092 154516
rect 351144 154504 351150 154556
rect 152642 154436 152648 154488
rect 152700 154476 152706 154488
rect 152700 154448 296714 154476
rect 152700 154436 152706 154448
rect 296686 154408 296714 154448
rect 299290 154436 299296 154488
rect 299348 154476 299354 154488
rect 353294 154476 353300 154488
rect 299348 154448 353300 154476
rect 299348 154436 299354 154448
rect 353294 154436 353300 154448
rect 353352 154436 353358 154488
rect 297910 154408 297916 154420
rect 296686 154380 297916 154408
rect 297910 154368 297916 154380
rect 297968 154408 297974 154420
rect 352190 154408 352196 154420
rect 297968 154380 352196 154408
rect 297968 154368 297974 154380
rect 352190 154368 352196 154380
rect 352248 154368 352254 154420
rect 154482 154300 154488 154352
rect 154540 154340 154546 154352
rect 297818 154340 297824 154352
rect 154540 154312 297824 154340
rect 154540 154300 154546 154312
rect 297818 154300 297824 154312
rect 297876 154340 297882 154352
rect 354398 154340 354404 154352
rect 297876 154312 354404 154340
rect 297876 154300 297882 154312
rect 354398 154300 354404 154312
rect 354456 154300 354462 154352
rect 155770 154232 155776 154284
rect 155828 154272 155834 154284
rect 286686 154272 286692 154284
rect 155828 154244 286692 154272
rect 155828 154232 155834 154244
rect 286686 154232 286692 154244
rect 286744 154272 286750 154284
rect 329190 154272 329196 154284
rect 286744 154244 329196 154272
rect 286744 154232 286750 154244
rect 329190 154232 329196 154244
rect 329248 154232 329254 154284
rect 151354 154164 151360 154216
rect 151412 154204 151418 154216
rect 278682 154204 278688 154216
rect 151412 154176 278688 154204
rect 151412 154164 151418 154176
rect 278682 154164 278688 154176
rect 278740 154164 278746 154216
rect 327350 154204 327356 154216
rect 280172 154176 327356 154204
rect 157058 154096 157064 154148
rect 157116 154136 157122 154148
rect 279970 154136 279976 154148
rect 157116 154108 279976 154136
rect 157116 154096 157122 154108
rect 279970 154096 279976 154108
rect 280028 154136 280034 154148
rect 280172 154136 280200 154176
rect 327350 154164 327356 154176
rect 327408 154164 327414 154216
rect 317690 154136 317696 154148
rect 280028 154108 280200 154136
rect 287026 154108 317696 154136
rect 280028 154096 280034 154108
rect 227714 154028 227720 154080
rect 227772 154068 227778 154080
rect 271138 154068 271144 154080
rect 227772 154040 271144 154068
rect 227772 154028 227778 154040
rect 271138 154028 271144 154040
rect 271196 154028 271202 154080
rect 193214 153960 193220 154012
rect 193272 154000 193278 154012
rect 265434 154000 265440 154012
rect 193272 153972 265440 154000
rect 193272 153960 193278 153972
rect 265434 153960 265440 153972
rect 265492 153960 265498 154012
rect 168374 153892 168380 153944
rect 168432 153932 168438 153944
rect 261386 153932 261392 153944
rect 168432 153904 261392 153932
rect 168432 153892 168438 153904
rect 261386 153892 261392 153904
rect 261444 153892 261450 153944
rect 133874 153824 133880 153876
rect 133932 153864 133938 153876
rect 254394 153864 254400 153876
rect 133932 153836 254400 153864
rect 133932 153824 133938 153836
rect 254394 153824 254400 153836
rect 254452 153824 254458 153876
rect 265618 153824 265624 153876
rect 265676 153864 265682 153876
rect 275002 153864 275008 153876
rect 265676 153836 275008 153864
rect 265676 153824 265682 153836
rect 275002 153824 275008 153836
rect 275060 153824 275066 153876
rect 275094 153824 275100 153876
rect 275152 153864 275158 153876
rect 280430 153864 280436 153876
rect 275152 153836 280436 153864
rect 275152 153824 275158 153836
rect 280430 153824 280436 153836
rect 280488 153824 280494 153876
rect 118234 153756 118240 153808
rect 118292 153796 118298 153808
rect 283926 153796 283932 153808
rect 118292 153768 283932 153796
rect 118292 153756 118298 153768
rect 283926 153756 283932 153768
rect 283984 153796 283990 153808
rect 287026 153796 287054 154108
rect 317690 154096 317696 154108
rect 317748 154096 317754 154148
rect 290090 153824 290096 153876
rect 290148 153864 290154 153876
rect 331214 153864 331220 153876
rect 290148 153836 331220 153864
rect 290148 153824 290154 153836
rect 331214 153824 331220 153836
rect 331272 153824 331278 153876
rect 283984 153768 287054 153796
rect 283984 153756 283990 153768
rect 153930 153688 153936 153740
rect 153988 153728 153994 153740
rect 298186 153728 298192 153740
rect 153988 153700 298192 153728
rect 153988 153688 153994 153700
rect 298186 153688 298192 153700
rect 298244 153728 298250 153740
rect 299290 153728 299296 153740
rect 298244 153700 299296 153728
rect 298244 153688 298250 153700
rect 299290 153688 299296 153700
rect 299348 153688 299354 153740
rect 136082 153144 136088 153196
rect 136140 153184 136146 153196
rect 271322 153184 271328 153196
rect 136140 153156 271328 153184
rect 136140 153144 136146 153156
rect 271322 153144 271328 153156
rect 271380 153144 271386 153196
rect 138934 153076 138940 153128
rect 138992 153116 138998 153128
rect 271414 153116 271420 153128
rect 138992 153088 271420 153116
rect 138992 153076 138998 153088
rect 271414 153076 271420 153088
rect 271472 153076 271478 153128
rect 141418 153008 141424 153060
rect 141476 153048 141482 153060
rect 271230 153048 271236 153060
rect 141476 153020 271236 153048
rect 141476 153008 141482 153020
rect 271230 153008 271236 153020
rect 271288 153008 271294 153060
rect 144362 152940 144368 152992
rect 144420 152980 144426 152992
rect 268562 152980 268568 152992
rect 144420 152952 268568 152980
rect 144420 152940 144426 152952
rect 268562 152940 268568 152952
rect 268620 152940 268626 152992
rect 146018 152872 146024 152924
rect 146076 152912 146082 152924
rect 268470 152912 268476 152924
rect 146076 152884 268476 152912
rect 146076 152872 146082 152884
rect 268470 152872 268476 152884
rect 268528 152872 268534 152924
rect 148410 152804 148416 152856
rect 148468 152844 148474 152856
rect 268378 152844 268384 152856
rect 148468 152816 268384 152844
rect 148468 152804 148474 152816
rect 268378 152804 268384 152816
rect 268436 152804 268442 152856
rect 150986 152736 150992 152788
rect 151044 152776 151050 152788
rect 268654 152776 268660 152788
rect 151044 152748 268660 152776
rect 151044 152736 151050 152748
rect 268654 152736 268660 152748
rect 268712 152736 268718 152788
rect 235994 152668 236000 152720
rect 236052 152708 236058 152720
rect 273714 152708 273720 152720
rect 236052 152680 273720 152708
rect 236052 152668 236058 152680
rect 273714 152668 273720 152680
rect 273772 152668 273778 152720
rect 207014 152600 207020 152652
rect 207072 152640 207078 152652
rect 268194 152640 268200 152652
rect 207072 152612 268200 152640
rect 207072 152600 207078 152612
rect 268194 152600 268200 152612
rect 268252 152600 268258 152652
rect 284386 152600 284392 152652
rect 284444 152640 284450 152652
rect 299566 152640 299572 152652
rect 284444 152612 299572 152640
rect 284444 152600 284450 152612
rect 299566 152600 299572 152612
rect 299624 152600 299630 152652
rect 171134 152532 171140 152584
rect 171192 152572 171198 152584
rect 261294 152572 261300 152584
rect 171192 152544 261300 152572
rect 171192 152532 171198 152544
rect 261294 152532 261300 152544
rect 261352 152532 261358 152584
rect 291654 152532 291660 152584
rect 291712 152572 291718 152584
rect 333974 152572 333980 152584
rect 291712 152544 333980 152572
rect 291712 152532 291718 152544
rect 333974 152532 333980 152544
rect 334032 152532 334038 152584
rect 135254 152464 135260 152516
rect 135312 152504 135318 152516
rect 254302 152504 254308 152516
rect 135312 152476 254308 152504
rect 135312 152464 135318 152476
rect 254302 152464 254308 152476
rect 254360 152464 254366 152516
rect 294598 152464 294604 152516
rect 294656 152504 294662 152516
rect 343634 152504 343640 152516
rect 294656 152476 343640 152504
rect 294656 152464 294662 152476
rect 343634 152464 343640 152476
rect 343692 152464 343698 152516
rect 209774 151172 209780 151224
rect 209832 151212 209838 151224
rect 268102 151212 268108 151224
rect 209832 151184 268108 151212
rect 209832 151172 209838 151184
rect 268102 151172 268108 151184
rect 268160 151172 268166 151224
rect 175274 151104 175280 151156
rect 175332 151144 175338 151156
rect 253198 151144 253204 151156
rect 175332 151116 253204 151144
rect 175332 151104 175338 151116
rect 253198 151104 253204 151116
rect 253256 151104 253262 151156
rect 146294 151036 146300 151088
rect 146352 151076 146358 151088
rect 257154 151076 257160 151088
rect 146352 151048 257160 151076
rect 146352 151036 146358 151048
rect 257154 151036 257160 151048
rect 257212 151036 257218 151088
rect 268194 151036 268200 151088
rect 268252 151076 268258 151088
rect 279142 151076 279148 151088
rect 268252 151048 279148 151076
rect 268252 151036 268258 151048
rect 279142 151036 279148 151048
rect 279200 151036 279206 151088
rect 291562 151036 291568 151088
rect 291620 151076 291626 151088
rect 338114 151076 338120 151088
rect 291620 151048 338120 151076
rect 291620 151036 291626 151048
rect 338114 151036 338120 151048
rect 338172 151036 338178 151088
rect 283282 149880 283288 149932
rect 283340 149920 283346 149932
rect 292942 149920 292948 149932
rect 283340 149892 292948 149920
rect 283340 149880 283346 149892
rect 292942 149880 292948 149892
rect 293000 149880 293006 149932
rect 218054 149812 218060 149864
rect 218112 149852 218118 149864
rect 269574 149852 269580 149864
rect 218112 149824 269580 149852
rect 218112 149812 218118 149824
rect 269574 149812 269580 149824
rect 269632 149812 269638 149864
rect 288802 149812 288808 149864
rect 288860 149852 288866 149864
rect 317414 149852 317420 149864
rect 288860 149824 317420 149852
rect 288860 149812 288866 149824
rect 317414 149812 317420 149824
rect 317472 149812 317478 149864
rect 184934 149744 184940 149796
rect 184992 149784 184998 149796
rect 264054 149784 264060 149796
rect 184992 149756 264060 149784
rect 184992 149744 184998 149756
rect 264054 149744 264060 149756
rect 264112 149744 264118 149796
rect 291470 149744 291476 149796
rect 291528 149784 291534 149796
rect 336734 149784 336740 149796
rect 291528 149756 336740 149784
rect 291528 149744 291534 149756
rect 336734 149744 336740 149756
rect 336792 149744 336798 149796
rect 153194 149676 153200 149728
rect 153252 149716 153258 149728
rect 249150 149716 249156 149728
rect 153252 149688 249156 149716
rect 153252 149676 153258 149688
rect 249150 149676 249156 149688
rect 249208 149676 249214 149728
rect 292850 149676 292856 149728
rect 292908 149716 292914 149728
rect 345014 149716 345020 149728
rect 292908 149688 345020 149716
rect 292908 149676 292914 149688
rect 345014 149676 345020 149688
rect 345072 149676 345078 149728
rect 201494 148452 201500 148504
rect 201552 148492 201558 148504
rect 266722 148492 266728 148504
rect 201552 148464 266728 148492
rect 201552 148452 201558 148464
rect 266722 148452 266728 148464
rect 266780 148452 266786 148504
rect 189074 148384 189080 148436
rect 189132 148424 189138 148436
rect 263962 148424 263968 148436
rect 189132 148396 263968 148424
rect 189132 148384 189138 148396
rect 263962 148384 263968 148396
rect 264020 148384 264026 148436
rect 132494 148316 132500 148368
rect 132552 148356 132558 148368
rect 251818 148356 251824 148368
rect 132552 148328 251824 148356
rect 132552 148316 132558 148328
rect 251818 148316 251824 148328
rect 251876 148316 251882 148368
rect 264330 148316 264336 148368
rect 264388 148356 264394 148368
rect 274910 148356 274916 148368
rect 264388 148328 274916 148356
rect 264388 148316 264394 148328
rect 274910 148316 274916 148328
rect 274968 148316 274974 148368
rect 295794 148316 295800 148368
rect 295852 148356 295858 148368
rect 357434 148356 357440 148368
rect 295852 148328 357440 148356
rect 295852 148316 295858 148328
rect 357434 148316 357440 148328
rect 357492 148316 357498 148368
rect 216674 147024 216680 147076
rect 216732 147064 216738 147076
rect 269482 147064 269488 147076
rect 216732 147036 269488 147064
rect 216732 147024 216738 147036
rect 269482 147024 269488 147036
rect 269540 147024 269546 147076
rect 285858 147024 285864 147076
rect 285916 147064 285922 147076
rect 303614 147064 303620 147076
rect 285916 147036 303620 147064
rect 285916 147024 285922 147036
rect 303614 147024 303620 147036
rect 303672 147024 303678 147076
rect 176654 146956 176660 147008
rect 176712 146996 176718 147008
rect 262398 146996 262404 147008
rect 176712 146968 262404 146996
rect 176712 146956 176718 146968
rect 262398 146956 262404 146968
rect 262456 146956 262462 147008
rect 293310 146956 293316 147008
rect 293368 146996 293374 147008
rect 328454 146996 328460 147008
rect 293368 146968 328460 146996
rect 293368 146956 293374 146968
rect 328454 146956 328460 146968
rect 328512 146956 328518 147008
rect 128354 146888 128360 146940
rect 128412 146928 128418 146940
rect 252738 146928 252744 146940
rect 128412 146900 252744 146928
rect 128412 146888 128418 146900
rect 252738 146888 252744 146900
rect 252796 146888 252802 146940
rect 253198 146888 253204 146940
rect 253256 146928 253262 146940
rect 273622 146928 273628 146940
rect 253256 146900 273628 146928
rect 253256 146888 253262 146900
rect 273622 146888 273628 146900
rect 273680 146888 273686 146940
rect 295702 146888 295708 146940
rect 295760 146928 295766 146940
rect 360194 146928 360200 146940
rect 295760 146900 360200 146928
rect 295760 146888 295766 146900
rect 360194 146888 360200 146900
rect 360252 146888 360258 146940
rect 229094 145664 229100 145716
rect 229152 145704 229158 145716
rect 272058 145704 272064 145716
rect 229152 145676 272064 145704
rect 229152 145664 229158 145676
rect 272058 145664 272064 145676
rect 272116 145664 272122 145716
rect 195974 145596 195980 145648
rect 196032 145636 196038 145648
rect 265342 145636 265348 145648
rect 196032 145608 265348 145636
rect 196032 145596 196038 145608
rect 265342 145596 265348 145608
rect 265400 145596 265406 145648
rect 287330 145596 287336 145648
rect 287388 145636 287394 145648
rect 310514 145636 310520 145648
rect 287388 145608 310520 145636
rect 287388 145596 287394 145608
rect 310514 145596 310520 145608
rect 310572 145596 310578 145648
rect 157334 145528 157340 145580
rect 157392 145568 157398 145580
rect 247678 145568 247684 145580
rect 157392 145540 247684 145568
rect 157392 145528 157398 145540
rect 247678 145528 247684 145540
rect 247736 145528 247742 145580
rect 289998 145528 290004 145580
rect 290056 145568 290062 145580
rect 332594 145568 332600 145580
rect 290056 145540 332600 145568
rect 290056 145528 290062 145540
rect 332594 145528 332600 145540
rect 332652 145528 332658 145580
rect 224954 144304 224960 144356
rect 225012 144344 225018 144356
rect 270862 144344 270868 144356
rect 225012 144316 270868 144344
rect 225012 144304 225018 144316
rect 270862 144304 270868 144316
rect 270920 144304 270926 144356
rect 154574 144236 154580 144288
rect 154632 144276 154638 144288
rect 258350 144276 258356 144288
rect 154632 144248 258356 144276
rect 154632 144236 154638 144248
rect 258350 144236 258356 144248
rect 258408 144236 258414 144288
rect 287238 144236 287244 144288
rect 287296 144276 287302 144288
rect 314654 144276 314660 144288
rect 287296 144248 314660 144276
rect 287296 144236 287302 144248
rect 314654 144236 314660 144248
rect 314712 144236 314718 144288
rect 150434 144168 150440 144220
rect 150492 144208 150498 144220
rect 257062 144208 257068 144220
rect 150492 144180 257068 144208
rect 150492 144168 150498 144180
rect 257062 144168 257068 144180
rect 257120 144168 257126 144220
rect 292758 144168 292764 144220
rect 292816 144208 292822 144220
rect 342254 144208 342260 144220
rect 292816 144180 342260 144208
rect 292816 144168 292822 144180
rect 342254 144168 342260 144180
rect 342312 144168 342318 144220
rect 285030 144032 285036 144084
rect 285088 144072 285094 144084
rect 287330 144072 287336 144084
rect 285088 144044 287336 144072
rect 285088 144032 285094 144044
rect 287330 144032 287336 144044
rect 287388 144032 287394 144084
rect 271138 143760 271144 143812
rect 271196 143800 271202 143812
rect 276198 143800 276204 143812
rect 271196 143772 276204 143800
rect 271196 143760 271202 143772
rect 276198 143760 276204 143772
rect 276256 143760 276262 143812
rect 193306 142876 193312 142928
rect 193364 142916 193370 142928
rect 265250 142916 265256 142928
rect 193364 142888 265256 142916
rect 193364 142876 193370 142888
rect 265250 142876 265256 142888
rect 265308 142876 265314 142928
rect 139394 142808 139400 142860
rect 139452 142848 139458 142860
rect 255774 142848 255780 142860
rect 139452 142820 255780 142848
rect 139452 142808 139458 142820
rect 255774 142808 255780 142820
rect 255832 142808 255838 142860
rect 265342 142808 265348 142860
rect 265400 142848 265406 142860
rect 277670 142848 277676 142860
rect 265400 142820 277676 142848
rect 265400 142808 265406 142820
rect 277670 142808 277676 142820
rect 277728 142808 277734 142860
rect 288710 142808 288716 142860
rect 288768 142848 288774 142860
rect 321554 142848 321560 142860
rect 288768 142820 321560 142848
rect 288768 142808 288774 142820
rect 321554 142808 321560 142820
rect 321612 142808 321618 142860
rect 223574 141516 223580 141568
rect 223632 141556 223638 141568
rect 270770 141556 270776 141568
rect 223632 141528 270776 141556
rect 223632 141516 223638 141528
rect 270770 141516 270776 141528
rect 270828 141516 270834 141568
rect 143534 141448 143540 141500
rect 143592 141488 143598 141500
rect 255682 141488 255688 141500
rect 143592 141460 255688 141488
rect 143592 141448 143598 141460
rect 255682 141448 255688 141460
rect 255740 141448 255746 141500
rect 129734 141380 129740 141432
rect 129792 141420 129798 141432
rect 254210 141420 254216 141432
rect 129792 141392 254216 141420
rect 129792 141380 129798 141392
rect 254210 141380 254216 141392
rect 254268 141380 254274 141432
rect 288618 141380 288624 141432
rect 288676 141420 288682 141432
rect 324406 141420 324412 141432
rect 288676 141392 324412 141420
rect 288676 141380 288682 141392
rect 324406 141380 324412 141392
rect 324464 141380 324470 141432
rect 197354 140088 197360 140140
rect 197412 140128 197418 140140
rect 266630 140128 266636 140140
rect 197412 140100 266636 140128
rect 197412 140088 197418 140100
rect 266630 140088 266636 140100
rect 266688 140088 266694 140140
rect 126974 140020 126980 140072
rect 127032 140060 127038 140072
rect 252646 140060 252652 140072
rect 127032 140032 252652 140060
rect 127032 140020 127038 140032
rect 252646 140020 252652 140032
rect 252704 140020 252710 140072
rect 291378 140020 291384 140072
rect 291436 140060 291442 140072
rect 335354 140060 335360 140072
rect 291436 140032 335360 140060
rect 291436 140020 291442 140032
rect 335354 140020 335360 140032
rect 335412 140020 335418 140072
rect 208394 138796 208400 138848
rect 208452 138836 208458 138848
rect 268010 138836 268016 138848
rect 208452 138808 268016 138836
rect 208452 138796 208458 138808
rect 268010 138796 268016 138808
rect 268068 138796 268074 138848
rect 283190 138796 283196 138848
rect 283248 138836 283254 138848
rect 291378 138836 291384 138848
rect 283248 138808 291384 138836
rect 283248 138796 283254 138808
rect 291378 138796 291384 138808
rect 291436 138796 291442 138848
rect 161474 138728 161480 138780
rect 161532 138768 161538 138780
rect 259822 138768 259828 138780
rect 161532 138740 259828 138768
rect 161532 138728 161538 138740
rect 259822 138728 259828 138740
rect 259880 138728 259886 138780
rect 114554 138660 114560 138712
rect 114612 138700 114618 138712
rect 250162 138700 250168 138712
rect 114612 138672 250168 138700
rect 114612 138660 114618 138672
rect 250162 138660 250168 138672
rect 250220 138660 250226 138712
rect 291286 138660 291292 138712
rect 291344 138700 291350 138712
rect 339494 138700 339500 138712
rect 291344 138672 339500 138700
rect 291344 138660 291350 138672
rect 339494 138660 339500 138672
rect 339552 138660 339558 138712
rect 3142 137912 3148 137964
rect 3200 137952 3206 137964
rect 82078 137952 82084 137964
rect 3200 137924 82084 137952
rect 3200 137912 3206 137924
rect 82078 137912 82084 137924
rect 82136 137912 82142 137964
rect 215294 137368 215300 137420
rect 215352 137408 215358 137420
rect 269390 137408 269396 137420
rect 215352 137380 269396 137408
rect 215352 137368 215358 137380
rect 269390 137368 269396 137380
rect 269448 137368 269454 137420
rect 165614 137300 165620 137352
rect 165672 137340 165678 137352
rect 259730 137340 259736 137352
rect 165672 137312 259736 137340
rect 165672 137300 165678 137312
rect 259730 137300 259736 137312
rect 259788 137300 259794 137352
rect 110414 137232 110420 137284
rect 110472 137272 110478 137284
rect 244918 137272 244924 137284
rect 110472 137244 244924 137272
rect 110472 137232 110478 137244
rect 244918 137232 244924 137244
rect 244976 137232 244982 137284
rect 292666 137232 292672 137284
rect 292724 137272 292730 137284
rect 346394 137272 346400 137284
rect 292724 137244 346400 137272
rect 292724 137232 292730 137244
rect 346394 137232 346400 137244
rect 346452 137232 346458 137284
rect 222194 136008 222200 136060
rect 222252 136048 222258 136060
rect 270678 136048 270684 136060
rect 222252 136020 270684 136048
rect 222252 136008 222258 136020
rect 270678 136008 270684 136020
rect 270736 136008 270742 136060
rect 168466 135940 168472 135992
rect 168524 135980 168530 135992
rect 261110 135980 261116 135992
rect 168524 135952 261116 135980
rect 168524 135940 168530 135952
rect 261110 135940 261116 135952
rect 261168 135940 261174 135992
rect 271230 135940 271236 135992
rect 271288 135980 271294 135992
rect 279050 135980 279056 135992
rect 271288 135952 279056 135980
rect 271288 135940 271294 135952
rect 279050 135940 279056 135952
rect 279108 135940 279114 135992
rect 103514 135872 103520 135924
rect 103572 135912 103578 135924
rect 243722 135912 243728 135924
rect 103572 135884 243728 135912
rect 103572 135872 103578 135884
rect 243722 135872 243728 135884
rect 243780 135872 243786 135924
rect 279510 135192 279516 135244
rect 279568 135232 279574 135244
rect 280338 135232 280344 135244
rect 279568 135204 280344 135232
rect 279568 135192 279574 135204
rect 280338 135192 280344 135204
rect 280396 135192 280402 135244
rect 172514 134580 172520 134632
rect 172572 134620 172578 134632
rect 261018 134620 261024 134632
rect 172572 134592 261024 134620
rect 172572 134580 172578 134592
rect 261018 134580 261024 134592
rect 261076 134580 261082 134632
rect 147674 134512 147680 134564
rect 147732 134552 147738 134564
rect 256970 134552 256976 134564
rect 147732 134524 256976 134552
rect 147732 134512 147738 134524
rect 256970 134512 256976 134524
rect 257028 134512 257034 134564
rect 261478 134512 261484 134564
rect 261536 134552 261542 134564
rect 276106 134552 276112 134564
rect 261536 134524 276112 134552
rect 261536 134512 261542 134524
rect 276106 134512 276112 134524
rect 276164 134512 276170 134564
rect 179414 133220 179420 133272
rect 179472 133260 179478 133272
rect 262306 133260 262312 133272
rect 179472 133232 262312 133260
rect 179472 133220 179478 133232
rect 262306 133220 262312 133232
rect 262364 133220 262370 133272
rect 158714 133152 158720 133204
rect 158772 133192 158778 133204
rect 258258 133192 258264 133204
rect 158772 133164 258264 133192
rect 158772 133152 158778 133164
rect 258258 133152 258264 133164
rect 258316 133152 258322 133204
rect 191834 131792 191840 131844
rect 191892 131832 191898 131844
rect 265158 131832 265164 131844
rect 191892 131804 265164 131832
rect 191892 131792 191898 131804
rect 265158 131792 265164 131804
rect 265216 131792 265222 131844
rect 183554 131724 183560 131776
rect 183612 131764 183618 131776
rect 263870 131764 263876 131776
rect 183612 131736 263876 131764
rect 183612 131724 183618 131736
rect 263870 131724 263876 131736
rect 263928 131724 263934 131776
rect 205634 130500 205640 130552
rect 205692 130540 205698 130552
rect 267918 130540 267924 130552
rect 205692 130512 267924 130540
rect 205692 130500 205698 130512
rect 267918 130500 267924 130512
rect 267976 130500 267982 130552
rect 186314 130432 186320 130484
rect 186372 130472 186378 130484
rect 263778 130472 263784 130484
rect 186372 130444 263784 130472
rect 186372 130432 186378 130444
rect 263778 130432 263784 130444
rect 263836 130432 263842 130484
rect 118694 130364 118700 130416
rect 118752 130404 118758 130416
rect 251450 130404 251456 130416
rect 118752 130376 251456 130404
rect 118752 130364 118758 130376
rect 251450 130364 251456 130376
rect 251508 130364 251514 130416
rect 288526 130364 288532 130416
rect 288584 130404 288590 130416
rect 318794 130404 318800 130416
rect 288584 130376 318800 130404
rect 288584 130364 288590 130376
rect 318794 130364 318800 130376
rect 318852 130364 318858 130416
rect 230474 129140 230480 129192
rect 230532 129180 230538 129192
rect 271966 129180 271972 129192
rect 230532 129152 271972 129180
rect 230532 129140 230538 129152
rect 271966 129140 271972 129152
rect 272024 129140 272030 129192
rect 190454 129072 190460 129124
rect 190512 129112 190518 129124
rect 265066 129112 265072 129124
rect 190512 129084 265072 129112
rect 190512 129072 190518 129084
rect 265066 129072 265072 129084
rect 265124 129072 265130 129124
rect 107654 129004 107660 129056
rect 107712 129044 107718 129056
rect 242342 129044 242348 129056
rect 107712 129016 242348 129044
rect 107712 129004 107718 129016
rect 242342 129004 242348 129016
rect 242400 129004 242406 129056
rect 289906 129004 289912 129056
rect 289964 129044 289970 129056
rect 325694 129044 325700 129056
rect 289964 129016 325700 129044
rect 289964 129004 289970 129016
rect 325694 129004 325700 129016
rect 325752 129004 325758 129056
rect 204254 127644 204260 127696
rect 204312 127684 204318 127696
rect 266538 127684 266544 127696
rect 204312 127656 266544 127684
rect 204312 127644 204318 127656
rect 266538 127644 266544 127656
rect 266596 127644 266602 127696
rect 100754 127576 100760 127628
rect 100812 127616 100818 127628
rect 246390 127616 246396 127628
rect 100812 127588 246396 127616
rect 100812 127576 100818 127588
rect 246390 127576 246396 127588
rect 246448 127576 246454 127628
rect 291194 127576 291200 127628
rect 291252 127616 291258 127628
rect 332686 127616 332692 127628
rect 291252 127588 332692 127616
rect 291252 127576 291258 127588
rect 332686 127576 332692 127588
rect 332744 127576 332750 127628
rect 211154 126284 211160 126336
rect 211212 126324 211218 126336
rect 267826 126324 267832 126336
rect 211212 126296 267832 126324
rect 211212 126284 211218 126296
rect 267826 126284 267832 126296
rect 267884 126284 267890 126336
rect 155954 126216 155960 126268
rect 156012 126256 156018 126268
rect 258166 126256 258172 126268
rect 156012 126228 258172 126256
rect 156012 126216 156018 126228
rect 258166 126216 258172 126228
rect 258224 126216 258230 126268
rect 267918 126216 267924 126268
rect 267976 126256 267982 126268
rect 278958 126256 278964 126268
rect 267976 126228 278964 126256
rect 267976 126216 267982 126228
rect 278958 126216 278964 126228
rect 279016 126216 279022 126268
rect 292574 126216 292580 126268
rect 292632 126256 292638 126268
rect 340966 126256 340972 126268
rect 292632 126228 340972 126256
rect 292632 126216 292638 126228
rect 340966 126216 340972 126228
rect 341024 126216 341030 126268
rect 218146 124924 218152 124976
rect 218204 124964 218210 124976
rect 269298 124964 269304 124976
rect 218204 124936 269304 124964
rect 218204 124924 218210 124936
rect 269298 124924 269304 124936
rect 269356 124924 269362 124976
rect 138014 124856 138020 124908
rect 138072 124896 138078 124908
rect 255590 124896 255596 124908
rect 138072 124868 255596 124896
rect 138072 124856 138078 124868
rect 255590 124856 255596 124868
rect 255648 124856 255654 124908
rect 296070 124856 296076 124908
rect 296128 124896 296134 124908
rect 354674 124896 354680 124908
rect 296128 124868 354680 124896
rect 296128 124856 296134 124868
rect 354674 124856 354680 124868
rect 354732 124856 354738 124908
rect 226334 123496 226340 123548
rect 226392 123536 226398 123548
rect 270586 123536 270592 123548
rect 226392 123508 270592 123536
rect 226392 123496 226398 123508
rect 270586 123496 270592 123508
rect 270644 123496 270650 123548
rect 173894 123428 173900 123480
rect 173952 123468 173958 123480
rect 260926 123468 260932 123480
rect 173952 123440 260932 123468
rect 173952 123428 173958 123440
rect 260926 123428 260932 123440
rect 260984 123428 260990 123480
rect 234706 122136 234712 122188
rect 234764 122176 234770 122188
rect 272334 122176 272340 122188
rect 234764 122148 272340 122176
rect 234764 122136 234770 122148
rect 272334 122136 272340 122148
rect 272392 122136 272398 122188
rect 136634 122068 136640 122120
rect 136692 122108 136698 122120
rect 254118 122108 254124 122120
rect 136692 122080 254124 122108
rect 136692 122068 136698 122080
rect 254118 122068 254124 122080
rect 254176 122068 254182 122120
rect 140774 120708 140780 120760
rect 140832 120748 140838 120760
rect 255498 120748 255504 120760
rect 140832 120720 255504 120748
rect 140832 120708 140838 120720
rect 255498 120708 255504 120720
rect 255556 120708 255562 120760
rect 255958 120708 255964 120760
rect 256016 120748 256022 120760
rect 274818 120748 274824 120760
rect 256016 120720 274824 120748
rect 256016 120708 256022 120720
rect 274818 120708 274824 120720
rect 274876 120708 274882 120760
rect 143626 119348 143632 119400
rect 143684 119388 143690 119400
rect 255406 119388 255412 119400
rect 143684 119360 255412 119388
rect 143684 119348 143690 119360
rect 255406 119348 255412 119360
rect 255464 119348 255470 119400
rect 151814 117920 151820 117972
rect 151872 117960 151878 117972
rect 256878 117960 256884 117972
rect 151872 117932 256884 117960
rect 151872 117920 151878 117932
rect 256878 117920 256884 117932
rect 256936 117920 256942 117972
rect 127066 116560 127072 116612
rect 127124 116600 127130 116612
rect 253014 116600 253020 116612
rect 127124 116572 253020 116600
rect 127124 116560 127130 116572
rect 253014 116560 253020 116572
rect 253072 116560 253078 116612
rect 162854 115200 162860 115252
rect 162912 115240 162918 115252
rect 259638 115240 259644 115252
rect 162912 115212 259644 115240
rect 162912 115200 162918 115212
rect 259638 115200 259644 115212
rect 259696 115200 259702 115252
rect 169754 113772 169760 113824
rect 169812 113812 169818 113824
rect 260834 113812 260840 113824
rect 169812 113784 260840 113812
rect 169812 113772 169818 113784
rect 260834 113772 260840 113784
rect 260892 113772 260898 113824
rect 442258 113092 442264 113144
rect 442316 113132 442322 113144
rect 579798 113132 579804 113144
rect 442316 113104 579804 113132
rect 442316 113092 442322 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 166994 112412 167000 112464
rect 167052 112452 167058 112464
rect 259546 112452 259552 112464
rect 167052 112424 259552 112452
rect 167052 112412 167058 112424
rect 259546 112412 259552 112424
rect 259604 112412 259610 112464
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 84838 111772 84844 111784
rect 3200 111744 84844 111772
rect 3200 111732 3206 111744
rect 84838 111732 84844 111744
rect 84896 111732 84902 111784
rect 180794 111052 180800 111104
rect 180852 111092 180858 111104
rect 262582 111092 262588 111104
rect 180852 111064 262588 111092
rect 180852 111052 180858 111064
rect 262582 111052 262588 111064
rect 262640 111052 262646 111104
rect 185026 109692 185032 109744
rect 185084 109732 185090 109744
rect 263686 109732 263692 109744
rect 185084 109704 263692 109732
rect 185084 109692 185090 109704
rect 263686 109692 263692 109704
rect 263744 109692 263750 109744
rect 187694 108264 187700 108316
rect 187752 108304 187758 108316
rect 263594 108304 263600 108316
rect 187752 108276 263600 108304
rect 187752 108264 187758 108276
rect 263594 108264 263600 108276
rect 263652 108264 263658 108316
rect 264422 108264 264428 108316
rect 264480 108304 264486 108316
rect 277578 108304 277584 108316
rect 264480 108276 277584 108304
rect 264480 108264 264486 108276
rect 277578 108264 277584 108276
rect 277636 108264 277642 108316
rect 131114 106904 131120 106956
rect 131172 106944 131178 106956
rect 254026 106944 254032 106956
rect 131172 106916 254032 106944
rect 131172 106904 131178 106916
rect 254026 106904 254032 106916
rect 254084 106904 254090 106956
rect 266538 106904 266544 106956
rect 266596 106944 266602 106956
rect 276658 106944 276664 106956
rect 266596 106916 276664 106944
rect 266596 106904 266602 106916
rect 276658 106904 276664 106916
rect 276716 106904 276722 106956
rect 198734 105544 198740 105596
rect 198792 105584 198798 105596
rect 266446 105584 266452 105596
rect 198792 105556 266452 105584
rect 198792 105544 198798 105556
rect 266446 105544 266452 105556
rect 266504 105544 266510 105596
rect 209866 104184 209872 104236
rect 209924 104224 209930 104236
rect 267734 104224 267740 104236
rect 209924 104196 267740 104224
rect 209924 104184 209930 104196
rect 267734 104184 267740 104196
rect 267792 104184 267798 104236
rect 106274 104116 106280 104168
rect 106332 104156 106338 104168
rect 248598 104156 248604 104168
rect 106332 104128 248604 104156
rect 106332 104116 106338 104128
rect 248598 104116 248604 104128
rect 248656 104116 248662 104168
rect 219434 102824 219440 102876
rect 219492 102864 219498 102876
rect 269206 102864 269212 102876
rect 219492 102836 269212 102864
rect 219492 102824 219498 102836
rect 269206 102824 269212 102836
rect 269264 102824 269270 102876
rect 111794 102756 111800 102808
rect 111852 102796 111858 102808
rect 250070 102796 250076 102808
rect 111852 102768 250076 102796
rect 111852 102756 111858 102768
rect 250070 102756 250076 102768
rect 250128 102756 250134 102808
rect 142154 101396 142160 101448
rect 142212 101436 142218 101448
rect 255314 101436 255320 101448
rect 142212 101408 255320 101436
rect 142212 101396 142218 101408
rect 255314 101396 255320 101408
rect 255372 101396 255378 101448
rect 149054 99968 149060 100020
rect 149112 100008 149118 100020
rect 256786 100008 256792 100020
rect 149112 99980 256792 100008
rect 149112 99968 149118 99980
rect 256786 99968 256792 99980
rect 256844 99968 256850 100020
rect 160186 98608 160192 98660
rect 160244 98648 160250 98660
rect 258442 98648 258448 98660
rect 160244 98620 258448 98648
rect 160244 98608 160250 98620
rect 258442 98608 258448 98620
rect 258500 98608 258506 98660
rect 121454 97248 121460 97300
rect 121512 97288 121518 97300
rect 251358 97288 251364 97300
rect 121512 97260 251364 97288
rect 121512 97248 121518 97260
rect 251358 97248 251364 97260
rect 251416 97248 251422 97300
rect 109034 94460 109040 94512
rect 109092 94500 109098 94512
rect 249978 94500 249984 94512
rect 109092 94472 249984 94500
rect 109092 94460 109098 94472
rect 249978 94460 249984 94472
rect 250036 94460 250042 94512
rect 115934 93100 115940 93152
rect 115992 93140 115998 93152
rect 249058 93140 249064 93152
rect 115992 93112 249064 93140
rect 115992 93100 115998 93112
rect 249058 93100 249064 93112
rect 249116 93100 249122 93152
rect 99374 91740 99380 91792
rect 99432 91780 99438 91792
rect 247310 91780 247316 91792
rect 99432 91752 247316 91780
rect 99432 91740 99438 91752
rect 247310 91740 247316 91752
rect 247368 91740 247374 91792
rect 113818 90312 113824 90364
rect 113876 90352 113882 90364
rect 249886 90352 249892 90364
rect 113876 90324 249892 90352
rect 113876 90312 113882 90324
rect 249886 90312 249892 90324
rect 249944 90312 249950 90364
rect 49694 88952 49700 89004
rect 49752 88992 49758 89004
rect 239306 88992 239312 89004
rect 49752 88964 239312 88992
rect 49752 88952 49758 88964
rect 239306 88952 239312 88964
rect 239364 88952 239370 89004
rect 120074 86232 120080 86284
rect 120132 86272 120138 86284
rect 242250 86272 242256 86284
rect 120132 86244 242256 86272
rect 120132 86232 120138 86244
rect 242250 86232 242256 86244
rect 242308 86232 242314 86284
rect 3418 85484 3424 85536
rect 3476 85524 3482 85536
rect 80698 85524 80704 85536
rect 3476 85496 80704 85524
rect 3476 85484 3482 85496
rect 80698 85484 80704 85496
rect 80756 85484 80762 85536
rect 104894 64132 104900 64184
rect 104952 64172 104958 64184
rect 248506 64172 248512 64184
rect 104952 64144 248512 64172
rect 104952 64132 104958 64144
rect 248506 64132 248512 64144
rect 248564 64132 248570 64184
rect 47578 33736 47584 33788
rect 47636 33776 47642 33788
rect 237466 33776 237472 33788
rect 47636 33748 237472 33776
rect 47636 33736 47642 33748
rect 237466 33736 237472 33748
rect 237524 33736 237530 33788
rect 526438 33056 526444 33108
rect 526496 33096 526502 33108
rect 580166 33096 580172 33108
rect 526496 33068 580172 33096
rect 526496 33056 526502 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 117958 25508 117964 25560
rect 118016 25548 118022 25560
rect 250254 25548 250260 25560
rect 118016 25520 250260 25548
rect 118016 25508 118022 25520
rect 250254 25508 250260 25520
rect 250312 25508 250318 25560
rect 151906 24080 151912 24132
rect 151964 24120 151970 24132
rect 257338 24120 257344 24132
rect 151964 24092 257344 24120
rect 151964 24080 151970 24092
rect 257338 24080 257344 24092
rect 257396 24080 257402 24132
rect 295978 24080 295984 24132
rect 296036 24120 296042 24132
rect 347774 24120 347780 24132
rect 296036 24092 347780 24120
rect 296036 24080 296042 24092
rect 347774 24080 347780 24092
rect 347832 24080 347838 24132
rect 144914 22720 144920 22772
rect 144972 22760 144978 22772
rect 256694 22760 256700 22772
rect 144972 22732 256700 22760
rect 144972 22720 144978 22732
rect 256694 22720 256700 22732
rect 256752 22720 256758 22772
rect 212534 21360 212540 21412
rect 212592 21400 212598 21412
rect 269114 21400 269120 21412
rect 212592 21372 269120 21400
rect 212592 21360 212598 21372
rect 269114 21360 269120 21372
rect 269172 21360 269178 21412
rect 201586 19932 201592 19984
rect 201644 19972 201650 19984
rect 266906 19972 266912 19984
rect 201644 19944 266912 19972
rect 201644 19932 201650 19944
rect 266906 19932 266912 19944
rect 266964 19932 266970 19984
rect 194594 18572 194600 18624
rect 194652 18612 194658 18624
rect 264974 18612 264980 18624
rect 194652 18584 264980 18612
rect 194652 18572 194658 18584
rect 264974 18572 264980 18584
rect 265032 18572 265038 18624
rect 295610 18572 295616 18624
rect 295668 18612 295674 18624
rect 361574 18612 361580 18624
rect 295668 18584 361580 18612
rect 295668 18572 295674 18584
rect 361574 18572 361580 18584
rect 361632 18572 361638 18624
rect 135346 17280 135352 17332
rect 135404 17320 135410 17332
rect 254486 17320 254492 17332
rect 135404 17292 254492 17320
rect 135404 17280 135410 17292
rect 254486 17280 254492 17292
rect 254544 17280 254550 17332
rect 254026 17212 254032 17264
rect 254084 17252 254090 17264
rect 275278 17252 275284 17264
rect 254084 17224 275284 17252
rect 254084 17212 254090 17224
rect 275278 17212 275284 17224
rect 275336 17212 275342 17264
rect 288434 17212 288440 17264
rect 288492 17252 288498 17264
rect 322934 17252 322940 17264
rect 288492 17224 322940 17252
rect 288492 17212 288498 17224
rect 322934 17212 322940 17224
rect 322992 17212 322998 17264
rect 242894 15852 242900 15904
rect 242952 15892 242958 15904
rect 273530 15892 273536 15904
rect 242952 15864 273536 15892
rect 242952 15852 242958 15864
rect 273530 15852 273536 15864
rect 273588 15852 273594 15904
rect 289814 15852 289820 15904
rect 289872 15892 289878 15904
rect 330386 15892 330392 15904
rect 289872 15864 330392 15892
rect 289872 15852 289878 15864
rect 330386 15852 330392 15864
rect 330444 15852 330450 15904
rect 42794 14424 42800 14476
rect 42852 14464 42858 14476
rect 237834 14464 237840 14476
rect 42852 14436 237840 14464
rect 42852 14424 42858 14436
rect 237834 14424 237840 14436
rect 237892 14424 237898 14476
rect 291838 14424 291844 14476
rect 291896 14464 291902 14476
rect 305546 14464 305552 14476
rect 291896 14436 305552 14464
rect 291896 14424 291902 14436
rect 305546 14424 305552 14436
rect 305604 14424 305610 14476
rect 273898 13948 273904 14000
rect 273956 13988 273962 14000
rect 278866 13988 278872 14000
rect 273956 13960 278872 13988
rect 273956 13948 273962 13960
rect 278866 13948 278872 13960
rect 278924 13948 278930 14000
rect 255866 13132 255872 13184
rect 255924 13172 255930 13184
rect 264238 13172 264244 13184
rect 255924 13144 264244 13172
rect 255924 13132 255930 13144
rect 264238 13132 264244 13144
rect 264296 13132 264302 13184
rect 81618 13064 81624 13116
rect 81676 13104 81682 13116
rect 242158 13104 242164 13116
rect 81676 13076 242164 13104
rect 81676 13064 81682 13076
rect 242158 13064 242164 13076
rect 242216 13064 242222 13116
rect 260006 13064 260012 13116
rect 260064 13104 260070 13116
rect 277486 13104 277492 13116
rect 260064 13076 277492 13104
rect 260064 13064 260070 13076
rect 277486 13064 277492 13076
rect 277544 13064 277550 13116
rect 287146 13064 287152 13116
rect 287204 13104 287210 13116
rect 312170 13104 312176 13116
rect 287204 13076 312176 13104
rect 287204 13064 287210 13076
rect 312170 13064 312176 13076
rect 312228 13064 312234 13116
rect 278130 12452 278136 12504
rect 278188 12492 278194 12504
rect 280246 12492 280252 12504
rect 278188 12464 280252 12492
rect 278188 12452 278194 12464
rect 280246 12452 280252 12464
rect 280304 12452 280310 12504
rect 280706 12452 280712 12504
rect 280764 12492 280770 12504
rect 281902 12492 281908 12504
rect 280764 12464 281908 12492
rect 280764 12452 280770 12464
rect 281902 12452 281908 12464
rect 281960 12452 281966 12504
rect 439130 11880 439136 11892
rect 439056 11852 439136 11880
rect 160094 11772 160100 11824
rect 160152 11812 160158 11824
rect 161290 11812 161296 11824
rect 160152 11784 161296 11812
rect 160152 11772 160158 11784
rect 161290 11772 161296 11784
rect 161348 11772 161354 11824
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 234614 11772 234620 11824
rect 234672 11812 234678 11824
rect 235810 11812 235816 11824
rect 234672 11784 235816 11812
rect 234672 11772 234678 11784
rect 235810 11772 235816 11784
rect 235868 11772 235874 11824
rect 102134 11704 102140 11756
rect 102192 11744 102198 11756
rect 246298 11744 246304 11756
rect 102192 11716 246304 11744
rect 102192 11704 102198 11716
rect 246298 11704 246304 11716
rect 246356 11704 246362 11756
rect 287054 11704 287060 11756
rect 287112 11744 287118 11756
rect 316218 11744 316224 11756
rect 287112 11716 316224 11744
rect 287112 11704 287118 11716
rect 316218 11704 316224 11716
rect 316276 11704 316282 11756
rect 439056 11688 439084 11852
rect 439130 11840 439136 11852
rect 439188 11840 439194 11892
rect 439038 11636 439044 11688
rect 439096 11636 439102 11688
rect 270770 10480 270776 10532
rect 270828 10520 270834 10532
rect 278038 10520 278044 10532
rect 270828 10492 278044 10520
rect 270828 10480 270834 10492
rect 278038 10480 278044 10492
rect 278096 10480 278102 10532
rect 237650 10344 237656 10396
rect 237708 10384 237714 10396
rect 273438 10384 273444 10396
rect 237708 10356 273444 10384
rect 237708 10344 237714 10356
rect 273438 10344 273444 10356
rect 273496 10344 273502 10396
rect 53006 10276 53012 10328
rect 53064 10316 53070 10328
rect 239214 10316 239220 10328
rect 53064 10288 239220 10316
rect 53064 10276 53070 10288
rect 239214 10276 239220 10288
rect 239272 10276 239278 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 283098 9120 283104 9172
rect 283156 9160 283162 9172
rect 292574 9160 292580 9172
rect 283156 9132 292580 9160
rect 283156 9120 283162 9132
rect 292574 9120 292580 9132
rect 292632 9120 292638 9172
rect 289354 9052 289360 9104
rect 289412 9092 289418 9104
rect 410794 9092 410800 9104
rect 289412 9064 410800 9092
rect 289412 9052 289418 9064
rect 410794 9052 410800 9064
rect 410852 9052 410858 9104
rect 241698 8984 241704 9036
rect 241756 9024 241762 9036
rect 273346 9024 273352 9036
rect 241756 8996 273352 9024
rect 241756 8984 241762 8996
rect 273346 8984 273352 8996
rect 273404 8984 273410 9036
rect 285398 8984 285404 9036
rect 285456 9024 285462 9036
rect 411898 9024 411904 9036
rect 285456 8996 411904 9024
rect 285456 8984 285462 8996
rect 411898 8984 411904 8996
rect 411956 8984 411962 9036
rect 123478 8916 123484 8968
rect 123536 8956 123542 8968
rect 243538 8956 243544 8968
rect 123536 8928 243544 8956
rect 123536 8916 123542 8928
rect 243538 8916 243544 8928
rect 243596 8916 243602 8968
rect 248782 8916 248788 8968
rect 248840 8956 248846 8968
rect 262858 8956 262864 8968
rect 248840 8928 262864 8956
rect 248840 8916 248846 8928
rect 262858 8916 262864 8928
rect 262916 8916 262922 8968
rect 288066 8916 288072 8968
rect 288124 8956 288130 8968
rect 414290 8956 414296 8968
rect 288124 8928 414296 8956
rect 288124 8916 288130 8928
rect 414290 8916 414296 8928
rect 414348 8916 414354 8968
rect 281810 8236 281816 8288
rect 281868 8276 281874 8288
rect 283098 8276 283104 8288
rect 281868 8248 283104 8276
rect 281868 8236 281874 8248
rect 283098 8236 283104 8248
rect 283156 8236 283162 8288
rect 240502 7624 240508 7676
rect 240560 7664 240566 7676
rect 273254 7664 273260 7676
rect 240560 7636 273260 7664
rect 240560 7624 240566 7636
rect 273254 7624 273260 7636
rect 273312 7624 273318 7676
rect 227530 7556 227536 7608
rect 227588 7596 227594 7608
rect 270494 7596 270500 7608
rect 227588 7568 270500 7596
rect 227588 7556 227594 7568
rect 270494 7556 270500 7568
rect 270552 7556 270558 7608
rect 276014 7556 276020 7608
rect 276072 7596 276078 7608
rect 280522 7596 280528 7608
rect 276072 7568 280528 7596
rect 276072 7556 276078 7568
rect 280522 7556 280528 7568
rect 280580 7556 280586 7608
rect 299566 7556 299572 7608
rect 299624 7596 299630 7608
rect 300762 7596 300768 7608
rect 299624 7568 300768 7596
rect 299624 7556 299630 7568
rect 300762 7556 300768 7568
rect 300820 7556 300826 7608
rect 283006 6944 283012 6996
rect 283064 6984 283070 6996
rect 288986 6984 288992 6996
rect 283064 6956 288992 6984
rect 283064 6944 283070 6956
rect 288986 6944 288992 6956
rect 289044 6944 289050 6996
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 40678 6848 40684 6860
rect 3476 6820 40684 6848
rect 3476 6808 3482 6820
rect 40678 6808 40684 6820
rect 40736 6808 40742 6860
rect 295518 6740 295524 6792
rect 295576 6780 295582 6792
rect 358722 6780 358728 6792
rect 295576 6752 358728 6780
rect 295576 6740 295582 6752
rect 358722 6740 358728 6752
rect 358780 6740 358786 6792
rect 291102 6672 291108 6724
rect 291160 6712 291166 6724
rect 378870 6712 378876 6724
rect 291160 6684 378876 6712
rect 291160 6672 291166 6684
rect 378870 6672 378876 6684
rect 378928 6672 378934 6724
rect 291010 6604 291016 6656
rect 291068 6644 291074 6656
rect 385954 6644 385960 6656
rect 291068 6616 385960 6644
rect 291068 6604 291074 6616
rect 385954 6604 385960 6616
rect 386012 6604 386018 6656
rect 287882 6536 287888 6588
rect 287940 6576 287946 6588
rect 400122 6576 400128 6588
rect 287940 6548 400128 6576
rect 287940 6536 287946 6548
rect 400122 6536 400128 6548
rect 400180 6536 400186 6588
rect 289722 6468 289728 6520
rect 289780 6508 289786 6520
rect 403618 6508 403624 6520
rect 289780 6480 403624 6508
rect 289780 6468 289786 6480
rect 403618 6468 403624 6480
rect 403676 6468 403682 6520
rect 284938 6400 284944 6452
rect 284996 6440 285002 6452
rect 294874 6440 294880 6452
rect 284996 6412 294880 6440
rect 284996 6400 285002 6412
rect 294874 6400 294880 6412
rect 294932 6400 294938 6452
rect 294966 6400 294972 6452
rect 295024 6440 295030 6452
rect 413094 6440 413100 6452
rect 295024 6412 413100 6440
rect 295024 6400 295030 6412
rect 413094 6400 413100 6412
rect 413152 6400 413158 6452
rect 287974 6332 287980 6384
rect 288032 6372 288038 6384
rect 407206 6372 407212 6384
rect 288032 6344 407212 6372
rect 288032 6332 288038 6344
rect 407206 6332 407212 6344
rect 407264 6332 407270 6384
rect 290642 6264 290648 6316
rect 290700 6304 290706 6316
rect 416682 6304 416688 6316
rect 290700 6276 416688 6304
rect 290700 6264 290706 6276
rect 416682 6264 416688 6276
rect 416740 6264 416746 6316
rect 247586 6196 247592 6248
rect 247644 6236 247650 6248
rect 274726 6236 274732 6248
rect 247644 6208 274732 6236
rect 247644 6196 247650 6208
rect 274726 6196 274732 6208
rect 274784 6196 274790 6248
rect 292482 6196 292488 6248
rect 292540 6236 292546 6248
rect 420178 6236 420184 6248
rect 292540 6208 420184 6236
rect 292540 6196 292546 6208
rect 420178 6196 420184 6208
rect 420236 6196 420242 6248
rect 119890 6128 119896 6180
rect 119948 6168 119954 6180
rect 251266 6168 251272 6180
rect 119948 6140 251272 6168
rect 119948 6128 119954 6140
rect 251266 6128 251272 6140
rect 251324 6128 251330 6180
rect 257062 6128 257068 6180
rect 257120 6168 257126 6180
rect 276290 6168 276296 6180
rect 257120 6140 276296 6168
rect 257120 6128 257126 6140
rect 276290 6128 276296 6140
rect 276348 6128 276354 6180
rect 286962 6128 286968 6180
rect 287020 6168 287026 6180
rect 415486 6168 415492 6180
rect 287020 6140 415492 6168
rect 287020 6128 287026 6140
rect 415486 6128 415492 6140
rect 415544 6128 415550 6180
rect 278314 5516 278320 5568
rect 278372 5556 278378 5568
rect 279418 5556 279424 5568
rect 278372 5528 279424 5556
rect 278372 5516 278378 5528
rect 279418 5516 279424 5528
rect 279476 5516 279482 5568
rect 284294 5176 284300 5228
rect 284352 5216 284358 5228
rect 298462 5216 298468 5228
rect 284352 5188 298468 5216
rect 284352 5176 284358 5188
rect 298462 5176 298468 5188
rect 298520 5176 298526 5228
rect 285766 5108 285772 5160
rect 285824 5148 285830 5160
rect 307938 5148 307944 5160
rect 285824 5120 307944 5148
rect 285824 5108 285830 5120
rect 307938 5108 307944 5120
rect 307996 5108 308002 5160
rect 294138 5040 294144 5092
rect 294196 5080 294202 5092
rect 350442 5080 350448 5092
rect 294196 5052 350448 5080
rect 294196 5040 294202 5052
rect 350442 5040 350448 5052
rect 350500 5040 350506 5092
rect 294230 4972 294236 5024
rect 294288 5012 294294 5024
rect 354030 5012 354036 5024
rect 294288 4984 354036 5012
rect 294288 4972 294294 4984
rect 354030 4972 354036 4984
rect 354088 4972 354094 5024
rect 296714 4904 296720 4956
rect 296772 4944 296778 4956
rect 364610 4944 364616 4956
rect 296772 4916 364616 4944
rect 296772 4904 296778 4916
rect 364610 4904 364616 4916
rect 364668 4904 364674 4956
rect 244090 4836 244096 4888
rect 244148 4876 244154 4888
rect 275186 4876 275192 4888
rect 244148 4848 275192 4876
rect 244148 4836 244154 4848
rect 275186 4836 275192 4848
rect 275244 4836 275250 4888
rect 298554 4836 298560 4888
rect 298612 4876 298618 4888
rect 371694 4876 371700 4888
rect 298612 4848 371700 4876
rect 298612 4836 298618 4848
rect 371694 4836 371700 4848
rect 371752 4836 371758 4888
rect 177850 4768 177856 4820
rect 177908 4808 177914 4820
rect 260098 4808 260104 4820
rect 177908 4780 260104 4808
rect 177908 4768 177914 4780
rect 260098 4768 260104 4780
rect 260156 4768 260162 4820
rect 264146 4768 264152 4820
rect 264204 4808 264210 4820
rect 277762 4808 277768 4820
rect 264204 4780 277768 4808
rect 264204 4768 264210 4780
rect 277762 4768 277768 4780
rect 277820 4768 277826 4820
rect 282914 4768 282920 4820
rect 282972 4808 282978 4820
rect 290182 4808 290188 4820
rect 282972 4780 290188 4808
rect 282972 4768 282978 4780
rect 290182 4768 290188 4780
rect 290240 4768 290246 4820
rect 299382 4768 299388 4820
rect 299440 4808 299446 4820
rect 377674 4808 377680 4820
rect 299440 4780 377680 4808
rect 299440 4768 299446 4780
rect 377674 4768 377680 4780
rect 377732 4768 377738 4820
rect 281718 4156 281724 4208
rect 281776 4196 281782 4208
rect 285398 4196 285404 4208
rect 281776 4168 285404 4196
rect 281776 4156 281782 4168
rect 285398 4156 285404 4168
rect 285456 4156 285462 4208
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 7558 4128 7564 4140
rect 2924 4100 7564 4128
rect 2924 4088 2930 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 46290 4128 46296 4140
rect 45520 4100 46296 4128
rect 45520 4088 45526 4100
rect 46290 4088 46296 4100
rect 46348 4088 46354 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 293310 4088 293316 4140
rect 293368 4128 293374 4140
rect 296070 4128 296076 4140
rect 293368 4100 296076 4128
rect 293368 4088 293374 4100
rect 296070 4088 296076 4100
rect 296128 4088 296134 4140
rect 349246 4128 349252 4140
rect 298204 4100 349252 4128
rect 239306 4020 239312 4072
rect 239364 4060 239370 4072
rect 253198 4060 253204 4072
rect 239364 4032 253204 4060
rect 239364 4020 239370 4032
rect 253198 4020 253204 4032
rect 253256 4020 253262 4072
rect 294046 4020 294052 4072
rect 294104 4060 294110 4072
rect 298204 4060 298232 4100
rect 349246 4088 349252 4100
rect 349304 4088 349310 4140
rect 430850 4088 430856 4140
rect 430908 4128 430914 4140
rect 437658 4128 437664 4140
rect 430908 4100 437664 4128
rect 430908 4088 430914 4100
rect 437658 4088 437664 4100
rect 437716 4088 437722 4140
rect 460198 4088 460204 4140
rect 460256 4128 460262 4140
rect 462774 4128 462780 4140
rect 460256 4100 462780 4128
rect 460256 4088 460262 4100
rect 462774 4088 462780 4100
rect 462832 4088 462838 4140
rect 468478 4088 468484 4140
rect 468536 4128 468542 4140
rect 471054 4128 471060 4140
rect 468536 4100 471060 4128
rect 468536 4088 468542 4100
rect 471054 4088 471060 4100
rect 471112 4088 471118 4140
rect 536190 4088 536196 4140
rect 536248 4128 536254 4140
rect 538398 4128 538404 4140
rect 536248 4100 538404 4128
rect 536248 4088 536254 4100
rect 538398 4088 538404 4100
rect 538456 4088 538462 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 569126 4128 569132 4140
rect 566516 4100 569132 4128
rect 566516 4088 566522 4100
rect 569126 4088 569132 4100
rect 569184 4088 569190 4140
rect 294104 4032 298232 4060
rect 294104 4020 294110 4032
rect 298278 4020 298284 4072
rect 298336 4060 298342 4072
rect 352834 4060 352840 4072
rect 298336 4032 352840 4060
rect 298336 4020 298342 4032
rect 352834 4020 352840 4032
rect 352892 4020 352898 4072
rect 429654 4020 429660 4072
rect 429712 4060 429718 4072
rect 438854 4060 438860 4072
rect 429712 4032 438860 4060
rect 429712 4020 429718 4032
rect 438854 4020 438860 4032
rect 438912 4020 438918 4072
rect 92750 3952 92756 4004
rect 92808 3992 92814 4004
rect 95878 3992 95884 4004
rect 92808 3964 95884 3992
rect 92808 3952 92814 3964
rect 95878 3952 95884 3964
rect 95936 3952 95942 4004
rect 135254 3952 135260 4004
rect 135312 3992 135318 4004
rect 136450 3992 136456 4004
rect 135312 3964 136456 3992
rect 135312 3952 135318 3964
rect 136450 3952 136456 3964
rect 136508 3952 136514 4004
rect 164878 3952 164884 4004
rect 164936 3992 164942 4004
rect 259454 3992 259460 4004
rect 164936 3964 259460 3992
rect 164936 3952 164942 3964
rect 259454 3952 259460 3964
rect 259512 3952 259518 4004
rect 273622 3952 273628 4004
rect 273680 3992 273686 4004
rect 279510 3992 279516 4004
rect 273680 3964 279516 3992
rect 273680 3952 273686 3964
rect 279510 3952 279516 3964
rect 279568 3952 279574 4004
rect 295334 3952 295340 4004
rect 295392 3992 295398 4004
rect 356330 3992 356336 4004
rect 295392 3964 298324 3992
rect 295392 3952 295398 3964
rect 110506 3884 110512 3936
rect 110564 3924 110570 3936
rect 113818 3924 113824 3936
rect 110564 3896 113824 3924
rect 110564 3884 110570 3896
rect 113818 3884 113824 3896
rect 113876 3884 113882 3936
rect 124674 3884 124680 3936
rect 124732 3924 124738 3936
rect 243630 3924 243636 3936
rect 124732 3896 243636 3924
rect 124732 3884 124738 3896
rect 243630 3884 243636 3896
rect 243688 3884 243694 3936
rect 293954 3884 293960 3936
rect 294012 3924 294018 3936
rect 298186 3924 298192 3936
rect 294012 3896 298192 3924
rect 294012 3884 294018 3896
rect 298186 3884 298192 3896
rect 298244 3884 298250 3936
rect 298296 3924 298324 3964
rect 298480 3964 356336 3992
rect 298480 3924 298508 3964
rect 356330 3952 356336 3964
rect 356388 3952 356394 4004
rect 428458 3952 428464 4004
rect 428516 3992 428522 4004
rect 439038 3992 439044 4004
rect 428516 3964 439044 3992
rect 428516 3952 428522 3964
rect 439038 3952 439044 3964
rect 439096 3952 439102 4004
rect 298296 3896 298508 3924
rect 298738 3884 298744 3936
rect 298796 3924 298802 3936
rect 365806 3924 365812 3936
rect 298796 3896 365812 3924
rect 298796 3884 298802 3896
rect 365806 3884 365812 3896
rect 365864 3884 365870 3936
rect 426158 3884 426164 3936
rect 426216 3924 426222 3936
rect 437566 3924 437572 3936
rect 426216 3896 437572 3924
rect 426216 3884 426222 3896
rect 437566 3884 437572 3896
rect 437624 3884 437630 3936
rect 476758 3884 476764 3936
rect 476816 3924 476822 3936
rect 480530 3924 480536 3936
rect 476816 3896 480536 3924
rect 476816 3884 476822 3896
rect 480530 3884 480536 3896
rect 480588 3884 480594 3936
rect 117590 3816 117596 3868
rect 117648 3856 117654 3868
rect 239398 3856 239404 3868
rect 117648 3828 239404 3856
rect 117648 3816 117654 3828
rect 239398 3816 239404 3828
rect 239456 3816 239462 3868
rect 245194 3816 245200 3868
rect 245252 3856 245258 3868
rect 255958 3856 255964 3868
rect 245252 3828 255964 3856
rect 245252 3816 245258 3828
rect 255958 3816 255964 3828
rect 256016 3816 256022 3868
rect 261478 3856 261484 3868
rect 258046 3828 261484 3856
rect 19426 3748 19432 3800
rect 19484 3788 19490 3800
rect 39298 3788 39304 3800
rect 19484 3760 39304 3788
rect 19484 3748 19490 3760
rect 39298 3748 39304 3760
rect 39356 3748 39362 3800
rect 102226 3748 102232 3800
rect 102284 3788 102290 3800
rect 248690 3788 248696 3800
rect 102284 3760 248696 3788
rect 102284 3748 102290 3760
rect 248690 3748 248696 3760
rect 248748 3748 248754 3800
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 46198 3720 46204 3732
rect 11204 3692 46204 3720
rect 11204 3680 11210 3692
rect 46198 3680 46204 3692
rect 46256 3680 46262 3732
rect 68278 3720 68284 3732
rect 55186 3692 68284 3720
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 50338 3652 50344 3664
rect 15988 3624 50344 3652
rect 15988 3612 15994 3624
rect 50338 3612 50344 3624
rect 50396 3612 50402 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 4798 3584 4804 3596
rect 1728 3556 4804 3584
rect 1728 3544 1734 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 10318 3584 10324 3596
rect 6886 3556 10324 3584
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 6886 3516 6914 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13078 3584 13084 3596
rect 12400 3556 13084 3584
rect 12400 3544 12406 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 55186 3584 55214 3692
rect 68278 3680 68284 3692
rect 68336 3680 68342 3732
rect 98638 3680 98644 3732
rect 98696 3720 98702 3732
rect 247402 3720 247408 3732
rect 98696 3692 247408 3720
rect 98696 3680 98702 3692
rect 247402 3680 247408 3692
rect 247460 3680 247466 3732
rect 64138 3652 64144 3664
rect 25372 3556 55214 3584
rect 55876 3624 64144 3652
rect 25372 3544 25378 3556
rect 4120 3488 6914 3516
rect 4120 3476 4126 3488
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8938 3516 8944 3528
rect 7708 3488 8944 3516
rect 7708 3476 7714 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 55876 3516 55904 3624
rect 64138 3612 64144 3624
rect 64196 3612 64202 3664
rect 74994 3612 75000 3664
rect 75052 3652 75058 3664
rect 88978 3652 88984 3664
rect 75052 3624 88984 3652
rect 75052 3612 75058 3624
rect 88978 3612 88984 3624
rect 89036 3612 89042 3664
rect 97442 3612 97448 3664
rect 97500 3652 97506 3664
rect 247218 3652 247224 3664
rect 97500 3624 247224 3652
rect 97500 3612 97506 3624
rect 247218 3612 247224 3624
rect 247276 3612 247282 3664
rect 251266 3612 251272 3664
rect 251324 3652 251330 3664
rect 258046 3652 258074 3828
rect 261478 3816 261484 3828
rect 261536 3816 261542 3868
rect 295426 3816 295432 3868
rect 295484 3856 295490 3868
rect 359918 3856 359924 3868
rect 295484 3828 359924 3856
rect 295484 3816 295490 3828
rect 359918 3816 359924 3828
rect 359976 3816 359982 3868
rect 427262 3816 427268 3868
rect 427320 3856 427326 3868
rect 439314 3856 439320 3868
rect 427320 3828 439320 3856
rect 427320 3816 427326 3828
rect 439314 3816 439320 3828
rect 439372 3816 439378 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 519538 3856 519544 3868
rect 516836 3828 519544 3856
rect 516836 3816 516842 3828
rect 519538 3816 519544 3828
rect 519596 3816 519602 3868
rect 574738 3816 574744 3868
rect 574796 3856 574802 3868
rect 577406 3856 577412 3868
rect 574796 3828 577412 3856
rect 574796 3816 574802 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 264330 3788 264336 3800
rect 251324 3624 258074 3652
rect 258184 3760 264336 3788
rect 251324 3612 251330 3624
rect 70302 3544 70308 3596
rect 70360 3584 70366 3596
rect 71038 3584 71044 3596
rect 70360 3556 71044 3584
rect 70360 3544 70366 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 82170 3584 82176 3596
rect 74506 3556 82176 3584
rect 20680 3488 55904 3516
rect 20680 3476 20686 3488
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 57238 3516 57244 3528
rect 56100 3488 57244 3516
rect 56100 3476 56106 3488
rect 57238 3476 57244 3488
rect 57296 3476 57302 3528
rect 60734 3476 60740 3528
rect 60792 3516 60798 3528
rect 61654 3516 61660 3528
rect 60792 3488 61660 3516
rect 60792 3476 60798 3488
rect 61654 3476 61660 3488
rect 61712 3476 61718 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66898 3516 66904 3528
rect 65576 3488 66904 3516
rect 65576 3476 65582 3488
rect 66898 3476 66904 3488
rect 66956 3476 66962 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 74506 3516 74534 3556
rect 82170 3544 82176 3556
rect 82228 3544 82234 3596
rect 96246 3544 96252 3596
rect 96304 3584 96310 3596
rect 97258 3584 97264 3596
rect 96304 3556 97264 3584
rect 96304 3544 96310 3556
rect 97258 3544 97264 3556
rect 97316 3544 97322 3596
rect 102134 3544 102140 3596
rect 102192 3584 102198 3596
rect 103330 3584 103336 3596
rect 102192 3556 103336 3584
rect 102192 3544 102198 3556
rect 103330 3544 103336 3556
rect 103388 3544 103394 3596
rect 103422 3544 103428 3596
rect 103480 3584 103486 3596
rect 247494 3584 247500 3596
rect 103480 3556 247500 3584
rect 103480 3544 103486 3556
rect 247494 3544 247500 3556
rect 247552 3544 247558 3596
rect 249978 3544 249984 3596
rect 250036 3584 250042 3596
rect 258184 3584 258212 3760
rect 264330 3748 264336 3760
rect 264388 3748 264394 3800
rect 288342 3748 288348 3800
rect 288400 3788 288406 3800
rect 367002 3788 367008 3800
rect 288400 3760 367008 3788
rect 288400 3748 288406 3760
rect 367002 3748 367008 3760
rect 367060 3748 367066 3800
rect 424962 3748 424968 3800
rect 425020 3788 425026 3800
rect 437474 3788 437480 3800
rect 425020 3760 437480 3788
rect 425020 3748 425026 3760
rect 437474 3748 437480 3760
rect 437532 3748 437538 3800
rect 259454 3680 259460 3732
rect 259512 3720 259518 3732
rect 269758 3720 269764 3732
rect 259512 3692 269764 3720
rect 259512 3680 259518 3692
rect 269758 3680 269764 3692
rect 269816 3680 269822 3732
rect 295242 3680 295248 3732
rect 295300 3720 295306 3732
rect 384758 3720 384764 3732
rect 295300 3692 384764 3720
rect 295300 3680 295306 3692
rect 384758 3680 384764 3692
rect 384816 3680 384822 3732
rect 423766 3680 423772 3732
rect 423824 3720 423830 3732
rect 437842 3720 437848 3732
rect 423824 3692 437848 3720
rect 423824 3680 423830 3692
rect 437842 3680 437848 3692
rect 437900 3680 437906 3732
rect 295150 3612 295156 3664
rect 295208 3652 295214 3664
rect 402514 3652 402520 3664
rect 295208 3624 402520 3652
rect 295208 3612 295214 3624
rect 402514 3612 402520 3624
rect 402572 3612 402578 3664
rect 422570 3612 422576 3664
rect 422628 3652 422634 3664
rect 438946 3652 438952 3664
rect 422628 3624 438952 3652
rect 422628 3612 422634 3624
rect 438946 3612 438952 3624
rect 439004 3612 439010 3664
rect 250036 3556 258212 3584
rect 250036 3544 250042 3556
rect 258258 3544 258264 3596
rect 258316 3584 258322 3596
rect 260190 3584 260196 3596
rect 258316 3556 260196 3584
rect 258316 3544 258322 3556
rect 260190 3544 260196 3556
rect 260248 3544 260254 3596
rect 267918 3544 267924 3596
rect 267976 3584 267982 3596
rect 268470 3584 268476 3596
rect 267976 3556 268476 3584
rect 267976 3544 267982 3556
rect 268470 3544 268476 3556
rect 268528 3544 268534 3596
rect 271138 3584 271144 3596
rect 269408 3556 271144 3584
rect 67968 3488 74534 3516
rect 67968 3476 67974 3488
rect 77294 3476 77300 3528
rect 77352 3516 77358 3528
rect 78214 3516 78220 3528
rect 77352 3488 78220 3516
rect 77352 3476 77358 3488
rect 78214 3476 78220 3488
rect 78272 3476 78278 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 244366 3516 244372 3528
rect 83332 3488 244372 3516
rect 83332 3476 83338 3488
rect 244366 3476 244372 3488
rect 244424 3476 244430 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252370 3516 252376 3528
rect 251232 3488 252376 3516
rect 251232 3476 251238 3488
rect 252370 3476 252376 3488
rect 252428 3476 252434 3528
rect 253474 3476 253480 3528
rect 253532 3516 253538 3528
rect 269408 3516 269436 3556
rect 271138 3544 271144 3556
rect 271196 3544 271202 3596
rect 286318 3544 286324 3596
rect 286376 3584 286382 3596
rect 297266 3584 297272 3596
rect 286376 3556 297272 3584
rect 286376 3544 286382 3556
rect 297266 3544 297272 3556
rect 297324 3544 297330 3596
rect 298002 3544 298008 3596
rect 298060 3584 298066 3596
rect 406010 3584 406016 3596
rect 298060 3556 406016 3584
rect 298060 3544 298066 3556
rect 406010 3544 406016 3556
rect 406068 3544 406074 3596
rect 421374 3544 421380 3596
rect 421432 3584 421438 3596
rect 434346 3584 434352 3596
rect 421432 3556 434352 3584
rect 421432 3544 421438 3556
rect 434346 3544 434352 3556
rect 434404 3544 434410 3596
rect 434438 3544 434444 3596
rect 434496 3584 434502 3596
rect 439130 3584 439136 3596
rect 434496 3556 439136 3584
rect 434496 3544 434502 3556
rect 439130 3544 439136 3556
rect 439188 3544 439194 3596
rect 442350 3544 442356 3596
rect 442408 3584 442414 3596
rect 447410 3584 447416 3596
rect 442408 3556 447416 3584
rect 442408 3544 442414 3556
rect 447410 3544 447416 3556
rect 447468 3544 447474 3596
rect 450538 3544 450544 3596
rect 450596 3584 450602 3596
rect 450596 3556 451274 3584
rect 450596 3544 450602 3556
rect 253532 3488 269436 3516
rect 253532 3476 253538 3488
rect 270034 3476 270040 3528
rect 270092 3516 270098 3528
rect 271230 3516 271236 3528
rect 270092 3488 271236 3516
rect 270092 3476 270098 3488
rect 271230 3476 271236 3488
rect 271288 3476 271294 3528
rect 272426 3476 272432 3528
rect 272484 3516 272490 3528
rect 273898 3516 273904 3528
rect 272484 3488 273904 3516
rect 272484 3476 272490 3488
rect 273898 3476 273904 3488
rect 273956 3476 273962 3528
rect 293862 3476 293868 3528
rect 293920 3516 293926 3528
rect 409598 3516 409604 3528
rect 293920 3488 409604 3516
rect 293920 3476 293926 3488
rect 409598 3476 409604 3488
rect 409656 3476 409662 3528
rect 418982 3476 418988 3528
rect 419040 3516 419046 3528
rect 438026 3516 438032 3528
rect 419040 3488 438032 3516
rect 419040 3476 419046 3488
rect 438026 3476 438032 3488
rect 438084 3476 438090 3528
rect 440326 3476 440332 3528
rect 440384 3516 440390 3528
rect 441522 3516 441528 3528
rect 440384 3488 441528 3516
rect 440384 3476 440390 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 448606 3476 448612 3528
rect 448664 3516 448670 3528
rect 449802 3516 449808 3528
rect 448664 3488 449808 3516
rect 448664 3476 448670 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 451246 3516 451274 3556
rect 453298 3544 453304 3596
rect 453356 3584 453362 3596
rect 455690 3584 455696 3596
rect 453356 3556 455696 3584
rect 453356 3544 453362 3556
rect 455690 3544 455696 3556
rect 455748 3544 455754 3596
rect 458818 3544 458824 3596
rect 458876 3584 458882 3596
rect 465166 3584 465172 3596
rect 458876 3556 465172 3584
rect 458876 3544 458882 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 469858 3584 469864 3596
rect 467156 3556 469864 3584
rect 467156 3544 467162 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 470566 3556 475240 3584
rect 454494 3516 454500 3528
rect 451246 3488 454500 3516
rect 454494 3476 454500 3488
rect 454552 3476 454558 3528
rect 456886 3476 456892 3528
rect 456944 3516 456950 3528
rect 458082 3516 458088 3528
rect 456944 3488 458088 3516
rect 456944 3476 456950 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 462958 3476 462964 3528
rect 463016 3516 463022 3528
rect 470566 3516 470594 3556
rect 463016 3488 470594 3516
rect 463016 3476 463022 3488
rect 471238 3476 471244 3528
rect 471296 3516 471302 3528
rect 473446 3516 473452 3528
rect 471296 3488 473452 3516
rect 471296 3476 471302 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 475212 3516 475240 3556
rect 475378 3544 475384 3596
rect 475436 3584 475442 3596
rect 476942 3584 476948 3596
rect 475436 3556 476948 3584
rect 475436 3544 475442 3556
rect 476942 3544 476948 3556
rect 477000 3544 477006 3596
rect 478230 3544 478236 3596
rect 478288 3584 478294 3596
rect 484026 3584 484032 3596
rect 478288 3556 484032 3584
rect 478288 3544 478294 3556
rect 484026 3544 484032 3556
rect 484084 3544 484090 3596
rect 500218 3544 500224 3596
rect 500276 3584 500282 3596
rect 501782 3584 501788 3596
rect 500276 3556 501788 3584
rect 500276 3544 500282 3556
rect 501782 3544 501788 3556
rect 501840 3544 501846 3596
rect 548518 3544 548524 3596
rect 548576 3584 548582 3596
rect 550266 3584 550272 3596
rect 548576 3556 550272 3584
rect 548576 3544 548582 3556
rect 550266 3544 550272 3556
rect 550324 3544 550330 3596
rect 479334 3516 479340 3528
rect 475212 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 496078 3476 496084 3528
rect 496136 3516 496142 3528
rect 497090 3516 497096 3528
rect 496136 3488 497096 3516
rect 496136 3476 496142 3488
rect 497090 3476 497096 3488
rect 497148 3476 497154 3528
rect 514018 3476 514024 3528
rect 514076 3516 514082 3528
rect 515950 3516 515956 3528
rect 514076 3488 515956 3516
rect 514076 3476 514082 3488
rect 515950 3476 515956 3488
rect 516008 3476 516014 3528
rect 522298 3476 522304 3528
rect 522356 3516 522362 3528
rect 524230 3516 524236 3528
rect 522356 3488 524236 3516
rect 522356 3476 522362 3488
rect 524230 3476 524236 3488
rect 524288 3476 524294 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 540790 3516 540796 3528
rect 538916 3488 540796 3516
rect 538916 3476 538922 3488
rect 540790 3476 540796 3488
rect 540848 3476 540854 3528
rect 549898 3476 549904 3528
rect 549956 3516 549962 3528
rect 551462 3516 551468 3528
rect 549956 3488 551468 3516
rect 549956 3476 549962 3488
rect 551462 3476 551468 3488
rect 551520 3476 551526 3528
rect 563698 3476 563704 3528
rect 563756 3516 563762 3528
rect 566826 3516 566832 3528
rect 563756 3488 566832 3516
rect 563756 3476 563762 3488
rect 566826 3476 566832 3488
rect 566884 3476 566890 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 581822 3516 581828 3528
rect 581052 3488 581828 3516
rect 581052 3476 581058 3488
rect 581822 3476 581828 3488
rect 581880 3476 581886 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 25498 3448 25504 3460
rect 624 3420 25504 3448
rect 624 3408 630 3420
rect 25498 3408 25504 3420
rect 25556 3408 25562 3460
rect 27614 3408 27620 3460
rect 27672 3448 27678 3460
rect 28534 3448 28540 3460
rect 27672 3420 28540 3448
rect 27672 3408 27678 3420
rect 28534 3408 28540 3420
rect 28592 3408 28598 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 35158 3448 35164 3460
rect 33652 3420 35164 3448
rect 33652 3408 33658 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 39390 3448 39396 3460
rect 38436 3420 39396 3448
rect 38436 3408 38442 3420
rect 39390 3408 39396 3420
rect 39448 3408 39454 3460
rect 39574 3408 39580 3460
rect 39632 3448 39638 3460
rect 43438 3448 43444 3460
rect 39632 3420 43444 3448
rect 39632 3408 39638 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 46658 3408 46664 3460
rect 46716 3448 46722 3460
rect 47578 3448 47584 3460
rect 46716 3420 47584 3448
rect 46716 3408 46722 3420
rect 47578 3408 47584 3420
rect 47636 3408 47642 3460
rect 47854 3408 47860 3460
rect 47912 3448 47918 3460
rect 48958 3448 48964 3460
rect 47912 3420 48964 3448
rect 47912 3408 47918 3420
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 79686 3408 79692 3460
rect 79744 3448 79750 3460
rect 244550 3448 244556 3460
rect 79744 3420 244556 3448
rect 79744 3408 79750 3420
rect 244550 3408 244556 3420
rect 244608 3408 244614 3460
rect 246390 3408 246396 3460
rect 246448 3448 246454 3460
rect 246448 3420 258074 3448
rect 246448 3408 246454 3420
rect 95142 3340 95148 3392
rect 95200 3380 95206 3392
rect 103422 3380 103428 3392
rect 95200 3352 103428 3380
rect 95200 3340 95206 3352
rect 103422 3340 103428 3352
rect 103480 3340 103486 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 258046 3380 258074 3420
rect 285582 3408 285588 3460
rect 285640 3448 285646 3460
rect 401318 3448 401324 3460
rect 285640 3420 401324 3448
rect 285640 3408 285646 3420
rect 401318 3408 401324 3420
rect 401376 3408 401382 3460
rect 417878 3408 417884 3460
rect 417936 3448 417942 3460
rect 437750 3448 437756 3460
rect 417936 3420 437756 3448
rect 417936 3408 417942 3420
rect 437750 3408 437756 3420
rect 437808 3408 437814 3460
rect 445110 3408 445116 3460
rect 445168 3448 445174 3460
rect 445168 3420 509234 3448
rect 445168 3408 445174 3420
rect 265618 3380 265624 3392
rect 258046 3352 265624 3380
rect 265618 3340 265624 3352
rect 265676 3340 265682 3392
rect 285674 3340 285680 3392
rect 285732 3380 285738 3392
rect 309042 3380 309048 3392
rect 285732 3352 309048 3380
rect 285732 3340 285738 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332686 3340 332692 3392
rect 332744 3380 332750 3392
rect 333882 3380 333888 3392
rect 332744 3352 333888 3380
rect 332744 3340 332750 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 434346 3340 434352 3392
rect 434404 3380 434410 3392
rect 439222 3380 439228 3392
rect 434404 3352 439228 3380
rect 434404 3340 434410 3352
rect 439222 3340 439228 3352
rect 439280 3340 439286 3392
rect 446398 3340 446404 3392
rect 446456 3380 446462 3392
rect 452102 3380 452108 3392
rect 446456 3352 452108 3380
rect 446456 3340 446462 3352
rect 452102 3340 452108 3352
rect 452160 3340 452166 3392
rect 493318 3340 493324 3392
rect 493376 3380 493382 3392
rect 499390 3380 499396 3392
rect 493376 3352 499396 3380
rect 493376 3340 493382 3352
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 509206 3380 509234 3420
rect 514110 3408 514116 3460
rect 514168 3448 514174 3460
rect 514754 3448 514760 3460
rect 514168 3420 514760 3448
rect 514168 3408 514174 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 520918 3408 520924 3460
rect 520976 3448 520982 3460
rect 523034 3448 523040 3460
rect 520976 3420 523040 3448
rect 520976 3408 520982 3420
rect 523034 3408 523040 3420
rect 523092 3408 523098 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 533706 3448 533712 3460
rect 527968 3420 533712 3448
rect 527968 3408 527974 3420
rect 533706 3408 533712 3420
rect 533764 3408 533770 3460
rect 542998 3408 543004 3460
rect 543056 3448 543062 3460
rect 549070 3448 549076 3460
rect 543056 3420 549076 3448
rect 543056 3408 543062 3420
rect 549070 3408 549076 3420
rect 549128 3408 549134 3460
rect 526622 3380 526628 3392
rect 509206 3352 526628 3380
rect 526622 3340 526628 3352
rect 526680 3340 526686 3392
rect 554038 3340 554044 3392
rect 554096 3380 554102 3392
rect 559742 3380 559748 3392
rect 554096 3352 559748 3380
rect 554096 3340 554102 3352
rect 559742 3340 559748 3352
rect 559800 3340 559806 3392
rect 262950 3272 262956 3324
rect 263008 3312 263014 3324
rect 264422 3312 264428 3324
rect 263008 3284 264428 3312
rect 263008 3272 263014 3284
rect 264422 3272 264428 3284
rect 264480 3272 264486 3324
rect 454678 3272 454684 3324
rect 454736 3312 454742 3324
rect 459186 3312 459192 3324
rect 454736 3284 459192 3312
rect 454736 3272 454742 3284
rect 459186 3272 459192 3284
rect 459244 3272 459250 3324
rect 509878 3272 509884 3324
rect 509936 3312 509942 3324
rect 513558 3312 513564 3324
rect 509936 3284 513564 3312
rect 509936 3272 509942 3284
rect 513558 3272 513564 3284
rect 513616 3272 513622 3324
rect 571978 3272 571984 3324
rect 572036 3312 572042 3324
rect 573910 3312 573916 3324
rect 572036 3284 573916 3312
rect 572036 3272 572042 3284
rect 573910 3272 573916 3284
rect 573968 3272 573974 3324
rect 6454 3204 6460 3256
rect 6512 3244 6518 3256
rect 7558 3244 7564 3256
rect 6512 3216 7564 3244
rect 6512 3204 6518 3216
rect 7558 3204 7564 3216
rect 7616 3204 7622 3256
rect 51350 3204 51356 3256
rect 51408 3244 51414 3256
rect 53098 3244 53104 3256
rect 51408 3216 53104 3244
rect 51408 3204 51414 3216
rect 53098 3204 53104 3216
rect 53156 3204 53162 3256
rect 85666 3136 85672 3188
rect 85724 3176 85730 3188
rect 93118 3176 93124 3188
rect 85724 3148 93124 3176
rect 85724 3136 85730 3148
rect 93118 3136 93124 3148
rect 93176 3136 93182 3188
rect 114002 3136 114008 3188
rect 114060 3176 114066 3188
rect 117958 3176 117964 3188
rect 114060 3148 117964 3176
rect 114060 3136 114066 3148
rect 117958 3136 117964 3148
rect 118016 3136 118022 3188
rect 277118 3136 277124 3188
rect 277176 3176 277182 3188
rect 278130 3176 278136 3188
rect 277176 3148 278136 3176
rect 277176 3136 277182 3148
rect 278130 3136 278136 3148
rect 278188 3136 278194 3188
rect 281626 3136 281632 3188
rect 281684 3176 281690 3188
rect 284294 3176 284300 3188
rect 281684 3148 284300 3176
rect 281684 3136 281690 3148
rect 284294 3136 284300 3148
rect 284352 3136 284358 3188
rect 485038 3136 485044 3188
rect 485096 3176 485102 3188
rect 487614 3176 487620 3188
rect 485096 3148 487620 3176
rect 485096 3136 485102 3148
rect 487614 3136 487620 3148
rect 487672 3136 487678 3188
rect 534718 3136 534724 3188
rect 534776 3176 534782 3188
rect 537202 3176 537208 3188
rect 534776 3148 537208 3176
rect 534776 3136 534782 3148
rect 537202 3136 537208 3148
rect 537260 3136 537266 3188
rect 560938 3136 560944 3188
rect 560996 3176 561002 3188
rect 563238 3176 563244 3188
rect 560996 3148 563244 3176
rect 560996 3136 561002 3148
rect 563238 3136 563244 3148
rect 563296 3136 563302 3188
rect 567838 3136 567844 3188
rect 567896 3176 567902 3188
rect 570322 3176 570328 3188
rect 567896 3148 570328 3176
rect 567896 3136 567902 3148
rect 570322 3136 570328 3148
rect 570380 3136 570386 3188
rect 570598 3068 570604 3120
rect 570656 3108 570662 3120
rect 572714 3108 572720 3120
rect 570656 3080 572720 3108
rect 570656 3068 570662 3080
rect 572714 3068 572720 3080
rect 572772 3068 572778 3120
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 503070 3000 503076 3052
rect 503128 3040 503134 3052
rect 505370 3040 505376 3052
rect 503128 3012 505376 3040
rect 503128 3000 503134 3012
rect 505370 3000 505376 3012
rect 505428 3000 505434 3052
rect 552750 3000 552756 3052
rect 552808 3040 552814 3052
rect 554958 3040 554964 3052
rect 552808 3012 554964 3040
rect 552808 3000 552814 3012
rect 554958 3000 554964 3012
rect 555016 3000 555022 3052
rect 563790 3000 563796 3052
rect 563848 3040 563854 3052
rect 565630 3040 565636 3052
rect 563848 3012 565636 3040
rect 563848 3000 563854 3012
rect 565630 3000 565636 3012
rect 565688 3000 565694 3052
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 14458 2972 14464 2984
rect 8812 2944 14464 2972
rect 8812 2932 8818 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 526530 2932 526536 2984
rect 526588 2972 526594 2984
rect 527818 2972 527824 2984
rect 526588 2944 527824 2972
rect 526588 2932 526594 2944
rect 527818 2932 527824 2944
rect 527876 2932 527882 2984
rect 540238 2932 540244 2984
rect 540296 2972 540302 2984
rect 541986 2972 541992 2984
rect 540296 2944 541992 2972
rect 540296 2932 540302 2944
rect 541986 2932 541992 2944
rect 542044 2932 542050 2984
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 348792 700544 348844 700596
rect 357624 700544 357676 700596
rect 332508 700476 332560 700528
rect 358820 700476 358872 700528
rect 300124 700408 300176 700460
rect 357532 700408 357584 700460
rect 283840 700340 283892 700392
rect 358912 700340 358964 700392
rect 8116 700272 8168 700324
rect 21364 700272 21416 700324
rect 217968 700272 218020 700324
rect 235172 700272 235224 700324
rect 267648 700272 267700 700324
rect 357440 700272 357492 700324
rect 359464 700272 359516 700324
rect 397460 700272 397512 700324
rect 467104 700272 467156 700324
rect 527180 700272 527232 700324
rect 527824 700272 527876 700324
rect 559656 700272 559708 700324
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 371884 696940 371936 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 3516 670692 3568 670744
rect 18604 670692 18656 670744
rect 360844 670692 360896 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 17224 656888 17276 656940
rect 367744 643084 367796 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 13084 632068 13136 632120
rect 373264 630640 373316 630692
rect 579988 630640 580040 630692
rect 378784 616836 378836 616888
rect 580172 616836 580224 616888
rect 3516 606024 3568 606076
rect 7564 606024 7616 606076
rect 363604 590656 363656 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 10324 579640 10376 579692
rect 369124 576852 369176 576904
rect 580172 576852 580224 576904
rect 381544 563048 381596 563100
rect 580172 563048 580224 563100
rect 3608 553392 3660 553444
rect 22744 553392 22796 553444
rect 498844 536800 498896 536852
rect 579896 536800 579948 536852
rect 2964 527144 3016 527196
rect 14464 527144 14516 527196
rect 3332 501304 3384 501356
rect 8944 501304 8996 501356
rect 480904 484372 480956 484424
rect 580172 484372 580224 484424
rect 217324 478864 217376 478916
rect 220084 478864 220136 478916
rect 219072 478252 219124 478304
rect 238760 478252 238812 478304
rect 217600 478184 217652 478236
rect 248512 478184 248564 478236
rect 309140 478184 309192 478236
rect 357624 478184 357676 478236
rect 218060 478116 218112 478168
rect 314752 478116 314804 478168
rect 245752 476960 245804 477012
rect 247040 476960 247092 477012
rect 258080 476960 258132 477012
rect 262220 476960 262272 477012
rect 217508 476756 217560 476808
rect 230480 476756 230532 476808
rect 233240 476688 233292 476740
rect 242900 476688 242952 476740
rect 247316 476688 247368 476740
rect 248420 476688 248472 476740
rect 258080 476688 258132 476740
rect 258724 476688 258776 476740
rect 291200 476688 291252 476740
rect 325792 476688 325844 476740
rect 278780 476620 278832 476672
rect 305000 476620 305052 476672
rect 240140 476552 240192 476604
rect 252560 476552 252612 476604
rect 252652 476552 252704 476604
rect 264980 476552 265032 476604
rect 280160 476552 280212 476604
rect 307760 476552 307812 476604
rect 233332 476484 233384 476536
rect 247040 476484 247092 476536
rect 248512 476484 248564 476536
rect 260840 476484 260892 476536
rect 260932 476484 260984 476536
rect 277952 476484 278004 476536
rect 281540 476484 281592 476536
rect 310520 476484 310572 476536
rect 237472 476416 237524 476468
rect 239128 476416 239180 476468
rect 241428 476416 241480 476468
rect 244280 476416 244332 476468
rect 255320 476416 255372 476468
rect 268016 476416 268068 476468
rect 282920 476416 282972 476468
rect 313280 476416 313332 476468
rect 231860 476280 231912 476332
rect 236000 476280 236052 476332
rect 236184 476280 236236 476332
rect 249800 476348 249852 476400
rect 251272 476348 251324 476400
rect 263600 476348 263652 476400
rect 284300 476348 284352 476400
rect 314660 476348 314712 476400
rect 242900 476280 242952 476332
rect 236092 476212 236144 476264
rect 234620 476144 234672 476196
rect 237380 476144 237432 476196
rect 238852 476212 238904 476264
rect 244648 476212 244700 476264
rect 256792 476280 256844 476332
rect 270500 476280 270552 476332
rect 285680 476280 285732 476332
rect 317420 476280 317472 476332
rect 255412 476212 255464 476264
rect 258172 476212 258224 476264
rect 273260 476212 273312 476264
rect 288440 476212 288492 476264
rect 320180 476212 320232 476264
rect 241428 476144 241480 476196
rect 241520 476144 241572 476196
rect 245660 476144 245712 476196
rect 252376 476144 252428 476196
rect 253940 476144 253992 476196
rect 259552 476144 259604 476196
rect 276020 476144 276072 476196
rect 289820 476144 289872 476196
rect 322940 476144 322992 476196
rect 234712 476076 234764 476128
rect 236000 476076 236052 476128
rect 236000 475940 236052 475992
rect 236184 476076 236236 476128
rect 242808 476076 242860 476128
rect 244280 476076 244332 476128
rect 245844 476076 245896 476128
rect 258264 476076 258316 476128
rect 277584 476076 277636 476128
rect 302240 476076 302292 476128
rect 219164 475328 219216 475380
rect 247132 475328 247184 475380
rect 267556 475328 267608 475380
rect 274640 475328 274692 475380
rect 301044 475328 301096 475380
rect 580264 475328 580316 475380
rect 3332 474716 3384 474768
rect 331220 474716 331272 474768
rect 217784 474036 217836 474088
rect 250444 474036 250496 474088
rect 276020 474036 276072 474088
rect 300860 474036 300912 474088
rect 320180 474036 320232 474088
rect 498844 474036 498896 474088
rect 21364 473968 21416 474020
rect 347872 473968 347924 474020
rect 217876 472676 217928 472728
rect 254032 472676 254084 472728
rect 269212 472676 269264 472728
rect 289912 472676 289964 472728
rect 71780 472608 71832 472660
rect 346492 472608 346544 472660
rect 298100 471316 298152 471368
rect 373264 471316 373316 471368
rect 14464 471248 14516 471300
rect 328460 471248 328512 471300
rect 267740 469888 267792 469940
rect 287060 469888 287112 469940
rect 10324 469820 10376 469872
rect 327080 469820 327132 469872
rect 334072 469820 334124 469872
rect 359464 469820 359516 469872
rect 266452 468528 266504 468580
rect 285772 468528 285824 468580
rect 13084 468460 13136 468512
rect 324320 468460 324372 468512
rect 329840 468460 329892 468512
rect 467104 468460 467156 468512
rect 295340 467168 295392 467220
rect 369124 467168 369176 467220
rect 4804 467100 4856 467152
rect 321560 467100 321612 467152
rect 169760 465672 169812 465724
rect 314752 465672 314804 465724
rect 327172 465672 327224 465724
rect 371884 465672 371936 465724
rect 305000 464380 305052 464432
rect 428464 464380 428516 464432
rect 22744 464312 22796 464364
rect 351920 464312 351972 464364
rect 271880 462952 271932 463004
rect 295432 462952 295484 463004
rect 332600 462952 332652 463004
rect 462320 462952 462372 463004
rect 3332 462340 3384 462392
rect 332692 462340 332744 462392
rect 273168 461728 273220 461780
rect 280344 461728 280396 461780
rect 277308 461660 277360 461712
rect 287060 461660 287112 461712
rect 219256 461592 219308 461644
rect 241612 461592 241664 461644
rect 263692 461592 263744 461644
rect 280252 461592 280304 461644
rect 317420 461592 317472 461644
rect 480904 461592 480956 461644
rect 322940 460232 322992 460284
rect 363604 460232 363656 460284
rect 17224 460164 17276 460216
rect 350080 460164 350132 460216
rect 308128 458872 308180 458924
rect 364340 458872 364392 458924
rect 7564 458804 7616 458856
rect 350816 458804 350868 458856
rect 303620 457512 303672 457564
rect 494060 457512 494112 457564
rect 8944 457444 8996 457496
rect 352288 457444 352340 457496
rect 270960 456084 271012 456136
rect 292580 456084 292632 456136
rect 300952 456084 301004 456136
rect 527824 456084 527876 456136
rect 18604 456016 18656 456068
rect 323584 456016 323636 456068
rect 269028 455336 269080 455388
rect 276480 455336 276532 455388
rect 274456 454724 274508 454776
rect 283012 454724 283064 454776
rect 278688 454656 278740 454708
rect 288808 454656 288860 454708
rect 298928 454656 298980 454708
rect 360844 454656 360896 454708
rect 274088 453364 274140 453416
rect 298192 453364 298244 453416
rect 217692 453296 217744 453348
rect 231952 453296 232004 453348
rect 267648 453296 267700 453348
rect 273260 453296 273312 453348
rect 275928 453296 275980 453348
rect 285772 453296 285824 453348
rect 296720 453296 296772 453348
rect 378784 453296 378836 453348
rect 271788 452752 271840 452804
rect 279424 452752 279476 452804
rect 270408 451936 270460 451988
rect 277492 451936 277544 451988
rect 280068 451936 280120 451988
rect 290280 451936 290332 451988
rect 219348 451868 219400 451920
rect 244648 451868 244700 451920
rect 266268 451868 266320 451920
rect 271972 451868 272024 451920
rect 274548 451868 274600 451920
rect 284392 451868 284444 451920
rect 294144 451868 294196 451920
rect 381544 451868 381596 451920
rect 265164 450576 265216 450628
rect 283104 450576 283156 450628
rect 325608 450576 325660 450628
rect 367744 450576 367796 450628
rect 3608 450508 3660 450560
rect 331036 450508 331088 450560
rect 307852 449624 307904 449676
rect 412640 449624 412692 449676
rect 153200 449556 153252 449608
rect 317144 449556 317196 449608
rect 305460 449488 305512 449540
rect 477500 449488 477552 449540
rect 88340 449420 88392 449472
rect 319444 449420 319496 449472
rect 303160 449352 303212 449404
rect 542360 449352 542412 449404
rect 23480 449284 23532 449336
rect 321744 449284 321796 449336
rect 3424 449216 3476 449268
rect 326436 449216 326488 449268
rect 3516 449148 3568 449200
rect 328736 449148 328788 449200
rect 201500 448060 201552 448112
rect 341892 448060 341944 448112
rect 136640 447992 136692 448044
rect 344192 447992 344244 448044
rect 104900 447924 104952 447976
rect 317880 447924 317932 447976
rect 40040 447856 40092 447908
rect 320180 447856 320232 447908
rect 2872 447788 2924 447840
rect 353484 447788 353536 447840
rect 255964 447040 256016 447092
rect 258264 447040 258316 447092
rect 262864 447040 262916 447092
rect 267556 447040 267608 447092
rect 231860 446972 231912 447024
rect 232412 446972 232464 447024
rect 236000 446972 236052 447024
rect 237012 446972 237064 447024
rect 241520 446972 241572 447024
rect 242348 446972 242400 447024
rect 248420 446972 248472 447024
rect 249340 446972 249392 447024
rect 250444 446972 250496 447024
rect 252008 446972 252060 447024
rect 253940 446972 253992 447024
rect 254860 446972 254912 447024
rect 256608 446972 256660 447024
rect 259736 446972 259788 447024
rect 261484 446972 261536 447024
rect 265992 446972 266044 447024
rect 271880 446972 271932 447024
rect 272708 446972 272760 447024
rect 277492 446972 277544 447024
rect 278044 446972 278096 447024
rect 282920 446972 282972 447024
rect 283380 446972 283432 447024
rect 284300 446972 284352 447024
rect 285036 446972 285088 447024
rect 285680 446972 285732 447024
rect 286508 446972 286560 447024
rect 300952 446972 301004 447024
rect 301228 446972 301280 447024
rect 264244 446904 264296 446956
rect 269120 446904 269172 446956
rect 217968 446632 218020 446684
rect 313188 446632 313240 446684
rect 339592 446632 339644 446684
rect 357440 446632 357492 446684
rect 260748 446564 260800 446616
rect 264428 446564 264480 446616
rect 302424 446564 302476 446616
rect 333980 446564 334032 446616
rect 337200 446564 337252 446616
rect 358820 446564 358872 446616
rect 312452 446496 312504 446548
rect 358912 446496 358964 446548
rect 220084 446428 220136 446480
rect 230388 446428 230440 446480
rect 265624 446428 265676 446480
rect 270592 446428 270644 446480
rect 310888 446428 310940 446480
rect 357532 446428 357584 446480
rect 311716 446360 311768 446412
rect 362224 446360 362276 446412
rect 307024 446292 307076 446344
rect 364984 446292 365036 446344
rect 253848 446224 253900 446276
rect 256700 446224 256752 446276
rect 258724 446224 258776 446276
rect 261300 446224 261352 446276
rect 304724 446224 304776 446276
rect 363604 446224 363656 446276
rect 293132 446156 293184 446208
rect 361028 446156 361080 446208
rect 292304 446088 292356 446140
rect 373264 446088 373316 446140
rect 243544 446020 243596 446072
rect 345020 446020 345072 446072
rect 229836 445952 229888 446004
rect 338028 445952 338080 446004
rect 229744 445884 229796 445936
rect 347320 445884 347372 445936
rect 228364 445816 228416 445868
rect 349620 445816 349672 445868
rect 293868 445748 293920 445800
rect 458824 445748 458876 445800
rect 228548 445204 228600 445256
rect 336464 445204 336516 445256
rect 7564 445136 7616 445188
rect 334164 445136 334216 445188
rect 225696 445068 225748 445120
rect 338764 445068 338816 445120
rect 333980 445000 334032 445052
rect 580264 445000 580316 445052
rect 224224 444932 224276 444984
rect 341156 444932 341208 444984
rect 228456 444864 228508 444916
rect 355876 444864 355928 444916
rect 300032 444796 300084 444848
rect 442264 444796 442316 444848
rect 295432 444728 295484 444780
rect 526444 444728 526496 444780
rect 93216 444660 93268 444712
rect 343456 444660 343508 444712
rect 86224 444592 86276 444644
rect 345756 444592 345808 444644
rect 84844 444524 84896 444576
rect 348056 444524 348108 444576
rect 82084 444456 82136 444508
rect 358176 444456 358228 444508
rect 314016 444388 314068 444440
rect 369124 444388 369176 444440
rect 3516 443640 3568 443692
rect 243544 443640 243596 443692
rect 309324 443640 309376 443692
rect 316316 443572 316368 443624
rect 362316 443572 362368 443624
rect 367744 443504 367796 443556
rect 226984 443436 227036 443488
rect 335544 443436 335596 443488
rect 225604 443368 225656 443420
rect 342260 443368 342312 443420
rect 221464 443300 221516 443352
rect 340052 443300 340104 443352
rect 228640 443232 228692 443284
rect 354036 443232 354088 443284
rect 220084 443164 220136 443216
rect 354772 443164 354824 443216
rect 98644 443096 98696 443148
rect 356244 443096 356296 443148
rect 95976 443028 96028 443080
rect 356980 443028 357032 443080
rect 80704 442960 80756 443012
rect 358820 442960 358872 443012
rect 3608 442212 3660 442264
rect 229836 442212 229888 442264
rect 361028 442212 361080 442264
rect 581000 442212 581052 442264
rect 3424 440852 3476 440904
rect 229744 440852 229796 440904
rect 458824 439492 458876 439544
rect 582380 439492 582432 439544
rect 362316 431876 362368 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 7564 423580 7616 423632
rect 3332 411204 3384 411256
rect 226984 411204 227036 411256
rect 3332 398760 3384 398812
rect 228640 398760 228692 398812
rect 369124 379448 369176 379500
rect 580172 379448 580224 379500
rect 3056 372512 3108 372564
rect 228548 372512 228600 372564
rect 3332 346332 3384 346384
rect 220084 346332 220136 346384
rect 362224 325592 362276 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 225696 320084 225748 320136
rect 224960 309068 225012 309120
rect 237196 309068 237248 309120
rect 290556 309068 290608 309120
rect 349436 309068 349488 309120
rect 354864 309068 354916 309120
rect 97264 309000 97316 309052
rect 247684 309000 247736 309052
rect 281448 309000 281500 309052
rect 68284 308932 68336 308984
rect 234620 308932 234672 308984
rect 242256 308932 242308 308984
rect 252192 308932 252244 308984
rect 50344 308864 50396 308916
rect 232872 308864 232924 308916
rect 64144 308796 64196 308848
rect 233792 308796 233844 308848
rect 249340 308796 249392 308848
rect 258264 308796 258316 308848
rect 46204 308728 46256 308780
rect 232044 308728 232096 308780
rect 252008 308728 252060 308780
rect 43444 308660 43496 308712
rect 224960 308660 225012 308712
rect 39304 308592 39356 308644
rect 233516 308592 233568 308644
rect 35900 308524 35952 308576
rect 236552 308660 236604 308712
rect 27620 308456 27672 308508
rect 235264 308524 235316 308576
rect 237104 308524 237156 308576
rect 241796 308592 241848 308644
rect 243544 308592 243596 308644
rect 252652 308660 252704 308712
rect 252744 308660 252796 308712
rect 253572 308660 253624 308712
rect 268384 308728 268436 308780
rect 275652 308728 275704 308780
rect 264244 308660 264296 308712
rect 276940 308660 276992 308712
rect 281356 308932 281408 308984
rect 287704 309000 287756 309052
rect 350816 309000 350868 309052
rect 281172 308864 281224 308916
rect 347320 308932 347372 308984
rect 347964 308864 348016 308916
rect 348608 308796 348660 308848
rect 354220 308796 354272 308848
rect 355600 308796 355652 308848
rect 438124 308864 438176 308916
rect 282736 308728 282788 308780
rect 353208 308728 353260 308780
rect 354680 308728 354732 308780
rect 355416 308728 355468 308780
rect 356244 308728 356296 308780
rect 356520 308728 356572 308780
rect 357440 308728 357492 308780
rect 357900 308728 357952 308780
rect 436836 308796 436888 308848
rect 439504 308728 439556 308780
rect 348792 308660 348844 308712
rect 352932 308660 352984 308712
rect 438032 308660 438084 308712
rect 253756 308592 253808 308644
rect 254400 308592 254452 308644
rect 256056 308592 256108 308644
rect 262864 308592 262916 308644
rect 283932 308592 283984 308644
rect 341064 308592 341116 308644
rect 353576 308592 353628 308644
rect 439412 308592 439464 308644
rect 238944 308524 238996 308576
rect 239588 308524 239640 308576
rect 253572 308524 253624 308576
rect 262220 308524 262272 308576
rect 262496 308524 262548 308576
rect 348148 308524 348200 308576
rect 352288 308524 352340 308576
rect 440424 308524 440476 308576
rect 234712 308456 234764 308508
rect 235908 308456 235960 308508
rect 238116 308456 238168 308508
rect 23480 308388 23532 308440
rect 234988 308388 235040 308440
rect 235540 308388 235592 308440
rect 236092 308388 236144 308440
rect 236644 308388 236696 308440
rect 237564 308388 237616 308440
rect 237932 308388 237984 308440
rect 238760 308388 238812 308440
rect 239128 308388 239180 308440
rect 240324 308388 240376 308440
rect 240968 308388 241020 308440
rect 242900 308388 242952 308440
rect 243452 308388 243504 308440
rect 247684 308388 247736 308440
rect 258908 308388 258960 308440
rect 260196 308388 260248 308440
rect 262588 308388 262640 308440
rect 350172 308456 350224 308508
rect 351644 308456 351696 308508
rect 439596 308456 439648 308508
rect 312084 308388 312136 308440
rect 313004 308388 313056 308440
rect 313372 308388 313424 308440
rect 313648 308388 313700 308440
rect 314660 308388 314712 308440
rect 315672 308388 315724 308440
rect 315764 308388 315816 308440
rect 234804 308320 234856 308372
rect 235448 308320 235500 308372
rect 237472 308320 237524 308372
rect 238392 308320 238444 308372
rect 238852 308320 238904 308372
rect 239404 308320 239456 308372
rect 242992 308320 243044 308372
rect 243728 308320 243780 308372
rect 251916 308320 251968 308372
rect 253756 308320 253808 308372
rect 262312 308320 262364 308372
rect 263048 308320 263100 308372
rect 284208 308320 284260 308372
rect 338396 308320 338448 308372
rect 234436 308252 234488 308304
rect 237656 308252 237708 308304
rect 238300 308252 238352 308304
rect 239220 308252 239272 308304
rect 239680 308252 239732 308304
rect 241612 308252 241664 308304
rect 242624 308252 242676 308304
rect 243084 308252 243136 308304
rect 243820 308252 243872 308304
rect 274824 308252 274876 308304
rect 276296 308252 276348 308304
rect 285496 308252 285548 308304
rect 337292 308252 337344 308304
rect 437480 308388 437532 308440
rect 350724 308320 350776 308372
rect 351828 308320 351880 308372
rect 352012 308320 352064 308372
rect 352564 308320 352616 308372
rect 356060 308320 356112 308372
rect 356612 308320 356664 308372
rect 358912 308320 358964 308372
rect 359740 308320 359792 308372
rect 351000 308252 351052 308304
rect 351276 308252 351328 308304
rect 353668 308252 353720 308304
rect 354312 308252 354364 308304
rect 355140 308252 355192 308304
rect 355968 308252 356020 308304
rect 356152 308252 356204 308304
rect 357256 308252 357308 308304
rect 357808 308252 357860 308304
rect 358360 308252 358412 308304
rect 359004 308252 359056 308304
rect 360108 308252 360160 308304
rect 238760 308184 238812 308236
rect 240048 308184 240100 308236
rect 250996 308184 251048 308236
rect 262496 308184 262548 308236
rect 234252 308116 234304 308168
rect 243176 308116 243228 308168
rect 262864 308116 262916 308168
rect 268384 308116 268436 308168
rect 242532 308048 242584 308100
rect 249800 308048 249852 308100
rect 282644 308048 282696 308100
rect 283564 308048 283616 308100
rect 243728 307980 243780 308032
rect 249156 307980 249208 308032
rect 278780 307980 278832 308032
rect 281264 307980 281316 308032
rect 244924 307912 244976 307964
rect 250444 307912 250496 307964
rect 276664 307912 276716 307964
rect 278872 307912 278924 307964
rect 291016 307912 291068 307964
rect 337568 308184 337620 308236
rect 353392 308184 353444 308236
rect 354036 308184 354088 308236
rect 312176 308116 312228 308168
rect 312360 308116 312412 308168
rect 313556 308116 313608 308168
rect 314292 308116 314344 308168
rect 314752 308116 314804 308168
rect 314936 308116 314988 308168
rect 316316 308116 316368 308168
rect 316868 308116 316920 308168
rect 317604 308116 317656 308168
rect 317788 308116 317840 308168
rect 319076 308116 319128 308168
rect 319720 308116 319772 308168
rect 320272 308116 320324 308168
rect 321008 308116 321060 308168
rect 341064 308116 341116 308168
rect 353852 308116 353904 308168
rect 356336 308116 356388 308168
rect 357072 308116 357124 308168
rect 357624 308116 357676 308168
rect 357992 308116 358044 308168
rect 358820 308116 358872 308168
rect 359280 308116 359332 308168
rect 311900 308048 311952 308100
rect 312544 308048 312596 308100
rect 313280 308048 313332 308100
rect 314476 308048 314528 308100
rect 316224 308048 316276 308100
rect 316960 308048 317012 308100
rect 317512 308048 317564 308100
rect 318432 308048 318484 308100
rect 357532 308048 357584 308100
rect 358452 308048 358504 308100
rect 359188 308048 359240 308100
rect 359464 308048 359516 308100
rect 312176 307980 312228 308032
rect 313188 307980 313240 308032
rect 314752 307980 314804 308032
rect 315580 307980 315632 308032
rect 316132 307980 316184 308032
rect 317328 307980 317380 308032
rect 317420 307980 317472 308032
rect 318616 307980 318668 308032
rect 318800 307980 318852 308032
rect 319260 307980 319312 308032
rect 354772 307980 354824 308032
rect 355784 307980 355836 308032
rect 308036 307912 308088 307964
rect 315764 307912 315816 307964
rect 358820 307912 358872 307964
rect 359648 307912 359700 307964
rect 246488 307844 246540 307896
rect 248972 307844 249024 307896
rect 278136 307844 278188 307896
rect 279792 307844 279844 307896
rect 282828 307844 282880 307896
rect 285128 307844 285180 307896
rect 286048 307844 286100 307896
rect 291844 307844 291896 307896
rect 318800 307844 318852 307896
rect 319904 307844 319956 307896
rect 236644 307776 236696 307828
rect 237104 307776 237156 307828
rect 245016 307776 245068 307828
rect 246856 307776 246908 307828
rect 248512 307776 248564 307828
rect 249064 307776 249116 307828
rect 251364 307776 251416 307828
rect 257344 307776 257396 307828
rect 258080 307776 258132 307828
rect 265624 307776 265676 307828
rect 266728 307776 266780 307828
rect 271144 307776 271196 307828
rect 271972 307776 272024 307828
rect 275376 307776 275428 307828
rect 276756 307776 276808 307828
rect 277124 307776 277176 307828
rect 278044 307776 278096 307828
rect 279516 307776 279568 307828
rect 281080 307776 281132 307828
rect 284116 307776 284168 307828
rect 284944 307776 284996 307828
rect 285036 307776 285088 307828
rect 286324 307776 286376 307828
rect 293224 307776 293276 307828
rect 294696 307776 294748 307828
rect 295156 307776 295208 307828
rect 296444 307776 296496 307828
rect 328644 307708 328696 307760
rect 329380 307708 329432 307760
rect 243268 307640 243320 307692
rect 244188 307640 244240 307692
rect 320364 307640 320416 307692
rect 320548 307640 320600 307692
rect 242164 307572 242216 307624
rect 320548 307504 320600 307556
rect 321468 307504 321520 307556
rect 326712 307232 326764 307284
rect 445024 307232 445076 307284
rect 80060 307164 80112 307216
rect 244832 307164 244884 307216
rect 316500 307164 316552 307216
rect 467104 307164 467156 307216
rect 57980 307096 58032 307148
rect 240692 307096 240744 307148
rect 318248 307096 318300 307148
rect 476764 307096 476816 307148
rect 25504 307028 25556 307080
rect 230112 307028 230164 307080
rect 251180 307028 251232 307080
rect 274824 307028 274876 307080
rect 284300 307028 284352 307080
rect 293224 307028 293276 307080
rect 322112 307028 322164 307080
rect 500224 307028 500276 307080
rect 272156 306960 272208 307012
rect 288900 306960 288952 307012
rect 245844 306824 245896 306876
rect 266360 306756 266412 306808
rect 266636 306756 266688 306808
rect 272064 306756 272116 306808
rect 288992 306756 289044 306808
rect 299480 306688 299532 306740
rect 299940 306688 299992 306740
rect 320180 306688 320232 306740
rect 320732 306688 320784 306740
rect 329840 306688 329892 306740
rect 330208 306688 330260 306740
rect 335820 306688 335872 306740
rect 336096 306688 336148 306740
rect 273444 306620 273496 306672
rect 273628 306620 273680 306672
rect 322940 306620 322992 306672
rect 323492 306620 323544 306672
rect 230940 306552 230992 306604
rect 245844 306552 245896 306604
rect 263876 306552 263928 306604
rect 283012 306552 283064 306604
rect 291660 306552 291712 306604
rect 320180 306552 320232 306604
rect 321100 306552 321152 306604
rect 323216 306552 323268 306604
rect 343640 306552 343692 306604
rect 344008 306552 344060 306604
rect 245936 306484 245988 306536
rect 246396 306484 246448 306536
rect 250076 306484 250128 306536
rect 250536 306484 250588 306536
rect 241520 306416 241572 306468
rect 241796 306416 241848 306468
rect 245752 306416 245804 306468
rect 246304 306416 246356 306468
rect 247316 306416 247368 306468
rect 248144 306416 248196 306468
rect 249892 306416 249944 306468
rect 250260 306416 250312 306468
rect 256976 306416 257028 306468
rect 257160 306416 257212 306468
rect 260840 306416 260892 306468
rect 261300 306416 261352 306468
rect 270684 306416 270736 306468
rect 270960 306416 271012 306468
rect 277584 306416 277636 306468
rect 278228 306416 278280 306468
rect 281540 306416 281592 306468
rect 281908 306416 281960 306468
rect 230940 306348 230992 306400
rect 232044 306348 232096 306400
rect 232964 306348 233016 306400
rect 247408 306348 247460 306400
rect 248052 306348 248104 306400
rect 248512 306348 248564 306400
rect 249248 306348 249300 306400
rect 252652 306348 252704 306400
rect 253296 306348 253348 306400
rect 255412 306348 255464 306400
rect 256516 306348 256568 306400
rect 256884 306348 256936 306400
rect 257712 306348 257764 306400
rect 258264 306348 258316 306400
rect 259000 306348 259052 306400
rect 259644 306348 259696 306400
rect 260012 306348 260064 306400
rect 263876 306348 263928 306400
rect 265348 306348 265400 306400
rect 266084 306348 266136 306400
rect 268108 306348 268160 306400
rect 268568 306348 268620 306400
rect 270500 306348 270552 306400
rect 271604 306348 271656 306400
rect 273352 306348 273404 306400
rect 274364 306348 274416 306400
rect 278964 306348 279016 306400
rect 279332 306348 279384 306400
rect 289820 306416 289872 306468
rect 290648 306416 290700 306468
rect 284392 306348 284444 306400
rect 285220 306348 285272 306400
rect 287244 306348 287296 306400
rect 287796 306348 287848 306400
rect 288624 306348 288676 306400
rect 289728 306348 289780 306400
rect 290096 306348 290148 306400
rect 290832 306348 290884 306400
rect 295616 306484 295668 306536
rect 296352 306484 296404 306536
rect 307760 306484 307812 306536
rect 308404 306484 308456 306536
rect 295432 306416 295484 306468
rect 296076 306416 296128 306468
rect 302240 306416 302292 306468
rect 302516 306416 302568 306468
rect 308036 306416 308088 306468
rect 308496 306416 308548 306468
rect 310520 306416 310572 306468
rect 311256 306416 311308 306468
rect 295708 306348 295760 306400
rect 296260 306348 296312 306400
rect 298284 306348 298336 306400
rect 299296 306348 299348 306400
rect 301044 306348 301096 306400
rect 302148 306348 302200 306400
rect 306656 306348 306708 306400
rect 307116 306348 307168 306400
rect 308128 306348 308180 306400
rect 308864 306348 308916 306400
rect 309324 306348 309376 306400
rect 309968 306348 310020 306400
rect 310704 306348 310756 306400
rect 311440 306348 311492 306400
rect 323124 306348 323176 306400
rect 325792 306484 325844 306536
rect 326896 306484 326948 306536
rect 327356 306484 327408 306536
rect 327908 306484 327960 306536
rect 328368 306484 328420 306536
rect 328920 306484 328972 306536
rect 325700 306416 325752 306468
rect 326436 306416 326488 306468
rect 327080 306416 327132 306468
rect 328184 306416 328236 306468
rect 331312 306416 331364 306468
rect 331680 306416 331732 306468
rect 334072 306416 334124 306468
rect 334348 306416 334400 306468
rect 323308 306348 323360 306400
rect 324044 306348 324096 306400
rect 324320 306348 324372 306400
rect 324596 306348 324648 306400
rect 325884 306348 325936 306400
rect 326252 306348 326304 306400
rect 327264 306348 327316 306400
rect 327724 306348 327776 306400
rect 3332 306280 3384 306332
rect 221464 306280 221516 306332
rect 230664 306280 230716 306332
rect 231584 306280 231636 306332
rect 231952 306280 232004 306332
rect 232504 306280 232556 306332
rect 244464 306280 244516 306332
rect 245476 306280 245528 306332
rect 247040 306280 247092 306332
rect 247592 306280 247644 306332
rect 248604 306280 248656 306332
rect 249616 306280 249668 306332
rect 252836 306280 252888 306332
rect 253020 306280 253072 306332
rect 253940 306280 253992 306332
rect 254216 306280 254268 306332
rect 254308 306280 254360 306332
rect 255044 306280 255096 306332
rect 255320 306280 255372 306332
rect 255964 306280 256016 306332
rect 256792 306280 256844 306332
rect 257252 306280 257304 306332
rect 258172 306280 258224 306332
rect 258724 306280 258776 306332
rect 259460 306280 259512 306332
rect 260104 306280 260156 306332
rect 261024 306280 261076 306332
rect 261760 306280 261812 306332
rect 262496 306280 262548 306332
rect 263508 306280 263560 306332
rect 263600 306280 263652 306332
rect 264428 306280 264480 306332
rect 265256 306280 265308 306332
rect 265532 306280 265584 306332
rect 268016 306280 268068 306332
rect 268292 306280 268344 306332
rect 269212 306280 269264 306332
rect 270408 306280 270460 306332
rect 270592 306280 270644 306332
rect 271512 306280 271564 306332
rect 273536 306280 273588 306332
rect 274548 306280 274600 306332
rect 274916 306280 274968 306332
rect 275836 306280 275888 306332
rect 277768 306280 277820 306332
rect 278320 306280 278372 306332
rect 278872 306280 278924 306332
rect 279976 306280 280028 306332
rect 283012 306280 283064 306332
rect 283656 306280 283708 306332
rect 284300 306280 284352 306332
rect 284760 306280 284812 306332
rect 287152 306280 287204 306332
rect 287428 306280 287480 306332
rect 288440 306280 288492 306332
rect 288808 306280 288860 306332
rect 290004 306280 290056 306332
rect 290924 306280 290976 306332
rect 291660 306280 291712 306332
rect 292672 306280 292724 306332
rect 293684 306280 293736 306332
rect 293960 306280 294012 306332
rect 294604 306280 294656 306332
rect 295524 306280 295576 306332
rect 295892 306280 295944 306332
rect 298192 306280 298244 306332
rect 298652 306280 298704 306332
rect 299848 306280 299900 306332
rect 300400 306280 300452 306332
rect 300952 306280 301004 306332
rect 301504 306280 301556 306332
rect 301596 306280 301648 306332
rect 331588 306348 331640 306400
rect 332508 306348 332560 306400
rect 333980 306348 334032 306400
rect 334900 306348 334952 306400
rect 338304 306348 338356 306400
rect 339132 306348 339184 306400
rect 341156 306348 341208 306400
rect 341616 306348 341668 306400
rect 345204 306348 345256 306400
rect 345756 306348 345808 306400
rect 230756 306212 230808 306264
rect 231032 306212 231084 306264
rect 246120 306212 246172 306264
rect 246764 306212 246816 306264
rect 247224 306212 247276 306264
rect 247868 306212 247920 306264
rect 259552 306212 259604 306264
rect 259920 306212 259972 306264
rect 263784 306212 263836 306264
rect 264336 306212 264388 306264
rect 264980 306212 265032 306264
rect 265900 306212 265952 306264
rect 266820 306212 266872 306264
rect 267372 306212 267424 306264
rect 267740 306212 267792 306264
rect 268476 306212 268528 306264
rect 270776 306212 270828 306264
rect 271052 306212 271104 306264
rect 272156 306212 272208 306264
rect 272800 306212 272852 306264
rect 273628 306212 273680 306264
rect 273904 306212 273956 306264
rect 275928 306212 275980 306264
rect 255504 306144 255556 306196
rect 255872 306144 255924 306196
rect 260932 306144 260984 306196
rect 261392 306144 261444 306196
rect 263968 306144 264020 306196
rect 264796 306144 264848 306196
rect 266544 306144 266596 306196
rect 267464 306144 267516 306196
rect 267832 306144 267884 306196
rect 268936 306144 268988 306196
rect 270868 306144 270920 306196
rect 271328 306144 271380 306196
rect 273260 306144 273312 306196
rect 273812 306144 273864 306196
rect 274732 306144 274784 306196
rect 275192 306144 275244 306196
rect 276296 306144 276348 306196
rect 277032 306144 277084 306196
rect 277676 306144 277728 306196
rect 278688 306144 278740 306196
rect 280252 306144 280304 306196
rect 280712 306144 280764 306196
rect 281632 306144 281684 306196
rect 282184 306144 282236 306196
rect 283104 306212 283156 306264
rect 283288 306212 283340 306264
rect 283748 306212 283800 306264
rect 285772 306212 285824 306264
rect 286508 306212 286560 306264
rect 288900 306212 288952 306264
rect 289544 306212 289596 306264
rect 291568 306212 291620 306264
rect 292120 306212 292172 306264
rect 292396 306212 292448 306264
rect 331128 306212 331180 306264
rect 331404 306212 331456 306264
rect 331956 306212 332008 306264
rect 332600 306212 332652 306264
rect 332968 306212 333020 306264
rect 334164 306212 334216 306264
rect 334716 306212 334768 306264
rect 335360 306212 335412 306264
rect 335728 306212 335780 306264
rect 339684 306212 339736 306264
rect 340328 306212 340380 306264
rect 341064 306280 341116 306332
rect 341432 306280 341484 306332
rect 342720 306280 342772 306332
rect 344100 306280 344152 306332
rect 344928 306280 344980 306332
rect 345296 306280 345348 306332
rect 345480 306280 345532 306332
rect 342536 306212 342588 306264
rect 343364 306212 343416 306264
rect 345020 306212 345072 306264
rect 345848 306212 345900 306264
rect 347964 306212 348016 306264
rect 348240 306212 348292 306264
rect 349344 306212 349396 306264
rect 349896 306212 349948 306264
rect 341892 306144 341944 306196
rect 345296 306144 345348 306196
rect 346216 306144 346268 306196
rect 349252 306144 349304 306196
rect 349620 306144 349672 306196
rect 230756 306076 230808 306128
rect 231768 306076 231820 306128
rect 255688 306076 255740 306128
rect 256332 306076 256384 306128
rect 257068 306076 257120 306128
rect 257620 306076 257672 306128
rect 259552 306076 259604 306128
rect 260656 306076 260708 306128
rect 279056 306076 279108 306128
rect 279332 306076 279384 306128
rect 281724 306076 281776 306128
rect 282368 306076 282420 306128
rect 254124 306008 254176 306060
rect 255228 306008 255280 306060
rect 259736 306008 259788 306060
rect 260472 306008 260524 306060
rect 260932 306008 260984 306060
rect 261944 306008 261996 306060
rect 273260 306008 273312 306060
rect 273996 306008 274048 306060
rect 274732 306008 274784 306060
rect 275284 306008 275336 306060
rect 277308 306008 277360 306060
rect 344468 306076 344520 306128
rect 349436 306076 349488 306128
rect 350356 306076 350408 306128
rect 287428 306008 287480 306060
rect 288256 306008 288308 306060
rect 288440 306008 288492 306060
rect 289176 306008 289228 306060
rect 291476 306008 291528 306060
rect 291936 306008 291988 306060
rect 292028 306008 292080 306060
rect 351184 306008 351236 306060
rect 281080 305940 281132 305992
rect 350632 305940 350684 305992
rect 282368 305872 282420 305924
rect 352012 305872 352064 305924
rect 282276 305804 282328 305856
rect 353760 305804 353812 305856
rect 282184 305736 282236 305788
rect 353392 305736 353444 305788
rect 281172 305668 281224 305720
rect 353668 305668 353720 305720
rect 82176 305600 82228 305652
rect 241980 305600 242032 305652
rect 278688 305600 278740 305652
rect 358820 305600 358872 305652
rect 291292 305532 291344 305584
rect 292212 305532 292264 305584
rect 292856 305532 292908 305584
rect 293316 305532 293368 305584
rect 294236 305532 294288 305584
rect 294972 305532 295024 305584
rect 298376 305532 298428 305584
rect 299112 305532 299164 305584
rect 300124 305532 300176 305584
rect 284024 305464 284076 305516
rect 292028 305464 292080 305516
rect 299572 305464 299624 305516
rect 300584 305464 300636 305516
rect 296628 305328 296680 305380
rect 296812 305328 296864 305380
rect 299204 305328 299256 305380
rect 331864 305464 331916 305516
rect 294972 305260 295024 305312
rect 300124 305260 300176 305312
rect 285680 305192 285732 305244
rect 286692 305192 286744 305244
rect 296628 305192 296680 305244
rect 301596 305192 301648 305244
rect 283932 305124 283984 305176
rect 284208 305124 284260 305176
rect 299480 305124 299532 305176
rect 300216 305124 300268 305176
rect 299296 305056 299348 305108
rect 302332 305328 302384 305380
rect 302792 305328 302844 305380
rect 306380 305328 306432 305380
rect 306840 305328 306892 305380
rect 307944 305328 307996 305380
rect 309048 305328 309100 305380
rect 310612 305328 310664 305380
rect 310888 305328 310940 305380
rect 321652 305328 321704 305380
rect 322296 305328 322348 305380
rect 323124 305328 323176 305380
rect 323860 305328 323912 305380
rect 324504 305328 324556 305380
rect 325148 305328 325200 305380
rect 328644 305328 328696 305380
rect 329472 305328 329524 305380
rect 330024 305328 330076 305380
rect 330576 305328 330628 305380
rect 331220 305328 331272 305380
rect 331772 305328 331824 305380
rect 302608 305260 302660 305312
rect 303436 305260 303488 305312
rect 306564 305260 306616 305312
rect 307576 305260 307628 305312
rect 324320 305260 324372 305312
rect 325424 305260 325476 305312
rect 328552 305260 328604 305312
rect 329564 305260 329616 305312
rect 330116 305260 330168 305312
rect 330852 305260 330904 305312
rect 302424 305192 302476 305244
rect 303068 305192 303120 305244
rect 306380 305192 306432 305244
rect 307208 305192 307260 305244
rect 310612 305192 310664 305244
rect 311532 305192 311584 305244
rect 321560 305192 321612 305244
rect 322388 305192 322440 305244
rect 329932 305192 329984 305244
rect 330760 305192 330812 305244
rect 332968 305532 333020 305584
rect 333704 305532 333756 305584
rect 334256 305532 334308 305584
rect 334992 305532 335044 305584
rect 335544 305532 335596 305584
rect 336648 305532 336700 305584
rect 339592 305532 339644 305584
rect 340420 305532 340472 305584
rect 332784 305464 332836 305516
rect 333244 305464 333296 305516
rect 335360 305464 335412 305516
rect 336280 305464 336332 305516
rect 332692 305396 332744 305448
rect 333612 305396 333664 305448
rect 332232 305328 332284 305380
rect 338580 305328 338632 305380
rect 337936 305260 337988 305312
rect 339960 305124 340012 305176
rect 305092 305056 305144 305108
rect 305828 305056 305880 305108
rect 331864 305056 331916 305108
rect 340788 305056 340840 305108
rect 269304 304988 269356 305040
rect 269672 304988 269724 305040
rect 331220 304988 331272 305040
rect 332324 304988 332376 305040
rect 304540 304512 304592 304564
rect 88984 304308 89036 304360
rect 242992 304308 243044 304360
rect 303620 304308 303672 304360
rect 304080 304308 304132 304360
rect 7564 304240 7616 304292
rect 230480 304240 230532 304292
rect 251456 304240 251508 304292
rect 251732 304240 251784 304292
rect 271972 304240 272024 304292
rect 272248 304240 272300 304292
rect 287060 304240 287112 304292
rect 287888 304240 287940 304292
rect 303620 304172 303672 304224
rect 315396 304444 315448 304496
rect 458824 304444 458876 304496
rect 319260 304376 319312 304428
rect 478144 304376 478196 304428
rect 324688 304308 324740 304360
rect 514024 304308 514076 304360
rect 305184 304240 305236 304292
rect 305460 304240 305512 304292
rect 309232 304240 309284 304292
rect 309600 304240 309652 304292
rect 310796 304240 310848 304292
rect 311072 304240 311124 304292
rect 334532 304240 334584 304292
rect 566464 304240 566516 304292
rect 250168 303696 250220 303748
rect 251088 303696 251140 303748
rect 280988 303560 281040 303612
rect 354680 303560 354732 303612
rect 268476 303492 268528 303544
rect 344744 303492 344796 303544
rect 268568 303424 268620 303476
rect 343824 303424 343876 303476
rect 279608 303356 279660 303408
rect 356060 303356 356112 303408
rect 279516 303288 279568 303340
rect 356152 303288 356204 303340
rect 268384 303220 268436 303272
rect 345572 303220 345624 303272
rect 276940 303152 276992 303204
rect 357532 303152 357584 303204
rect 85580 303016 85632 303068
rect 245660 303084 245712 303136
rect 251364 303084 251416 303136
rect 252284 303084 252336 303136
rect 276848 303084 276900 303136
rect 357440 303084 357492 303136
rect 244372 303016 244424 303068
rect 276756 303016 276808 303068
rect 359372 303016 359424 303068
rect 77300 302948 77352 303000
rect 274088 302948 274140 303000
rect 358912 302948 358964 303000
rect 8944 302880 8996 302932
rect 231400 302880 231452 302932
rect 244372 302880 244424 302932
rect 245108 302880 245160 302932
rect 273904 302880 273956 302932
rect 360568 302880 360620 302932
rect 271236 302812 271288 302864
rect 342996 302812 343048 302864
rect 271420 302744 271472 302796
rect 342076 302744 342128 302796
rect 251272 302676 251324 302728
rect 251824 302676 251876 302728
rect 271328 302676 271380 302728
rect 340972 302676 341024 302728
rect 269304 302336 269356 302388
rect 270224 302336 270276 302388
rect 343824 302200 343876 302252
rect 344284 302200 344336 302252
rect 292764 301996 292816 302048
rect 293040 301996 293092 302048
rect 95884 301588 95936 301640
rect 247592 301588 247644 301640
rect 316592 301588 316644 301640
rect 468484 301588 468536 301640
rect 93860 301520 93912 301572
rect 247132 301520 247184 301572
rect 320640 301520 320692 301572
rect 494060 301520 494112 301572
rect 48964 301452 49016 301504
rect 239128 301452 239180 301504
rect 329380 301452 329432 301504
rect 534724 301452 534776 301504
rect 288716 301248 288768 301300
rect 289084 301248 289136 301300
rect 290924 300772 290976 300824
rect 342444 300772 342496 300824
rect 289544 300704 289596 300756
rect 341064 300704 341116 300756
rect 286784 300636 286836 300688
rect 338304 300636 338356 300688
rect 289452 300568 289504 300620
rect 344192 300568 344244 300620
rect 283932 300500 283984 300552
rect 338212 300500 338264 300552
rect 286600 300432 286652 300484
rect 343180 300432 343232 300484
rect 286876 300364 286928 300416
rect 346584 300364 346636 300416
rect 285312 300296 285364 300348
rect 345020 300296 345072 300348
rect 282736 300228 282788 300280
rect 352472 300228 352524 300280
rect 53104 300160 53156 300212
rect 238852 300160 238904 300212
rect 278412 300160 278464 300212
rect 349528 300160 349580 300212
rect 40040 300092 40092 300144
rect 237380 300092 237432 300144
rect 278504 300092 278556 300144
rect 349344 300092 349396 300144
rect 288256 300024 288308 300076
rect 339684 300024 339736 300076
rect 285128 299956 285180 300008
rect 337108 299956 337160 300008
rect 292212 299888 292264 299940
rect 340144 299888 340196 299940
rect 322756 298868 322808 298920
rect 502984 298868 503036 298920
rect 53840 298800 53892 298852
rect 238760 298800 238812 298852
rect 331772 298800 331824 298852
rect 549904 298800 549956 298852
rect 10324 298732 10376 298784
rect 231032 298732 231084 298784
rect 239404 298732 239456 298784
rect 251548 298732 251600 298784
rect 334348 298732 334400 298784
rect 563704 298732 563756 298784
rect 298008 297984 298060 298036
rect 356336 297984 356388 298036
rect 297916 297916 297968 297968
rect 356244 297916 356296 297968
rect 277216 297848 277268 297900
rect 338396 297848 338448 297900
rect 278320 297780 278372 297832
rect 341524 297780 341576 297832
rect 284852 297712 284904 297764
rect 360292 297712 360344 297764
rect 279976 297644 280028 297696
rect 359096 297644 359148 297696
rect 317972 297576 318024 297628
rect 462964 297576 463016 297628
rect 316224 297508 316276 297560
rect 473452 297508 473504 297560
rect 60740 297440 60792 297492
rect 241336 297440 241388 297492
rect 285864 297440 285916 297492
rect 323400 297440 323452 297492
rect 507860 297440 507912 297492
rect 62120 297372 62172 297424
rect 241796 297372 241848 297424
rect 333152 297372 333204 297424
rect 561680 297372 561732 297424
rect 285956 297236 286008 297288
rect 323308 296080 323360 296132
rect 512000 296080 512052 296132
rect 71044 296012 71096 296064
rect 243452 296012 243504 296064
rect 330116 296012 330168 296064
rect 548524 296012 548576 296064
rect 66904 295944 66956 295996
rect 241704 295944 241756 295996
rect 334256 295944 334308 295996
rect 570604 295944 570656 295996
rect 321836 294720 321888 294772
rect 493324 294720 493376 294772
rect 325976 294652 326028 294704
rect 521660 294652 521712 294704
rect 69020 294584 69072 294636
rect 241612 294584 241664 294636
rect 327540 294584 327592 294636
rect 529940 294584 529992 294636
rect 3332 293904 3384 293956
rect 228456 293904 228508 293956
rect 325884 293360 325936 293412
rect 522304 293360 522356 293412
rect 327448 293292 327500 293344
rect 527824 293292 527876 293344
rect 86960 293224 87012 293276
rect 246028 293224 246080 293276
rect 335820 293224 335872 293276
rect 578240 293224 578292 293276
rect 71780 291864 71832 291916
rect 243176 291864 243228 291916
rect 328828 291864 328880 291916
rect 536104 291864 536156 291916
rect 30380 291796 30432 291848
rect 234988 291796 235040 291848
rect 328920 291796 328972 291848
rect 538864 291796 538916 291848
rect 75920 290504 75972 290556
rect 243084 290504 243136 290556
rect 330024 290504 330076 290556
rect 547972 290504 548024 290556
rect 41420 290436 41472 290488
rect 237748 290436 237800 290488
rect 243636 290436 243688 290488
rect 252928 290436 252980 290488
rect 334164 290436 334216 290488
rect 567844 290436 567896 290488
rect 310980 289212 311032 289264
rect 440240 289212 440292 289264
rect 56600 289144 56652 289196
rect 240416 289144 240468 289196
rect 331680 289144 331732 289196
rect 552664 289144 552716 289196
rect 13084 289076 13136 289128
rect 232136 289076 232188 289128
rect 335728 289076 335780 289128
rect 571984 289076 572036 289128
rect 313924 287716 313976 287768
rect 449900 287716 449952 287768
rect 9680 287648 9732 287700
rect 230756 287648 230808 287700
rect 331588 287648 331640 287700
rect 557540 287648 557592 287700
rect 312268 286492 312320 286544
rect 448520 286492 448572 286544
rect 318064 286424 318116 286476
rect 456892 286424 456944 286476
rect 89720 286356 89772 286408
rect 245936 286356 245988 286408
rect 313648 286356 313700 286408
rect 456800 286356 456852 286408
rect 46296 286288 46348 286340
rect 237656 286288 237708 286340
rect 332968 286288 333020 286340
rect 563796 286288 563848 286340
rect 310796 285064 310848 285116
rect 440332 285064 440384 285116
rect 324688 284996 324740 285048
rect 516140 284996 516192 285048
rect 34520 284928 34572 284980
rect 236276 284928 236328 284980
rect 328736 284928 328788 284980
rect 535460 284928 535512 284980
rect 310704 283704 310756 283756
rect 443000 283704 443052 283756
rect 60832 283636 60884 283688
rect 240324 283636 240376 283688
rect 313556 283636 313608 283688
rect 454684 283636 454736 283688
rect 16580 283568 16632 283620
rect 232044 283568 232096 283620
rect 332876 283568 332928 283620
rect 554044 283568 554096 283620
rect 313464 282276 313516 282328
rect 450544 282276 450596 282328
rect 70400 282208 70452 282260
rect 233884 282208 233936 282260
rect 317696 282208 317748 282260
rect 475384 282208 475436 282260
rect 20720 282140 20772 282192
rect 233424 282140 233476 282192
rect 335636 282140 335688 282192
rect 574744 282140 574796 282192
rect 312176 280916 312228 280968
rect 452660 280916 452712 280968
rect 93124 280848 93176 280900
rect 245844 280848 245896 280900
rect 319076 280848 319128 280900
rect 488540 280848 488592 280900
rect 26240 280780 26292 280832
rect 234896 280780 234948 280832
rect 334072 280780 334124 280832
rect 567200 280780 567252 280832
rect 314936 279556 314988 279608
rect 460940 279556 460992 279608
rect 88340 279488 88392 279540
rect 245752 279488 245804 279540
rect 315028 279488 315080 279540
rect 463700 279488 463752 279540
rect 29000 279420 29052 279472
rect 234804 279420 234856 279472
rect 320456 279420 320508 279472
rect 491300 279420 491352 279472
rect 318984 278060 319036 278112
rect 485780 278060 485832 278112
rect 35164 277992 35216 278044
rect 236184 277992 236236 278044
rect 323216 277992 323268 278044
rect 506480 277992 506532 278044
rect 317604 276700 317656 276752
rect 477500 276700 477552 276752
rect 35992 276632 36044 276684
rect 236092 276632 236144 276684
rect 324596 276632 324648 276684
rect 509884 276632 509936 276684
rect 320364 275340 320416 275392
rect 492680 275340 492732 275392
rect 44180 275272 44232 275324
rect 237564 275272 237616 275324
rect 325792 275272 325844 275324
rect 526536 275272 526588 275324
rect 310612 274048 310664 274100
rect 444380 274048 444432 274100
rect 321744 273980 321796 274032
rect 499580 273980 499632 274032
rect 14464 273912 14516 273964
rect 230664 273912 230716 273964
rect 327356 273912 327408 273964
rect 531320 273912 531372 273964
rect 367744 273164 367796 273216
rect 579896 273164 579948 273216
rect 48320 272484 48372 272536
rect 239036 272484 239088 272536
rect 324504 272484 324556 272536
rect 517520 272484 517572 272536
rect 312084 271260 312136 271312
rect 446404 271260 446456 271312
rect 323124 271192 323176 271244
rect 510620 271192 510672 271244
rect 52460 271124 52512 271176
rect 238944 271124 238996 271176
rect 328644 271124 328696 271176
rect 540244 271124 540296 271176
rect 313372 269900 313424 269952
rect 453304 269900 453356 269952
rect 325700 269832 325752 269884
rect 524420 269832 524472 269884
rect 57244 269764 57296 269816
rect 240232 269764 240284 269816
rect 329932 269764 329984 269816
rect 543004 269764 543056 269816
rect 314844 268472 314896 268524
rect 460204 268472 460256 268524
rect 327264 268404 327316 268456
rect 531412 268404 531464 268456
rect 59360 268336 59412 268388
rect 240508 268336 240560 268388
rect 331496 268336 331548 268388
rect 552020 268336 552072 268388
rect 2964 267656 3016 267708
rect 224224 267656 224276 267708
rect 314752 267180 314804 267232
rect 464344 267180 464396 267232
rect 328552 267112 328604 267164
rect 542360 267112 542412 267164
rect 331404 267044 331456 267096
rect 556160 267044 556212 267096
rect 99288 266976 99340 267028
rect 335544 266976 335596 267028
rect 238208 265820 238260 265872
rect 351000 265820 351052 265872
rect 317512 265752 317564 265804
rect 481640 265752 481692 265804
rect 329840 265684 329892 265736
rect 546500 265684 546552 265736
rect 66260 265616 66312 265668
rect 241888 265616 241940 265668
rect 332784 265616 332836 265668
rect 560944 265616 560996 265668
rect 317420 264256 317472 264308
rect 481732 264256 481784 264308
rect 75184 264188 75236 264240
rect 243360 264188 243412 264240
rect 318892 264188 318944 264240
rect 484400 264188 484452 264240
rect 77392 262896 77444 262948
rect 243268 262896 243320 262948
rect 318800 262896 318852 262948
rect 490012 262896 490064 262948
rect 4160 262828 4212 262880
rect 230940 262828 230992 262880
rect 320272 262828 320324 262880
rect 495440 262828 495492 262880
rect 84200 261536 84252 261588
rect 244464 261536 244516 261588
rect 320180 261536 320232 261588
rect 496084 261536 496136 261588
rect 31760 261468 31812 261520
rect 234712 261468 234764 261520
rect 321652 261468 321704 261520
rect 502340 261468 502392 261520
rect 311992 260244 312044 260296
rect 445760 260244 445812 260296
rect 91100 260176 91152 260228
rect 246120 260176 246172 260228
rect 364984 260176 365036 260228
rect 580448 260176 580500 260228
rect 13820 260108 13872 260160
rect 231952 260108 232004 260160
rect 332692 260108 332744 260160
rect 564532 260108 564584 260160
rect 314660 258816 314712 258868
rect 466460 258816 466512 258868
rect 319444 258748 319496 258800
rect 471980 258748 472032 258800
rect 63500 258680 63552 258732
rect 236644 258680 236696 258732
rect 363604 258680 363656 258732
rect 580356 258680 580408 258732
rect 373264 257320 373316 257372
rect 581092 257320 581144 257372
rect 3148 255212 3200 255264
rect 225604 255212 225656 255264
rect 299388 254736 299440 254788
rect 336924 254736 336976 254788
rect 297548 254668 297600 254720
rect 342628 254668 342680 254720
rect 316040 254600 316092 254652
rect 467840 254600 467892 254652
rect 316132 254532 316184 254584
rect 474740 254532 474792 254584
rect 297640 253444 297692 253496
rect 339592 253444 339644 253496
rect 297180 253376 297232 253428
rect 343824 253376 343876 253428
rect 309508 253308 309560 253360
rect 436744 253308 436796 253360
rect 333980 253240 334032 253292
rect 571340 253240 571392 253292
rect 27712 253172 27764 253224
rect 235080 253172 235132 253224
rect 335452 253172 335504 253224
rect 574100 253172 574152 253224
rect 297456 252016 297508 252068
rect 341156 252016 341208 252068
rect 321560 251948 321612 252000
rect 503720 251948 503772 252000
rect 323032 251880 323084 251932
rect 506572 251880 506624 251932
rect 12440 251812 12492 251864
rect 232228 251812 232280 251864
rect 332600 251812 332652 251864
rect 560300 251812 560352 251864
rect 238392 250588 238444 250640
rect 355140 250588 355192 250640
rect 310520 250520 310572 250572
rect 441620 250520 441672 250572
rect 39396 250452 39448 250504
rect 236368 250452 236420 250504
rect 324412 250452 324464 250504
rect 514116 250452 514168 250504
rect 313280 249092 313332 249144
rect 459560 249092 459612 249144
rect 4804 249024 4856 249076
rect 229192 249024 229244 249076
rect 331312 249024 331364 249076
rect 553400 249024 553452 249076
rect 289360 248344 289412 248396
rect 303804 248344 303856 248396
rect 298652 248276 298704 248328
rect 345480 248276 345532 248328
rect 296536 248208 296588 248260
rect 344100 248208 344152 248260
rect 292304 248140 292356 248192
rect 345204 248140 345256 248192
rect 359004 248140 359056 248192
rect 438216 248140 438268 248192
rect 293684 248072 293736 248124
rect 350908 248072 350960 248124
rect 356428 248072 356480 248124
rect 436928 248072 436980 248124
rect 290740 248004 290792 248056
rect 347964 248004 348016 248056
rect 357716 248004 357768 248056
rect 440516 248004 440568 248056
rect 288164 247936 288216 247988
rect 348332 247936 348384 247988
rect 359280 247936 359332 247988
rect 441712 247936 441764 247988
rect 285588 247868 285640 247920
rect 304080 247868 304132 247920
rect 308220 247868 308272 247920
rect 437572 247868 437624 247920
rect 287980 247800 288032 247852
rect 305368 247800 305420 247852
rect 308128 247800 308180 247852
rect 438860 247800 438912 247852
rect 287888 247732 287940 247784
rect 303988 247732 304040 247784
rect 322940 247732 322992 247784
rect 509240 247732 509292 247784
rect 3700 247664 3752 247716
rect 228364 247664 228416 247716
rect 289176 247664 289228 247716
rect 305276 247664 305328 247716
rect 327172 247664 327224 247716
rect 528560 247664 528612 247716
rect 284760 247596 284812 247648
rect 305184 247596 305236 247648
rect 286968 247528 287020 247580
rect 303896 247528 303948 247580
rect 286692 247460 286744 247512
rect 305460 247460 305512 247512
rect 300768 246644 300820 246696
rect 346492 246644 346544 246696
rect 297272 246576 297324 246628
rect 349436 246576 349488 246628
rect 289636 246508 289688 246560
rect 349252 246508 349304 246560
rect 311900 246440 311952 246492
rect 448612 246440 448664 246492
rect 327080 246372 327132 246424
rect 534080 246372 534132 246424
rect 7656 246304 7708 246356
rect 230848 246304 230900 246356
rect 331220 246304 331272 246356
rect 556252 246304 556304 246356
rect 292120 245556 292172 245608
rect 302332 245556 302384 245608
rect 357624 245556 357676 245608
rect 440608 245556 440660 245608
rect 307944 245488 307996 245540
rect 437664 245488 437716 245540
rect 291752 245420 291804 245472
rect 306656 245420 306708 245472
rect 309232 245420 309284 245472
rect 439044 245420 439096 245472
rect 293408 245352 293460 245404
rect 305000 245352 305052 245404
rect 307852 245352 307904 245404
rect 437848 245352 437900 245404
rect 295064 245284 295116 245336
rect 305092 245284 305144 245336
rect 308036 245284 308088 245336
rect 439136 245284 439188 245336
rect 293776 245216 293828 245268
rect 302424 245216 302476 245268
rect 306748 245216 306800 245268
rect 437940 245216 437992 245268
rect 295248 245148 295300 245200
rect 299572 245148 299624 245200
rect 306472 245148 306524 245200
rect 437756 245148 437808 245200
rect 288348 245080 288400 245132
rect 296904 245080 296956 245132
rect 307760 245080 307812 245132
rect 439320 245080 439372 245132
rect 295156 245012 295208 245064
rect 303712 245012 303764 245064
rect 306564 245012 306616 245064
rect 438952 245012 439004 245064
rect 22100 244944 22152 244996
rect 233516 244944 233568 244996
rect 291108 244944 291160 244996
rect 299756 244944 299808 244996
rect 306380 244944 306432 244996
rect 439228 244944 439280 244996
rect 17960 244876 18012 244928
rect 233332 244876 233384 244928
rect 291016 244876 291068 244928
rect 300860 244876 300912 244928
rect 324320 244876 324372 244928
rect 520280 244876 520332 244928
rect 298928 244808 298980 244860
rect 339868 244808 339920 244860
rect 359188 244808 359240 244860
rect 441804 244808 441856 244860
rect 297732 244740 297784 244792
rect 335360 244740 335412 244792
rect 356520 244740 356572 244792
rect 438308 244740 438360 244792
rect 290648 244672 290700 244724
rect 306840 244672 306892 244724
rect 360384 244672 360436 244724
rect 439688 244672 439740 244724
rect 298836 244604 298888 244656
rect 342536 244604 342588 244656
rect 97908 244332 97960 244384
rect 297180 244332 297232 244384
rect 297364 244332 297416 244384
rect 297824 244332 297876 244384
rect 303620 244332 303672 244384
rect 3608 244264 3660 244316
rect 299112 244264 299164 244316
rect 295064 243924 295116 243976
rect 300768 243924 300820 243976
rect 299020 243856 299072 243908
rect 344008 243856 344060 243908
rect 299112 243788 299164 243840
rect 345388 243788 345440 243840
rect 293776 243720 293828 243772
rect 348056 243720 348108 243772
rect 297824 243652 297876 243704
rect 357900 243652 357952 243704
rect 285220 243584 285272 243636
rect 346860 243584 346912 243636
rect 286692 243516 286744 243568
rect 357808 243516 357860 243568
rect 97816 243380 97868 243432
rect 298652 243380 298704 243432
rect 3240 241408 3292 241460
rect 98644 241408 98696 241460
rect 3148 215228 3200 215280
rect 93216 215228 93268 215280
rect 293684 197276 293736 197328
rect 297180 197276 297232 197328
rect 297272 196392 297324 196444
rect 298560 196392 298612 196444
rect 3148 188980 3200 189032
rect 95976 188980 96028 189032
rect 285128 171028 285180 171080
rect 298008 171028 298060 171080
rect 238300 170348 238352 170400
rect 285128 170348 285180 170400
rect 295064 169260 295116 169312
rect 297272 169260 297324 169312
rect 238484 167628 238536 167680
rect 297732 167628 297784 167680
rect 3516 164160 3568 164212
rect 86224 164160 86276 164212
rect 261208 162120 261260 162172
rect 277032 162120 277084 162172
rect 97908 159876 97960 159928
rect 298836 159876 298888 159928
rect 97540 159808 97592 159860
rect 297640 159808 297692 159860
rect 97724 159740 97776 159792
rect 297456 159740 297508 159792
rect 97816 159672 97868 159724
rect 297364 159672 297416 159724
rect 97356 159604 97408 159656
rect 238484 159604 238536 159656
rect 298928 159604 298980 159656
rect 299296 159604 299348 159656
rect 97448 159536 97500 159588
rect 238300 159536 238352 159588
rect 286324 159536 286376 159588
rect 299480 159536 299532 159588
rect 287520 159468 287572 159520
rect 313280 159468 313332 159520
rect 288992 159400 289044 159452
rect 320180 159400 320232 159452
rect 234620 159332 234672 159384
rect 273812 159332 273864 159384
rect 296536 159332 296588 159384
rect 345940 159332 345992 159384
rect 297272 159264 297324 159316
rect 351000 159264 351052 159316
rect 292304 159196 292356 159248
rect 348240 159196 348292 159248
rect 163504 159128 163556 159180
rect 290464 159128 290516 159180
rect 293776 159128 293828 159180
rect 356060 159128 356112 159180
rect 203432 159060 203484 159112
rect 274088 159060 274140 159112
rect 290740 159060 290792 159112
rect 358452 159060 358504 159112
rect 165988 158992 166040 159044
rect 238116 158992 238168 159044
rect 298560 158992 298612 159044
rect 365904 158992 365956 159044
rect 160928 158924 160980 158976
rect 251916 158924 251968 158976
rect 285220 158924 285272 158976
rect 353576 158924 353628 158976
rect 158536 158856 158588 158908
rect 250444 158856 250496 158908
rect 297180 158856 297232 158908
rect 368204 158856 368256 158908
rect 168288 158788 168340 158840
rect 287704 158788 287756 158840
rect 288164 158788 288216 158840
rect 360844 158788 360896 158840
rect 289636 158720 289688 158772
rect 363420 158720 363472 158772
rect 393504 158720 393556 158772
rect 440516 158720 440568 158772
rect 119712 158652 119764 158704
rect 286140 158652 286192 158704
rect 290924 158652 290976 158704
rect 338396 158652 338448 158704
rect 371056 158652 371108 158704
rect 439596 158652 439648 158704
rect 131304 158584 131356 158636
rect 276020 158584 276072 158636
rect 280896 158584 280948 158636
rect 281172 158584 281224 158636
rect 294972 158584 295024 158636
rect 328276 158584 328328 158636
rect 373448 158584 373500 158636
rect 440424 158584 440476 158636
rect 130200 158516 130252 158568
rect 299020 158516 299072 158568
rect 299296 158516 299348 158568
rect 299572 158516 299624 158568
rect 332232 158516 332284 158568
rect 376024 158516 376076 158568
rect 438032 158516 438084 158568
rect 121184 158380 121236 158432
rect 288256 158448 288308 158500
rect 320548 158448 320600 158500
rect 378600 158448 378652 158500
rect 439412 158448 439464 158500
rect 289452 158380 289504 158432
rect 343548 158380 343600 158432
rect 380992 158380 381044 158432
rect 436836 158380 436888 158432
rect 286600 158312 286652 158364
rect 340972 158312 341024 158364
rect 383568 158312 383620 158364
rect 438124 158312 438176 158364
rect 122104 158244 122156 158296
rect 289636 158244 289688 158296
rect 292212 158244 292264 158296
rect 333612 158244 333664 158296
rect 385960 158244 386012 158296
rect 439504 158244 439556 158296
rect 295892 158176 295944 158228
rect 296628 158176 296680 158228
rect 328644 158176 328696 158228
rect 388536 158176 388588 158228
rect 436928 158176 436980 158228
rect 133512 158108 133564 158160
rect 284576 158108 284628 158160
rect 286140 158108 286192 158160
rect 286784 158108 286836 158160
rect 319444 158108 319496 158160
rect 391480 158108 391532 158160
rect 438308 158108 438360 158160
rect 127624 158040 127676 158092
rect 274640 158040 274692 158092
rect 278320 158040 278372 158092
rect 336004 158040 336056 158092
rect 395896 158040 395948 158092
rect 440608 158040 440660 158092
rect 277216 157972 277268 158024
rect 330484 157972 330536 158024
rect 398472 157972 398524 158024
rect 441712 157972 441764 158024
rect 159824 157904 159876 157956
rect 284668 157904 284720 157956
rect 299296 157904 299348 157956
rect 329932 157904 329984 157956
rect 401416 157904 401468 157956
rect 441804 157904 441856 157956
rect 158168 157836 158220 157888
rect 278688 157836 278740 157888
rect 191104 157768 191156 157820
rect 279608 157768 279660 157820
rect 128728 157700 128780 157752
rect 295892 157700 295944 157752
rect 97632 157632 97684 157684
rect 297548 157632 297600 157684
rect 126520 157564 126572 157616
rect 299204 157564 299256 157616
rect 326436 157836 326488 157888
rect 403808 157836 403860 157888
rect 438216 157836 438268 157888
rect 320088 157768 320140 157820
rect 325148 157768 325200 157820
rect 406752 157768 406804 157820
rect 439688 157768 439740 157820
rect 132408 157496 132460 157548
rect 299112 157496 299164 157548
rect 329196 157428 329248 157480
rect 355232 157428 355284 157480
rect 327356 157360 327408 157412
rect 356980 157360 357032 157412
rect 280988 157292 281040 157344
rect 281172 157292 281224 157344
rect 349804 157292 349856 157344
rect 125324 157224 125376 157276
rect 292396 157224 292448 157276
rect 324228 157224 324280 157276
rect 123208 157156 123260 157208
rect 290832 157156 290884 157208
rect 323124 157156 323176 157208
rect 278136 157088 278188 157140
rect 278412 157088 278464 157140
rect 338764 157088 338816 157140
rect 134892 157020 134944 157072
rect 286876 157020 286928 157072
rect 334532 157020 334584 157072
rect 135904 156952 135956 157004
rect 281448 156952 281500 157004
rect 335636 156952 335688 157004
rect 137008 156884 137060 156936
rect 281356 156884 281408 156936
rect 139216 156816 139268 156868
rect 284484 156884 284536 156936
rect 286324 156884 286376 156936
rect 336832 156884 336884 156936
rect 140688 156748 140740 156800
rect 278136 156748 278188 156800
rect 281264 156748 281316 156800
rect 338120 156816 338172 156868
rect 286600 156748 286652 156800
rect 316040 156748 316092 156800
rect 150256 156680 150308 156732
rect 281172 156680 281224 156732
rect 285956 156680 286008 156732
rect 302240 156680 302292 156732
rect 178960 156612 179012 156664
rect 282276 156612 282328 156664
rect 293500 156612 293552 156664
rect 327080 156612 327132 156664
rect 181720 156544 181772 156596
rect 282184 156544 282236 156596
rect 287428 156544 287480 156596
rect 316040 156544 316092 156596
rect 198464 156476 198516 156528
rect 276940 156476 276992 156528
rect 231860 156408 231912 156460
rect 272248 156408 272300 156460
rect 117320 156340 117372 156392
rect 284116 156340 284168 156392
rect 316684 156476 316736 156528
rect 116860 156272 116912 156324
rect 285496 156272 285548 156324
rect 286600 156272 286652 156324
rect 125416 155864 125468 155916
rect 298928 155864 298980 155916
rect 320088 155864 320140 155916
rect 283564 155796 283616 155848
rect 285956 155796 286008 155848
rect 141792 155728 141844 155780
rect 281080 155728 281132 155780
rect 281448 155728 281500 155780
rect 282368 155728 282420 155780
rect 282828 155728 282880 155780
rect 346400 155796 346452 155848
rect 286140 155728 286192 155780
rect 348700 155728 348752 155780
rect 140596 155660 140648 155712
rect 278504 155660 278556 155712
rect 278688 155660 278740 155712
rect 280068 155660 280120 155712
rect 343916 155660 343968 155712
rect 145288 155592 145340 155644
rect 282736 155592 282788 155644
rect 345112 155592 345164 155644
rect 144276 155524 144328 155576
rect 280068 155524 280120 155576
rect 283380 155524 283432 155576
rect 284208 155524 284260 155576
rect 346860 155524 346912 155576
rect 281448 155456 281500 155508
rect 341156 155456 341208 155508
rect 146392 155388 146444 155440
rect 282368 155388 282420 155440
rect 283472 155388 283524 155440
rect 284024 155388 284076 155440
rect 342812 155388 342864 155440
rect 148784 155320 148836 155372
rect 280896 155320 280948 155372
rect 286140 155320 286192 155372
rect 288900 155320 288952 155372
rect 324320 155320 324372 155372
rect 193956 155252 194008 155304
rect 279516 155252 279568 155304
rect 292948 155252 293000 155304
rect 340880 155252 340932 155304
rect 195888 155184 195940 155236
rect 276848 155184 276900 155236
rect 294328 155184 294380 155236
rect 350540 155184 350592 155236
rect 201040 155116 201092 155168
rect 276756 155116 276808 155168
rect 286048 155116 286100 155168
rect 306380 155116 306432 155168
rect 206284 155048 206336 155100
rect 273904 155048 273956 155100
rect 278688 155048 278740 155100
rect 339500 155048 339552 155100
rect 233240 154980 233292 155032
rect 272156 154980 272208 155032
rect 147772 154912 147824 154964
rect 283380 154912 283432 154964
rect 143080 154844 143132 154896
rect 283472 154844 283524 154896
rect 278688 154504 278740 154556
rect 351092 154504 351144 154556
rect 152648 154436 152700 154488
rect 299296 154436 299348 154488
rect 353300 154436 353352 154488
rect 297916 154368 297968 154420
rect 352196 154368 352248 154420
rect 154488 154300 154540 154352
rect 297824 154300 297876 154352
rect 354404 154300 354456 154352
rect 155776 154232 155828 154284
rect 286692 154232 286744 154284
rect 329196 154232 329248 154284
rect 151360 154164 151412 154216
rect 278688 154164 278740 154216
rect 157064 154096 157116 154148
rect 279976 154096 280028 154148
rect 327356 154164 327408 154216
rect 227720 154028 227772 154080
rect 271144 154028 271196 154080
rect 193220 153960 193272 154012
rect 265440 153960 265492 154012
rect 168380 153892 168432 153944
rect 261392 153892 261444 153944
rect 133880 153824 133932 153876
rect 254400 153824 254452 153876
rect 265624 153824 265676 153876
rect 275008 153824 275060 153876
rect 275100 153824 275152 153876
rect 280436 153824 280488 153876
rect 118240 153756 118292 153808
rect 283932 153756 283984 153808
rect 317696 154096 317748 154148
rect 290096 153824 290148 153876
rect 331220 153824 331272 153876
rect 153936 153688 153988 153740
rect 298192 153688 298244 153740
rect 299296 153688 299348 153740
rect 136088 153144 136140 153196
rect 271328 153144 271380 153196
rect 138940 153076 138992 153128
rect 271420 153076 271472 153128
rect 141424 153008 141476 153060
rect 271236 153008 271288 153060
rect 144368 152940 144420 152992
rect 268568 152940 268620 152992
rect 146024 152872 146076 152924
rect 268476 152872 268528 152924
rect 148416 152804 148468 152856
rect 268384 152804 268436 152856
rect 150992 152736 151044 152788
rect 268660 152736 268712 152788
rect 236000 152668 236052 152720
rect 273720 152668 273772 152720
rect 207020 152600 207072 152652
rect 268200 152600 268252 152652
rect 284392 152600 284444 152652
rect 299572 152600 299624 152652
rect 171140 152532 171192 152584
rect 261300 152532 261352 152584
rect 291660 152532 291712 152584
rect 333980 152532 334032 152584
rect 135260 152464 135312 152516
rect 254308 152464 254360 152516
rect 294604 152464 294656 152516
rect 343640 152464 343692 152516
rect 209780 151172 209832 151224
rect 268108 151172 268160 151224
rect 175280 151104 175332 151156
rect 253204 151104 253256 151156
rect 146300 151036 146352 151088
rect 257160 151036 257212 151088
rect 268200 151036 268252 151088
rect 279148 151036 279200 151088
rect 291568 151036 291620 151088
rect 338120 151036 338172 151088
rect 283288 149880 283340 149932
rect 292948 149880 293000 149932
rect 218060 149812 218112 149864
rect 269580 149812 269632 149864
rect 288808 149812 288860 149864
rect 317420 149812 317472 149864
rect 184940 149744 184992 149796
rect 264060 149744 264112 149796
rect 291476 149744 291528 149796
rect 336740 149744 336792 149796
rect 153200 149676 153252 149728
rect 249156 149676 249208 149728
rect 292856 149676 292908 149728
rect 345020 149676 345072 149728
rect 201500 148452 201552 148504
rect 266728 148452 266780 148504
rect 189080 148384 189132 148436
rect 263968 148384 264020 148436
rect 132500 148316 132552 148368
rect 251824 148316 251876 148368
rect 264336 148316 264388 148368
rect 274916 148316 274968 148368
rect 295800 148316 295852 148368
rect 357440 148316 357492 148368
rect 216680 147024 216732 147076
rect 269488 147024 269540 147076
rect 285864 147024 285916 147076
rect 303620 147024 303672 147076
rect 176660 146956 176712 147008
rect 262404 146956 262456 147008
rect 293316 146956 293368 147008
rect 328460 146956 328512 147008
rect 128360 146888 128412 146940
rect 252744 146888 252796 146940
rect 253204 146888 253256 146940
rect 273628 146888 273680 146940
rect 295708 146888 295760 146940
rect 360200 146888 360252 146940
rect 229100 145664 229152 145716
rect 272064 145664 272116 145716
rect 195980 145596 196032 145648
rect 265348 145596 265400 145648
rect 287336 145596 287388 145648
rect 310520 145596 310572 145648
rect 157340 145528 157392 145580
rect 247684 145528 247736 145580
rect 290004 145528 290056 145580
rect 332600 145528 332652 145580
rect 224960 144304 225012 144356
rect 270868 144304 270920 144356
rect 154580 144236 154632 144288
rect 258356 144236 258408 144288
rect 287244 144236 287296 144288
rect 314660 144236 314712 144288
rect 150440 144168 150492 144220
rect 257068 144168 257120 144220
rect 292764 144168 292816 144220
rect 342260 144168 342312 144220
rect 285036 144032 285088 144084
rect 287336 144032 287388 144084
rect 271144 143760 271196 143812
rect 276204 143760 276256 143812
rect 193312 142876 193364 142928
rect 265256 142876 265308 142928
rect 139400 142808 139452 142860
rect 255780 142808 255832 142860
rect 265348 142808 265400 142860
rect 277676 142808 277728 142860
rect 288716 142808 288768 142860
rect 321560 142808 321612 142860
rect 223580 141516 223632 141568
rect 270776 141516 270828 141568
rect 143540 141448 143592 141500
rect 255688 141448 255740 141500
rect 129740 141380 129792 141432
rect 254216 141380 254268 141432
rect 288624 141380 288676 141432
rect 324412 141380 324464 141432
rect 197360 140088 197412 140140
rect 266636 140088 266688 140140
rect 126980 140020 127032 140072
rect 252652 140020 252704 140072
rect 291384 140020 291436 140072
rect 335360 140020 335412 140072
rect 208400 138796 208452 138848
rect 268016 138796 268068 138848
rect 283196 138796 283248 138848
rect 291384 138796 291436 138848
rect 161480 138728 161532 138780
rect 259828 138728 259880 138780
rect 114560 138660 114612 138712
rect 250168 138660 250220 138712
rect 291292 138660 291344 138712
rect 339500 138660 339552 138712
rect 3148 137912 3200 137964
rect 82084 137912 82136 137964
rect 215300 137368 215352 137420
rect 269396 137368 269448 137420
rect 165620 137300 165672 137352
rect 259736 137300 259788 137352
rect 110420 137232 110472 137284
rect 244924 137232 244976 137284
rect 292672 137232 292724 137284
rect 346400 137232 346452 137284
rect 222200 136008 222252 136060
rect 270684 136008 270736 136060
rect 168472 135940 168524 135992
rect 261116 135940 261168 135992
rect 271236 135940 271288 135992
rect 279056 135940 279108 135992
rect 103520 135872 103572 135924
rect 243728 135872 243780 135924
rect 279516 135192 279568 135244
rect 280344 135192 280396 135244
rect 172520 134580 172572 134632
rect 261024 134580 261076 134632
rect 147680 134512 147732 134564
rect 256976 134512 257028 134564
rect 261484 134512 261536 134564
rect 276112 134512 276164 134564
rect 179420 133220 179472 133272
rect 262312 133220 262364 133272
rect 158720 133152 158772 133204
rect 258264 133152 258316 133204
rect 191840 131792 191892 131844
rect 265164 131792 265216 131844
rect 183560 131724 183612 131776
rect 263876 131724 263928 131776
rect 205640 130500 205692 130552
rect 267924 130500 267976 130552
rect 186320 130432 186372 130484
rect 263784 130432 263836 130484
rect 118700 130364 118752 130416
rect 251456 130364 251508 130416
rect 288532 130364 288584 130416
rect 318800 130364 318852 130416
rect 230480 129140 230532 129192
rect 271972 129140 272024 129192
rect 190460 129072 190512 129124
rect 265072 129072 265124 129124
rect 107660 129004 107712 129056
rect 242348 129004 242400 129056
rect 289912 129004 289964 129056
rect 325700 129004 325752 129056
rect 204260 127644 204312 127696
rect 266544 127644 266596 127696
rect 100760 127576 100812 127628
rect 246396 127576 246448 127628
rect 291200 127576 291252 127628
rect 332692 127576 332744 127628
rect 211160 126284 211212 126336
rect 267832 126284 267884 126336
rect 155960 126216 156012 126268
rect 258172 126216 258224 126268
rect 267924 126216 267976 126268
rect 278964 126216 279016 126268
rect 292580 126216 292632 126268
rect 340972 126216 341024 126268
rect 218152 124924 218204 124976
rect 269304 124924 269356 124976
rect 138020 124856 138072 124908
rect 255596 124856 255648 124908
rect 296076 124856 296128 124908
rect 354680 124856 354732 124908
rect 226340 123496 226392 123548
rect 270592 123496 270644 123548
rect 173900 123428 173952 123480
rect 260932 123428 260984 123480
rect 234712 122136 234764 122188
rect 272340 122136 272392 122188
rect 136640 122068 136692 122120
rect 254124 122068 254176 122120
rect 140780 120708 140832 120760
rect 255504 120708 255556 120760
rect 255964 120708 256016 120760
rect 274824 120708 274876 120760
rect 143632 119348 143684 119400
rect 255412 119348 255464 119400
rect 151820 117920 151872 117972
rect 256884 117920 256936 117972
rect 127072 116560 127124 116612
rect 253020 116560 253072 116612
rect 162860 115200 162912 115252
rect 259644 115200 259696 115252
rect 169760 113772 169812 113824
rect 260840 113772 260892 113824
rect 442264 113092 442316 113144
rect 579804 113092 579856 113144
rect 167000 112412 167052 112464
rect 259552 112412 259604 112464
rect 3148 111732 3200 111784
rect 84844 111732 84896 111784
rect 180800 111052 180852 111104
rect 262588 111052 262640 111104
rect 185032 109692 185084 109744
rect 263692 109692 263744 109744
rect 187700 108264 187752 108316
rect 263600 108264 263652 108316
rect 264428 108264 264480 108316
rect 277584 108264 277636 108316
rect 131120 106904 131172 106956
rect 254032 106904 254084 106956
rect 266544 106904 266596 106956
rect 276664 106904 276716 106956
rect 198740 105544 198792 105596
rect 266452 105544 266504 105596
rect 209872 104184 209924 104236
rect 267740 104184 267792 104236
rect 106280 104116 106332 104168
rect 248604 104116 248656 104168
rect 219440 102824 219492 102876
rect 269212 102824 269264 102876
rect 111800 102756 111852 102808
rect 250076 102756 250128 102808
rect 142160 101396 142212 101448
rect 255320 101396 255372 101448
rect 149060 99968 149112 100020
rect 256792 99968 256844 100020
rect 160192 98608 160244 98660
rect 258448 98608 258500 98660
rect 121460 97248 121512 97300
rect 251364 97248 251416 97300
rect 109040 94460 109092 94512
rect 249984 94460 250036 94512
rect 115940 93100 115992 93152
rect 249064 93100 249116 93152
rect 99380 91740 99432 91792
rect 247316 91740 247368 91792
rect 113824 90312 113876 90364
rect 249892 90312 249944 90364
rect 49700 88952 49752 89004
rect 239312 88952 239364 89004
rect 120080 86232 120132 86284
rect 242256 86232 242308 86284
rect 3424 85484 3476 85536
rect 80704 85484 80756 85536
rect 104900 64132 104952 64184
rect 248512 64132 248564 64184
rect 47584 33736 47636 33788
rect 237472 33736 237524 33788
rect 526444 33056 526496 33108
rect 580172 33056 580224 33108
rect 117964 25508 118016 25560
rect 250260 25508 250312 25560
rect 151912 24080 151964 24132
rect 257344 24080 257396 24132
rect 295984 24080 296036 24132
rect 347780 24080 347832 24132
rect 144920 22720 144972 22772
rect 256700 22720 256752 22772
rect 212540 21360 212592 21412
rect 269120 21360 269172 21412
rect 201592 19932 201644 19984
rect 266912 19932 266964 19984
rect 194600 18572 194652 18624
rect 264980 18572 265032 18624
rect 295616 18572 295668 18624
rect 361580 18572 361632 18624
rect 135352 17280 135404 17332
rect 254492 17280 254544 17332
rect 254032 17212 254084 17264
rect 275284 17212 275336 17264
rect 288440 17212 288492 17264
rect 322940 17212 322992 17264
rect 242900 15852 242952 15904
rect 273536 15852 273588 15904
rect 289820 15852 289872 15904
rect 330392 15852 330444 15904
rect 42800 14424 42852 14476
rect 237840 14424 237892 14476
rect 291844 14424 291896 14476
rect 305552 14424 305604 14476
rect 273904 13948 273956 14000
rect 278872 13948 278924 14000
rect 255872 13132 255924 13184
rect 264244 13132 264296 13184
rect 81624 13064 81676 13116
rect 242164 13064 242216 13116
rect 260012 13064 260064 13116
rect 277492 13064 277544 13116
rect 287152 13064 287204 13116
rect 312176 13064 312228 13116
rect 278136 12452 278188 12504
rect 280252 12452 280304 12504
rect 280712 12452 280764 12504
rect 281908 12452 281960 12504
rect 160100 11772 160152 11824
rect 161296 11772 161348 11824
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 234620 11772 234672 11824
rect 235816 11772 235868 11824
rect 102140 11704 102192 11756
rect 246304 11704 246356 11756
rect 287060 11704 287112 11756
rect 316224 11704 316276 11756
rect 439136 11840 439188 11892
rect 439044 11636 439096 11688
rect 270776 10480 270828 10532
rect 278044 10480 278096 10532
rect 237656 10344 237708 10396
rect 273444 10344 273496 10396
rect 53012 10276 53064 10328
rect 239220 10276 239272 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 283104 9120 283156 9172
rect 292580 9120 292632 9172
rect 289360 9052 289412 9104
rect 410800 9052 410852 9104
rect 241704 8984 241756 9036
rect 273352 8984 273404 9036
rect 285404 8984 285456 9036
rect 411904 8984 411956 9036
rect 123484 8916 123536 8968
rect 243544 8916 243596 8968
rect 248788 8916 248840 8968
rect 262864 8916 262916 8968
rect 288072 8916 288124 8968
rect 414296 8916 414348 8968
rect 281816 8236 281868 8288
rect 283104 8236 283156 8288
rect 240508 7624 240560 7676
rect 273260 7624 273312 7676
rect 227536 7556 227588 7608
rect 270500 7556 270552 7608
rect 276020 7556 276072 7608
rect 280528 7556 280580 7608
rect 299572 7556 299624 7608
rect 300768 7556 300820 7608
rect 283012 6944 283064 6996
rect 288992 6944 289044 6996
rect 3424 6808 3476 6860
rect 40684 6808 40736 6860
rect 295524 6740 295576 6792
rect 358728 6740 358780 6792
rect 291108 6672 291160 6724
rect 378876 6672 378928 6724
rect 291016 6604 291068 6656
rect 385960 6604 386012 6656
rect 287888 6536 287940 6588
rect 400128 6536 400180 6588
rect 289728 6468 289780 6520
rect 403624 6468 403676 6520
rect 284944 6400 284996 6452
rect 294880 6400 294932 6452
rect 294972 6400 295024 6452
rect 413100 6400 413152 6452
rect 287980 6332 288032 6384
rect 407212 6332 407264 6384
rect 290648 6264 290700 6316
rect 416688 6264 416740 6316
rect 247592 6196 247644 6248
rect 274732 6196 274784 6248
rect 292488 6196 292540 6248
rect 420184 6196 420236 6248
rect 119896 6128 119948 6180
rect 251272 6128 251324 6180
rect 257068 6128 257120 6180
rect 276296 6128 276348 6180
rect 286968 6128 287020 6180
rect 415492 6128 415544 6180
rect 278320 5516 278372 5568
rect 279424 5516 279476 5568
rect 284300 5176 284352 5228
rect 298468 5176 298520 5228
rect 285772 5108 285824 5160
rect 307944 5108 307996 5160
rect 294144 5040 294196 5092
rect 350448 5040 350500 5092
rect 294236 4972 294288 5024
rect 354036 4972 354088 5024
rect 296720 4904 296772 4956
rect 364616 4904 364668 4956
rect 244096 4836 244148 4888
rect 275192 4836 275244 4888
rect 298560 4836 298612 4888
rect 371700 4836 371752 4888
rect 177856 4768 177908 4820
rect 260104 4768 260156 4820
rect 264152 4768 264204 4820
rect 277768 4768 277820 4820
rect 282920 4768 282972 4820
rect 290188 4768 290240 4820
rect 299388 4768 299440 4820
rect 377680 4768 377732 4820
rect 281724 4156 281776 4208
rect 285404 4156 285456 4208
rect 2872 4088 2924 4140
rect 7564 4088 7616 4140
rect 45468 4088 45520 4140
rect 46296 4088 46348 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 293316 4088 293368 4140
rect 296076 4088 296128 4140
rect 239312 4020 239364 4072
rect 253204 4020 253256 4072
rect 294052 4020 294104 4072
rect 349252 4088 349304 4140
rect 430856 4088 430908 4140
rect 437664 4088 437716 4140
rect 460204 4088 460256 4140
rect 462780 4088 462832 4140
rect 468484 4088 468536 4140
rect 471060 4088 471112 4140
rect 536196 4088 536248 4140
rect 538404 4088 538456 4140
rect 566464 4088 566516 4140
rect 569132 4088 569184 4140
rect 298284 4020 298336 4072
rect 352840 4020 352892 4072
rect 429660 4020 429712 4072
rect 438860 4020 438912 4072
rect 92756 3952 92808 4004
rect 95884 3952 95936 4004
rect 135260 3952 135312 4004
rect 136456 3952 136508 4004
rect 164884 3952 164936 4004
rect 259460 3952 259512 4004
rect 273628 3952 273680 4004
rect 279516 3952 279568 4004
rect 295340 3952 295392 4004
rect 110512 3884 110564 3936
rect 113824 3884 113876 3936
rect 124680 3884 124732 3936
rect 243636 3884 243688 3936
rect 293960 3884 294012 3936
rect 298192 3884 298244 3936
rect 356336 3952 356388 4004
rect 428464 3952 428516 4004
rect 439044 3952 439096 4004
rect 298744 3884 298796 3936
rect 365812 3884 365864 3936
rect 426164 3884 426216 3936
rect 437572 3884 437624 3936
rect 476764 3884 476816 3936
rect 480536 3884 480588 3936
rect 117596 3816 117648 3868
rect 239404 3816 239456 3868
rect 245200 3816 245252 3868
rect 255964 3816 256016 3868
rect 19432 3748 19484 3800
rect 39304 3748 39356 3800
rect 102232 3748 102284 3800
rect 248696 3748 248748 3800
rect 11152 3680 11204 3732
rect 46204 3680 46256 3732
rect 15936 3612 15988 3664
rect 50344 3612 50396 3664
rect 1676 3544 1728 3596
rect 4804 3544 4856 3596
rect 4068 3476 4120 3528
rect 10324 3544 10376 3596
rect 12348 3544 12400 3596
rect 13084 3544 13136 3596
rect 25320 3544 25372 3596
rect 68284 3680 68336 3732
rect 98644 3680 98696 3732
rect 247408 3680 247460 3732
rect 7656 3476 7708 3528
rect 8944 3476 8996 3528
rect 20628 3476 20680 3528
rect 64144 3612 64196 3664
rect 75000 3612 75052 3664
rect 88984 3612 89036 3664
rect 97448 3612 97500 3664
rect 247224 3612 247276 3664
rect 251272 3612 251324 3664
rect 261484 3816 261536 3868
rect 295432 3816 295484 3868
rect 359924 3816 359976 3868
rect 427268 3816 427320 3868
rect 439320 3816 439372 3868
rect 516784 3816 516836 3868
rect 519544 3816 519596 3868
rect 574744 3816 574796 3868
rect 577412 3816 577464 3868
rect 70308 3544 70360 3596
rect 71044 3544 71096 3596
rect 56048 3476 56100 3528
rect 57244 3476 57296 3528
rect 60740 3476 60792 3528
rect 61660 3476 61712 3528
rect 65524 3476 65576 3528
rect 66904 3476 66956 3528
rect 67916 3476 67968 3528
rect 82176 3544 82228 3596
rect 96252 3544 96304 3596
rect 97264 3544 97316 3596
rect 102140 3544 102192 3596
rect 103336 3544 103388 3596
rect 103428 3544 103480 3596
rect 247500 3544 247552 3596
rect 249984 3544 250036 3596
rect 264336 3748 264388 3800
rect 288348 3748 288400 3800
rect 367008 3748 367060 3800
rect 424968 3748 425020 3800
rect 437480 3748 437532 3800
rect 259460 3680 259512 3732
rect 269764 3680 269816 3732
rect 295248 3680 295300 3732
rect 384764 3680 384816 3732
rect 423772 3680 423824 3732
rect 437848 3680 437900 3732
rect 295156 3612 295208 3664
rect 402520 3612 402572 3664
rect 422576 3612 422628 3664
rect 438952 3612 439004 3664
rect 258264 3544 258316 3596
rect 260196 3544 260248 3596
rect 267924 3544 267976 3596
rect 268476 3544 268528 3596
rect 77300 3476 77352 3528
rect 78220 3476 78272 3528
rect 83280 3476 83332 3528
rect 244372 3476 244424 3528
rect 251180 3476 251232 3528
rect 252376 3476 252428 3528
rect 253480 3476 253532 3528
rect 271144 3544 271196 3596
rect 286324 3544 286376 3596
rect 297272 3544 297324 3596
rect 298008 3544 298060 3596
rect 406016 3544 406068 3596
rect 421380 3544 421432 3596
rect 434352 3544 434404 3596
rect 434444 3544 434496 3596
rect 439136 3544 439188 3596
rect 442356 3544 442408 3596
rect 447416 3544 447468 3596
rect 450544 3544 450596 3596
rect 270040 3476 270092 3528
rect 271236 3476 271288 3528
rect 272432 3476 272484 3528
rect 273904 3476 273956 3528
rect 293868 3476 293920 3528
rect 409604 3476 409656 3528
rect 418988 3476 419040 3528
rect 438032 3476 438084 3528
rect 440332 3476 440384 3528
rect 441528 3476 441580 3528
rect 448612 3476 448664 3528
rect 449808 3476 449860 3528
rect 453304 3544 453356 3596
rect 455696 3544 455748 3596
rect 458824 3544 458876 3596
rect 465172 3544 465224 3596
rect 467104 3544 467156 3596
rect 469864 3544 469916 3596
rect 454500 3476 454552 3528
rect 456892 3476 456944 3528
rect 458088 3476 458140 3528
rect 462964 3476 463016 3528
rect 471244 3476 471296 3528
rect 473452 3476 473504 3528
rect 475384 3544 475436 3596
rect 476948 3544 477000 3596
rect 478236 3544 478288 3596
rect 484032 3544 484084 3596
rect 500224 3544 500276 3596
rect 501788 3544 501840 3596
rect 548524 3544 548576 3596
rect 550272 3544 550324 3596
rect 479340 3476 479392 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 496084 3476 496136 3528
rect 497096 3476 497148 3528
rect 514024 3476 514076 3528
rect 515956 3476 516008 3528
rect 522304 3476 522356 3528
rect 524236 3476 524288 3528
rect 538864 3476 538916 3528
rect 540796 3476 540848 3528
rect 549904 3476 549956 3528
rect 551468 3476 551520 3528
rect 563704 3476 563756 3528
rect 566832 3476 566884 3528
rect 581000 3476 581052 3528
rect 581828 3476 581880 3528
rect 572 3408 624 3460
rect 25504 3408 25556 3460
rect 27620 3408 27672 3460
rect 28540 3408 28592 3460
rect 33600 3408 33652 3460
rect 35164 3408 35216 3460
rect 38384 3408 38436 3460
rect 39396 3408 39448 3460
rect 39580 3408 39632 3460
rect 43444 3408 43496 3460
rect 46664 3408 46716 3460
rect 47584 3408 47636 3460
rect 47860 3408 47912 3460
rect 48964 3408 49016 3460
rect 79692 3408 79744 3460
rect 244556 3408 244608 3460
rect 246396 3408 246448 3460
rect 95148 3340 95200 3392
rect 103428 3340 103480 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 285588 3408 285640 3460
rect 401324 3408 401376 3460
rect 417884 3408 417936 3460
rect 437756 3408 437808 3460
rect 445116 3408 445168 3460
rect 265624 3340 265676 3392
rect 285680 3340 285732 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332692 3340 332744 3392
rect 333888 3340 333940 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 434352 3340 434404 3392
rect 439228 3340 439280 3392
rect 446404 3340 446456 3392
rect 452108 3340 452160 3392
rect 493324 3340 493376 3392
rect 499396 3340 499448 3392
rect 514116 3408 514168 3460
rect 514760 3408 514812 3460
rect 520924 3408 520976 3460
rect 523040 3408 523092 3460
rect 527916 3408 527968 3460
rect 533712 3408 533764 3460
rect 543004 3408 543056 3460
rect 549076 3408 549128 3460
rect 526628 3340 526680 3392
rect 554044 3340 554096 3392
rect 559748 3340 559800 3392
rect 262956 3272 263008 3324
rect 264428 3272 264480 3324
rect 454684 3272 454736 3324
rect 459192 3272 459244 3324
rect 509884 3272 509936 3324
rect 513564 3272 513616 3324
rect 571984 3272 572036 3324
rect 573916 3272 573968 3324
rect 6460 3204 6512 3256
rect 7564 3204 7616 3256
rect 51356 3204 51408 3256
rect 53104 3204 53156 3256
rect 85672 3136 85724 3188
rect 93124 3136 93176 3188
rect 114008 3136 114060 3188
rect 117964 3136 118016 3188
rect 277124 3136 277176 3188
rect 278136 3136 278188 3188
rect 281632 3136 281684 3188
rect 284300 3136 284352 3188
rect 485044 3136 485096 3188
rect 487620 3136 487672 3188
rect 534724 3136 534776 3188
rect 537208 3136 537260 3188
rect 560944 3136 560996 3188
rect 563244 3136 563296 3188
rect 567844 3136 567896 3188
rect 570328 3136 570380 3188
rect 570604 3068 570656 3120
rect 572720 3068 572772 3120
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 503076 3000 503128 3052
rect 505376 3000 505428 3052
rect 552756 3000 552808 3052
rect 554964 3000 555016 3052
rect 563796 3000 563848 3052
rect 565636 3000 565688 3052
rect 8760 2932 8812 2984
rect 14464 2932 14516 2984
rect 526536 2932 526588 2984
rect 527824 2932 527876 2984
rect 540244 2932 540296 2984
rect 541992 2932 542044 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 21364 700324 21416 700330
rect 21364 700266 21416 700272
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501362 3372 501735
rect 3332 501356 3384 501362
rect 3332 501298 3384 501304
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 2870 449576 2926 449585
rect 2870 449511 2926 449520
rect 2884 447846 2912 449511
rect 3436 449274 3464 619103
rect 3514 606112 3570 606121
rect 3514 606047 3516 606056
rect 3568 606047 3570 606056
rect 3516 606018 3568 606024
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3424 449268 3476 449274
rect 3424 449210 3476 449216
rect 3528 449206 3556 566879
rect 3606 553888 3662 553897
rect 3606 553823 3662 553832
rect 3620 553450 3648 553823
rect 3608 553444 3660 553450
rect 3608 553386 3660 553392
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3620 450566 3648 514791
rect 4816 467158 4844 683674
rect 18604 670744 18656 670750
rect 18604 670686 18656 670692
rect 17224 656940 17276 656946
rect 17224 656882 17276 656888
rect 13084 632120 13136 632126
rect 13084 632062 13136 632068
rect 7564 606076 7616 606082
rect 7564 606018 7616 606024
rect 4804 467152 4856 467158
rect 4804 467094 4856 467100
rect 7576 458862 7604 606018
rect 10324 579692 10376 579698
rect 10324 579634 10376 579640
rect 8944 501356 8996 501362
rect 8944 501298 8996 501304
rect 7564 458856 7616 458862
rect 7564 458798 7616 458804
rect 8956 457502 8984 501298
rect 10336 469878 10364 579634
rect 10324 469872 10376 469878
rect 10324 469814 10376 469820
rect 13096 468518 13124 632062
rect 14464 527196 14516 527202
rect 14464 527138 14516 527144
rect 14476 471306 14504 527138
rect 14464 471300 14516 471306
rect 14464 471242 14516 471248
rect 13084 468512 13136 468518
rect 13084 468454 13136 468460
rect 17236 460222 17264 656882
rect 17224 460216 17276 460222
rect 17224 460158 17276 460164
rect 8944 457496 8996 457502
rect 8944 457438 8996 457444
rect 18616 456074 18644 670686
rect 21376 474026 21404 700266
rect 22744 553444 22796 553450
rect 22744 553386 22796 553392
rect 21364 474020 21416 474026
rect 21364 473962 21416 473968
rect 22756 464370 22784 553386
rect 22744 464364 22796 464370
rect 22744 464306 22796 464312
rect 18604 456068 18656 456074
rect 18604 456010 18656 456016
rect 3608 450560 3660 450566
rect 3608 450502 3660 450508
rect 23492 449342 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 23480 449336 23532 449342
rect 23480 449278 23532 449284
rect 3516 449200 3568 449206
rect 3516 449142 3568 449148
rect 40052 447914 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 472666 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 71780 472660 71832 472666
rect 71780 472602 71832 472608
rect 88352 449478 88380 702406
rect 88340 449472 88392 449478
rect 88340 449414 88392 449420
rect 104912 447982 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 448050 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 449614 153240 702406
rect 169772 465730 169800 702406
rect 169760 465724 169812 465730
rect 169760 465666 169812 465672
rect 153200 449608 153252 449614
rect 153200 449550 153252 449556
rect 201512 448118 201540 702986
rect 217968 700324 218020 700330
rect 217968 700266 218020 700272
rect 217874 516896 217930 516905
rect 217874 516831 217930 516840
rect 217782 515944 217838 515953
rect 217782 515879 217838 515888
rect 217598 513768 217654 513777
rect 217598 513703 217654 513712
rect 217322 488336 217378 488345
rect 217322 488271 217378 488280
rect 217336 478922 217364 488271
rect 217506 488064 217562 488073
rect 217506 487999 217562 488008
rect 217324 478916 217376 478922
rect 217324 478858 217376 478864
rect 217520 476814 217548 487999
rect 217612 478242 217640 513703
rect 217690 489968 217746 489977
rect 217690 489903 217746 489912
rect 217600 478236 217652 478242
rect 217600 478178 217652 478184
rect 217508 476808 217560 476814
rect 217508 476750 217560 476756
rect 217704 453354 217732 489903
rect 217796 474094 217824 515879
rect 217784 474088 217836 474094
rect 217784 474030 217836 474036
rect 217888 472734 217916 516831
rect 217876 472728 217928 472734
rect 217876 472670 217928 472676
rect 217692 453348 217744 453354
rect 217692 453290 217744 453296
rect 201500 448112 201552 448118
rect 201500 448054 201552 448060
rect 136640 448044 136692 448050
rect 136640 447986 136692 447992
rect 104900 447976 104952 447982
rect 104900 447918 104952 447924
rect 40040 447908 40092 447914
rect 40040 447850 40092 447856
rect 2872 447840 2924 447846
rect 2872 447782 2924 447788
rect 217980 446690 218008 700266
rect 218072 478174 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700330 235212 703520
rect 267660 700330 267688 703520
rect 283852 700398 283880 703520
rect 300136 700466 300164 703520
rect 332520 700534 332548 703520
rect 348804 700602 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 357624 700596 357676 700602
rect 357624 700538 357676 700544
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 357532 700460 357584 700466
rect 357532 700402 357584 700408
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 357440 700324 357492 700330
rect 357440 700266 357492 700272
rect 219162 512816 219218 512825
rect 219162 512751 219218 512760
rect 219070 508192 219126 508201
rect 219070 508127 219126 508136
rect 219084 478310 219112 508127
rect 219072 478304 219124 478310
rect 219072 478246 219124 478252
rect 218060 478168 218112 478174
rect 218060 478110 218112 478116
rect 219176 475386 219204 512751
rect 219346 511048 219402 511057
rect 219346 510983 219402 510992
rect 219254 509960 219310 509969
rect 219254 509895 219310 509904
rect 219164 475380 219216 475386
rect 219164 475322 219216 475328
rect 219268 461650 219296 509895
rect 219256 461644 219308 461650
rect 219256 461586 219308 461592
rect 219360 451926 219388 510983
rect 220084 478916 220136 478922
rect 220084 478858 220136 478864
rect 219348 451920 219400 451926
rect 219348 451862 219400 451868
rect 217968 446684 218020 446690
rect 217968 446626 218020 446632
rect 220096 446486 220124 478858
rect 238760 478304 238812 478310
rect 238760 478246 238812 478252
rect 238772 476898 238800 478246
rect 248512 478236 248564 478242
rect 248512 478178 248564 478184
rect 309140 478236 309192 478242
rect 309140 478178 309192 478184
rect 247038 477456 247094 477465
rect 247038 477391 247094 477400
rect 242898 477048 242954 477057
rect 247052 477018 247080 477391
rect 248418 477048 248474 477057
rect 242898 476983 242954 476992
rect 245752 477012 245804 477018
rect 238680 476870 238800 476898
rect 230480 476808 230532 476814
rect 230480 476750 230532 476756
rect 230492 460934 230520 476750
rect 233240 476740 233292 476746
rect 233240 476682 233292 476688
rect 231860 476332 231912 476338
rect 231860 476274 231912 476280
rect 230492 460906 230704 460934
rect 220084 446480 220136 446486
rect 220084 446422 220136 446428
rect 230388 446480 230440 446486
rect 230388 446422 230440 446428
rect 229836 446004 229888 446010
rect 229836 445946 229888 445952
rect 229744 445936 229796 445942
rect 229744 445878 229796 445884
rect 228364 445868 228416 445874
rect 228364 445810 228416 445816
rect 7564 445188 7616 445194
rect 7564 445130 7616 445136
rect 3516 443692 3568 443698
rect 3516 443634 3568 443640
rect 3424 440904 3476 440910
rect 3424 440846 3476 440852
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3056 372564 3108 372570
rect 3056 372506 3108 372512
rect 3068 371385 3096 372506
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3148 215280 3200 215286
rect 3148 215222 3200 215228
rect 3160 214985 3188 215222
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3436 149841 3464 440846
rect 3528 201929 3556 443634
rect 3608 442264 3660 442270
rect 3608 442206 3660 442212
rect 3620 358465 3648 442206
rect 7576 423638 7604 445130
rect 225696 445120 225748 445126
rect 225696 445062 225748 445068
rect 224224 444984 224276 444990
rect 224224 444926 224276 444932
rect 93216 444712 93268 444718
rect 93216 444654 93268 444660
rect 86224 444644 86276 444650
rect 86224 444586 86276 444592
rect 84844 444576 84896 444582
rect 84844 444518 84896 444524
rect 82084 444508 82136 444514
rect 82084 444450 82136 444456
rect 80704 443012 80756 443018
rect 80704 442954 80756 442960
rect 7564 423632 7616 423638
rect 7564 423574 7616 423580
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 68284 308984 68336 308990
rect 68284 308926 68336 308932
rect 50344 308916 50396 308922
rect 50344 308858 50396 308864
rect 46204 308780 46256 308786
rect 46204 308722 46256 308728
rect 43444 308712 43496 308718
rect 43444 308654 43496 308660
rect 39304 308644 39356 308650
rect 39304 308586 39356 308592
rect 35900 308576 35952 308582
rect 35900 308518 35952 308524
rect 27620 308508 27672 308514
rect 27620 308450 27672 308456
rect 23480 308440 23532 308446
rect 23480 308382 23532 308388
rect 7564 304292 7616 304298
rect 7564 304234 7616 304240
rect 4160 262880 4212 262886
rect 4160 262822 4212 262828
rect 3700 247716 3752 247722
rect 3700 247658 3752 247664
rect 3608 244316 3660 244322
rect 3608 244258 3660 244264
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 164212 3568 164218
rect 3516 164154 3568 164160
rect 3528 162897 3556 164154
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3148 137964 3200 137970
rect 3148 137906 3200 137912
rect 3160 136785 3188 137906
rect 3146 136776 3202 136785
rect 3146 136711 3202 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3424 85536 3476 85542
rect 3424 85478 3476 85484
rect 3436 84697 3464 85478
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3620 45529 3648 244258
rect 3712 97617 3740 247658
rect 3698 97608 3754 97617
rect 3698 97543 3754 97552
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 4172 16574 4200 262822
rect 4804 249076 4856 249082
rect 4804 249018 4856 249024
rect 4172 16546 4752 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 2884 480 2912 4082
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4724 3482 4752 16546
rect 4816 3602 4844 249018
rect 7576 4146 7604 304234
rect 8944 302932 8996 302938
rect 8944 302874 8996 302880
rect 7656 246356 7708 246362
rect 7656 246298 7708 246304
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 3618 7696 246298
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 7576 3590 7696 3618
rect 4080 480 4108 3470
rect 4724 3454 5304 3482
rect 5276 480 5304 3454
rect 7576 3262 7604 3590
rect 8956 3534 8984 302874
rect 10324 298784 10376 298790
rect 10324 298726 10376 298732
rect 9680 287700 9732 287706
rect 9680 287642 9732 287648
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 6460 3256 6512 3262
rect 6460 3198 6512 3204
rect 7564 3256 7616 3262
rect 7564 3198 7616 3204
rect 6472 480 6500 3198
rect 7668 480 7696 3470
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8772 480 8800 2926
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 287642
rect 10336 3602 10364 298726
rect 13084 289128 13136 289134
rect 13084 289070 13136 289076
rect 12440 251864 12492 251870
rect 12440 251806 12492 251812
rect 12452 16574 12480 251806
rect 12452 16546 13032 16574
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11164 480 11192 3674
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13004 3482 13032 16546
rect 13096 3602 13124 289070
rect 16580 283620 16632 283626
rect 16580 283562 16632 283568
rect 14464 273964 14516 273970
rect 14464 273906 14516 273912
rect 13820 260160 13872 260166
rect 13820 260102 13872 260108
rect 13832 16574 13860 260102
rect 13832 16546 14320 16574
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13004 3454 13584 3482
rect 13556 480 13584 3454
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2990 14504 273906
rect 16592 16574 16620 283562
rect 20720 282192 20772 282198
rect 20720 282134 20772 282140
rect 17960 244928 18012 244934
rect 17960 244870 18012 244876
rect 16592 16546 17080 16574
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 15948 480 15976 3606
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 244870
rect 20732 16574 20760 282134
rect 22100 244996 22152 245002
rect 22100 244938 22152 244944
rect 22112 16574 22140 244938
rect 23492 16574 23520 308382
rect 25504 307080 25556 307086
rect 25504 307022 25556 307028
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 19432 3800 19484 3806
rect 19432 3742 19484 3748
rect 19444 480 19472 3742
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 480 20668 3470
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 480 25360 3538
rect 25516 3466 25544 307022
rect 26240 280832 26292 280838
rect 26240 280774 26292 280780
rect 25504 3460 25556 3466
rect 25504 3402 25556 3408
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 280774
rect 27632 3466 27660 308450
rect 30380 291848 30432 291854
rect 30380 291790 30432 291796
rect 29000 279472 29052 279478
rect 29000 279414 29052 279420
rect 27712 253224 27764 253230
rect 27712 253166 27764 253172
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27724 480 27752 253166
rect 29012 16574 29040 279414
rect 30392 16574 30420 291790
rect 34520 284980 34572 284986
rect 34520 284922 34572 284928
rect 31760 261520 31812 261526
rect 31760 261462 31812 261468
rect 31772 16574 31800 261462
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3402
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 480 33640 3402
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 284922
rect 35164 278044 35216 278050
rect 35164 277986 35216 277992
rect 35176 3466 35204 277986
rect 35912 6914 35940 308518
rect 35992 276684 36044 276690
rect 35992 276626 36044 276632
rect 36004 16574 36032 276626
rect 36004 16546 36768 16574
rect 35912 6886 36032 6914
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 39316 3806 39344 308586
rect 40682 305688 40738 305697
rect 40682 305623 40738 305632
rect 40040 300144 40092 300150
rect 40040 300086 40092 300092
rect 39396 250504 39448 250510
rect 39396 250446 39448 250452
rect 39304 3800 39356 3806
rect 39304 3742 39356 3748
rect 39408 3466 39436 250446
rect 40052 16574 40080 300086
rect 40052 16546 40264 16574
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 39396 3460 39448 3466
rect 39396 3402 39448 3408
rect 39580 3460 39632 3466
rect 39580 3402 39632 3408
rect 38396 480 38424 3402
rect 39592 480 39620 3402
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 40696 6866 40724 305623
rect 41420 290488 41472 290494
rect 41420 290430 41472 290436
rect 41432 16574 41460 290430
rect 41432 16546 41920 16574
rect 40684 6860 40736 6866
rect 40684 6802 40736 6808
rect 41892 480 41920 16546
rect 42800 14476 42852 14482
rect 42800 14418 42852 14424
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 14418
rect 43456 3466 43484 308654
rect 44180 275324 44232 275330
rect 44180 275266 44232 275272
rect 44192 16574 44220 275266
rect 44192 16546 44312 16574
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 44284 480 44312 16546
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 45480 480 45508 4082
rect 46216 3738 46244 308722
rect 48964 301504 49016 301510
rect 48964 301446 49016 301452
rect 46296 286340 46348 286346
rect 46296 286282 46348 286288
rect 46308 4146 46336 286282
rect 48320 272536 48372 272542
rect 48320 272478 48372 272484
rect 47584 33788 47636 33794
rect 47584 33730 47636 33736
rect 46296 4140 46348 4146
rect 46296 4082 46348 4088
rect 46204 3732 46256 3738
rect 46204 3674 46256 3680
rect 47596 3466 47624 33730
rect 48332 16574 48360 272478
rect 48332 16546 48544 16574
rect 46664 3460 46716 3466
rect 46664 3402 46716 3408
rect 47584 3460 47636 3466
rect 47584 3402 47636 3408
rect 47860 3460 47912 3466
rect 47860 3402 47912 3408
rect 46676 480 46704 3402
rect 47872 480 47900 3402
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 48976 3466 49004 301446
rect 49700 89004 49752 89010
rect 49700 88946 49752 88952
rect 49712 16574 49740 88946
rect 49712 16546 50200 16574
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 50172 480 50200 16546
rect 50356 3670 50384 308858
rect 64144 308848 64196 308854
rect 64144 308790 64196 308796
rect 57980 307148 58032 307154
rect 57980 307090 58032 307096
rect 53104 300212 53156 300218
rect 53104 300154 53156 300160
rect 52460 271176 52512 271182
rect 52460 271118 52512 271124
rect 52472 16574 52500 271118
rect 52472 16546 52592 16574
rect 50344 3664 50396 3670
rect 50344 3606 50396 3612
rect 51356 3256 51408 3262
rect 51356 3198 51408 3204
rect 51368 480 51396 3198
rect 52564 480 52592 16546
rect 53012 10328 53064 10334
rect 53012 10270 53064 10276
rect 53024 490 53052 10270
rect 53116 3262 53144 300154
rect 53840 298852 53892 298858
rect 53840 298794 53892 298800
rect 53852 16574 53880 298794
rect 56600 289196 56652 289202
rect 56600 289138 56652 289144
rect 56612 16574 56640 289138
rect 57244 269816 57296 269822
rect 57244 269758 57296 269764
rect 53852 16546 54984 16574
rect 56612 16546 56824 16574
rect 53104 3256 53156 3262
rect 53104 3198 53156 3204
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53024 462 53328 490
rect 54956 480 54984 16546
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56060 480 56088 3470
rect 53300 354 53328 462
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3534 57284 269758
rect 57992 16574 58020 307090
rect 60740 297492 60792 297498
rect 60740 297434 60792 297440
rect 59360 268388 59412 268394
rect 59360 268330 59412 268336
rect 57992 16546 58480 16574
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 268330
rect 60752 3534 60780 297434
rect 62120 297424 62172 297430
rect 62120 297366 62172 297372
rect 60832 283688 60884 283694
rect 60832 283630 60884 283636
rect 60740 3528 60792 3534
rect 60740 3470 60792 3476
rect 60844 480 60872 283630
rect 62132 16574 62160 297366
rect 63500 258732 63552 258738
rect 63500 258674 63552 258680
rect 63512 16574 63540 258674
rect 62132 16546 63264 16574
rect 63512 16546 64092 16574
rect 61660 3528 61712 3534
rect 61660 3470 61712 3476
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3470
rect 63236 480 63264 16546
rect 64064 3482 64092 16546
rect 64156 3670 64184 308790
rect 66904 295996 66956 296002
rect 66904 295938 66956 295944
rect 66260 265668 66312 265674
rect 66260 265610 66312 265616
rect 66272 16574 66300 265610
rect 66272 16546 66760 16574
rect 64144 3664 64196 3670
rect 64144 3606 64196 3612
rect 65524 3528 65576 3534
rect 64064 3454 64368 3482
rect 65524 3470 65576 3476
rect 64340 480 64368 3454
rect 65536 480 65564 3470
rect 66732 480 66760 16546
rect 66916 3534 66944 295938
rect 68296 3738 68324 308926
rect 80060 307216 80112 307222
rect 80060 307158 80112 307164
rect 77300 303000 77352 303006
rect 77300 302942 77352 302948
rect 71044 296064 71096 296070
rect 71044 296006 71096 296012
rect 69020 294636 69072 294642
rect 69020 294578 69072 294584
rect 69032 16574 69060 294578
rect 70400 282260 70452 282266
rect 70400 282202 70452 282208
rect 70412 16574 70440 282202
rect 69032 16546 69152 16574
rect 70412 16546 70992 16574
rect 68284 3732 68336 3738
rect 68284 3674 68336 3680
rect 66904 3528 66956 3534
rect 66904 3470 66956 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 67928 480 67956 3470
rect 69124 480 69152 16546
rect 70308 3596 70360 3602
rect 70308 3538 70360 3544
rect 70320 480 70348 3538
rect 70964 3482 70992 16546
rect 71056 3602 71084 296006
rect 71780 291916 71832 291922
rect 71780 291858 71832 291864
rect 71792 16574 71820 291858
rect 75920 290556 75972 290562
rect 75920 290498 75972 290504
rect 75184 264240 75236 264246
rect 75184 264182 75236 264188
rect 71792 16546 72648 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 75196 4146 75224 264182
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 73816 480 73844 4082
rect 75000 3664 75052 3670
rect 75000 3606 75052 3612
rect 75012 480 75040 3606
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 290498
rect 77312 3534 77340 302942
rect 77392 262948 77444 262954
rect 77392 262890 77444 262896
rect 77300 3528 77352 3534
rect 77300 3470 77352 3476
rect 77404 480 77432 262890
rect 80072 16574 80100 307158
rect 80716 85542 80744 442954
rect 82096 137970 82124 444450
rect 82176 305652 82228 305658
rect 82176 305594 82228 305600
rect 82084 137964 82136 137970
rect 82084 137906 82136 137912
rect 80704 85536 80756 85542
rect 80704 85478 80756 85484
rect 80072 16546 80928 16574
rect 78220 3528 78272 3534
rect 78220 3470 78272 3476
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3470
rect 79692 3460 79744 3466
rect 79692 3402 79744 3408
rect 79704 480 79732 3402
rect 80900 480 80928 16546
rect 81624 13116 81676 13122
rect 81624 13058 81676 13064
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 13058
rect 82188 3602 82216 305594
rect 84200 261588 84252 261594
rect 84200 261530 84252 261536
rect 82176 3596 82228 3602
rect 82176 3538 82228 3544
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 83292 480 83320 3470
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 261530
rect 84856 111790 84884 444518
rect 85580 303068 85632 303074
rect 85580 303010 85632 303016
rect 84844 111784 84896 111790
rect 84844 111726 84896 111732
rect 85592 16574 85620 303010
rect 86236 164218 86264 444586
rect 88984 304360 89036 304366
rect 88984 304302 89036 304308
rect 86960 293276 87012 293282
rect 86960 293218 87012 293224
rect 86224 164212 86276 164218
rect 86224 164154 86276 164160
rect 86972 16574 87000 293218
rect 88340 279540 88392 279546
rect 88340 279482 88392 279488
rect 88352 16574 88380 279482
rect 85592 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 88932 16574
rect 85672 3188 85724 3194
rect 85672 3130 85724 3136
rect 85684 480 85712 3130
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 88904 3482 88932 16546
rect 88996 3670 89024 304302
rect 89720 286408 89772 286414
rect 89720 286350 89772 286356
rect 89732 16574 89760 286350
rect 93124 280900 93176 280906
rect 93124 280842 93176 280848
rect 91100 260228 91152 260234
rect 91100 260170 91152 260176
rect 91112 16574 91140 260170
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 88984 3664 89036 3670
rect 88984 3606 89036 3612
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92756 4004 92808 4010
rect 92756 3946 92808 3952
rect 92768 480 92796 3946
rect 93136 3194 93164 280842
rect 93228 215286 93256 444654
rect 221464 443352 221516 443358
rect 221464 443294 221516 443300
rect 220084 443216 220136 443222
rect 220084 443158 220136 443164
rect 98644 443148 98696 443154
rect 98644 443090 98696 443096
rect 95976 443080 96028 443086
rect 95976 443022 96028 443028
rect 95884 301640 95936 301646
rect 95884 301582 95936 301588
rect 93860 301572 93912 301578
rect 93860 301514 93912 301520
rect 93216 215280 93268 215286
rect 93216 215222 93268 215228
rect 93872 16574 93900 301514
rect 93872 16546 93992 16574
rect 93124 3188 93176 3194
rect 93124 3130 93176 3136
rect 93964 480 93992 16546
rect 95896 4010 95924 301582
rect 95988 189038 96016 443022
rect 97264 309052 97316 309058
rect 97264 308994 97316 309000
rect 95976 189032 96028 189038
rect 95976 188974 96028 188980
rect 95884 4004 95936 4010
rect 95884 3946 95936 3952
rect 97276 3602 97304 308994
rect 97908 244384 97960 244390
rect 97908 244326 97960 244332
rect 97816 243432 97868 243438
rect 97816 243374 97868 243380
rect 97828 196897 97856 243374
rect 97814 196888 97870 196897
rect 97814 196823 97870 196832
rect 97920 195945 97948 244326
rect 98656 241466 98684 443090
rect 220096 346390 220124 443158
rect 220084 346384 220136 346390
rect 220084 346326 220136 346332
rect 221476 306338 221504 443294
rect 221464 306332 221516 306338
rect 221464 306274 221516 306280
rect 224236 267714 224264 444926
rect 225604 443420 225656 443426
rect 225604 443362 225656 443368
rect 224960 309120 225012 309126
rect 224960 309062 225012 309068
rect 224972 308718 225000 309062
rect 224960 308712 225012 308718
rect 224960 308654 225012 308660
rect 224224 267708 224276 267714
rect 224224 267650 224276 267656
rect 99288 267028 99340 267034
rect 99288 266970 99340 266976
rect 98644 241460 98696 241466
rect 98644 241402 98696 241408
rect 97906 195936 97962 195945
rect 97906 195871 97962 195880
rect 97906 193760 97962 193769
rect 97906 193695 97962 193704
rect 97814 192808 97870 192817
rect 97814 192743 97870 192752
rect 97722 191040 97778 191049
rect 97722 190975 97778 190984
rect 97630 189952 97686 189961
rect 97630 189887 97686 189896
rect 97538 188184 97594 188193
rect 97538 188119 97594 188128
rect 97446 169960 97502 169969
rect 97446 169895 97502 169904
rect 97354 168328 97410 168337
rect 97354 168263 97410 168272
rect 97368 159662 97396 168263
rect 97356 159656 97408 159662
rect 97356 159598 97408 159604
rect 97460 159594 97488 169895
rect 97552 159866 97580 188119
rect 97540 159860 97592 159866
rect 97540 159802 97592 159808
rect 97448 159588 97500 159594
rect 97448 159530 97500 159536
rect 97644 157690 97672 189887
rect 97736 159798 97764 190975
rect 97724 159792 97776 159798
rect 97724 159734 97776 159740
rect 97828 159730 97856 192743
rect 97920 159934 97948 193695
rect 99300 168065 99328 266970
rect 225616 255270 225644 443362
rect 225708 320142 225736 445062
rect 226984 443488 227036 443494
rect 226984 443430 227036 443436
rect 226996 411262 227024 443430
rect 226984 411256 227036 411262
rect 226984 411198 227036 411204
rect 225696 320136 225748 320142
rect 225696 320078 225748 320084
rect 225604 255264 225656 255270
rect 225604 255206 225656 255212
rect 228376 247722 228404 445810
rect 228548 445256 228600 445262
rect 228548 445198 228600 445204
rect 228456 444916 228508 444922
rect 228456 444858 228508 444864
rect 228468 293962 228496 444858
rect 228560 372570 228588 445198
rect 228640 443284 228692 443290
rect 228640 443226 228692 443232
rect 228652 398818 228680 443226
rect 229756 440910 229784 445878
rect 229848 442270 229876 445946
rect 230400 443292 230428 446422
rect 230676 443306 230704 460906
rect 231872 447030 231900 476274
rect 231952 453348 232004 453354
rect 231952 453290 232004 453296
rect 231860 447024 231912 447030
rect 231860 446966 231912 446972
rect 231964 443306 231992 453290
rect 232412 447024 232464 447030
rect 232412 446966 232464 446972
rect 230676 443278 231150 443306
rect 231886 443278 231992 443306
rect 232424 443306 232452 446966
rect 233252 443306 233280 476682
rect 233332 476536 233384 476542
rect 233332 476478 233384 476484
rect 233344 460934 233372 476478
rect 237472 476468 237524 476474
rect 237472 476410 237524 476416
rect 235998 476368 236054 476377
rect 235998 476303 236000 476312
rect 236052 476303 236054 476312
rect 236184 476332 236236 476338
rect 236000 476274 236052 476280
rect 236184 476274 236236 476280
rect 236092 476264 236144 476270
rect 235998 476232 236054 476241
rect 234620 476196 234672 476202
rect 236092 476206 236144 476212
rect 235998 476167 236054 476176
rect 234620 476138 234672 476144
rect 233344 460906 233832 460934
rect 233804 443306 233832 460906
rect 234632 443306 234660 476138
rect 236012 476134 236040 476167
rect 234712 476128 234764 476134
rect 234712 476070 234764 476076
rect 236000 476128 236052 476134
rect 236000 476070 236052 476076
rect 234724 460934 234752 476070
rect 236000 475992 236052 475998
rect 236000 475934 236052 475940
rect 234724 460906 235304 460934
rect 235276 443306 235304 460906
rect 236012 447030 236040 475934
rect 236104 460934 236132 476206
rect 236196 476134 236224 476274
rect 237378 476232 237434 476241
rect 237378 476167 237380 476176
rect 237432 476167 237434 476176
rect 237380 476138 237432 476144
rect 236184 476128 236236 476134
rect 236184 476070 236236 476076
rect 237484 460934 237512 476410
rect 238680 476354 238708 476870
rect 242912 476746 242940 476983
rect 245752 476954 245804 476960
rect 247040 477012 247092 477018
rect 248418 476983 248474 476992
rect 247040 476954 247092 476960
rect 244646 476912 244702 476921
rect 244646 476847 244702 476856
rect 242900 476740 242952 476746
rect 242900 476682 242952 476688
rect 240140 476604 240192 476610
rect 240140 476546 240192 476552
rect 239126 476504 239182 476513
rect 239126 476439 239128 476448
rect 239180 476439 239182 476448
rect 239128 476410 239180 476416
rect 238680 476326 238800 476354
rect 236104 460906 236224 460934
rect 237484 460906 237696 460934
rect 236000 447024 236052 447030
rect 236000 446966 236052 446972
rect 236196 443306 236224 460906
rect 237012 447024 237064 447030
rect 237012 446966 237064 446972
rect 237024 443306 237052 446966
rect 237668 443306 237696 460906
rect 238772 443306 238800 476326
rect 238852 476264 238904 476270
rect 238852 476206 238904 476212
rect 238864 460934 238892 476206
rect 238864 460906 239352 460934
rect 239324 443306 239352 460906
rect 240152 443306 240180 476546
rect 244278 476504 244334 476513
rect 241428 476468 241480 476474
rect 244278 476439 244280 476448
rect 241428 476410 241480 476416
rect 244332 476439 244334 476448
rect 244280 476410 244332 476416
rect 240230 476232 240286 476241
rect 241440 476202 241468 476410
rect 242900 476332 242952 476338
rect 242900 476274 242952 476280
rect 242806 476232 242862 476241
rect 240230 476167 240286 476176
rect 241428 476196 241480 476202
rect 240244 460934 240272 476167
rect 241428 476138 241480 476144
rect 241520 476196 241572 476202
rect 242806 476167 242862 476176
rect 241520 476138 241572 476144
rect 240244 460906 240824 460934
rect 240796 443306 240824 460906
rect 241532 447030 241560 476138
rect 242820 476134 242848 476167
rect 242808 476128 242860 476134
rect 242808 476070 242860 476076
rect 241612 461644 241664 461650
rect 241612 461586 241664 461592
rect 241520 447024 241572 447030
rect 241520 446966 241572 446972
rect 241624 443306 241652 461586
rect 242912 460934 242940 476274
rect 244660 476270 244688 476847
rect 244648 476264 244700 476270
rect 244648 476206 244700 476212
rect 245658 476232 245714 476241
rect 245658 476167 245660 476176
rect 245712 476167 245714 476176
rect 245660 476138 245712 476144
rect 244280 476128 244332 476134
rect 244280 476070 244332 476076
rect 242912 460906 243216 460934
rect 242348 447024 242400 447030
rect 242348 446966 242400 446972
rect 242360 443306 242388 446966
rect 243188 443306 243216 460906
rect 243544 446072 243596 446078
rect 243544 446014 243596 446020
rect 243556 443698 243584 446014
rect 243544 443692 243596 443698
rect 243544 443634 243596 443640
rect 232424 443278 232714 443306
rect 233252 443278 233450 443306
rect 233804 443278 234278 443306
rect 234632 443278 235014 443306
rect 235276 443278 235750 443306
rect 236196 443278 236578 443306
rect 237024 443278 237314 443306
rect 237668 443278 238142 443306
rect 238772 443278 238878 443306
rect 239324 443278 239706 443306
rect 240152 443278 240442 443306
rect 240796 443278 241178 443306
rect 241624 443278 242006 443306
rect 242360 443278 242742 443306
rect 243188 443278 243570 443306
rect 244292 443292 244320 476070
rect 244648 451920 244700 451926
rect 244648 451862 244700 451868
rect 244660 443306 244688 451862
rect 245764 443306 245792 476954
rect 248432 476746 248460 476983
rect 247316 476740 247368 476746
rect 247316 476682 247368 476688
rect 248420 476740 248472 476746
rect 248420 476682 248472 476688
rect 247038 476640 247094 476649
rect 247038 476575 247094 476584
rect 247052 476542 247080 476575
rect 247040 476536 247092 476542
rect 247040 476478 247092 476484
rect 245844 476128 245896 476134
rect 245844 476070 245896 476076
rect 245856 460934 245884 476070
rect 247132 475380 247184 475386
rect 247132 475322 247184 475328
rect 245856 460906 246160 460934
rect 246132 443306 246160 460906
rect 247144 443306 247172 475322
rect 247328 460934 247356 476682
rect 248524 476626 248552 478178
rect 249890 477456 249946 477465
rect 249890 477391 249946 477400
rect 252466 477456 252522 477465
rect 252466 477391 252522 477400
rect 253846 477456 253902 477465
rect 253846 477391 253902 477400
rect 248432 476598 248552 476626
rect 247328 460906 247816 460934
rect 247788 443306 247816 460906
rect 248432 447030 248460 476598
rect 248512 476536 248564 476542
rect 248512 476478 248564 476484
rect 249798 476504 249854 476513
rect 248420 447024 248472 447030
rect 248420 446966 248472 446972
rect 248524 443306 248552 476478
rect 249798 476439 249854 476448
rect 249812 476406 249840 476439
rect 249800 476400 249852 476406
rect 249800 476342 249852 476348
rect 249904 460934 249932 477391
rect 251272 476400 251324 476406
rect 251272 476342 251324 476348
rect 250444 474088 250496 474094
rect 250444 474030 250496 474036
rect 249904 460906 250024 460934
rect 249340 447024 249392 447030
rect 249340 446966 249392 446972
rect 249352 443306 249380 446966
rect 249996 443306 250024 460906
rect 250456 447030 250484 474030
rect 250444 447024 250496 447030
rect 250444 446966 250496 446972
rect 244660 443278 245042 443306
rect 245764 443278 245870 443306
rect 246132 443278 246606 443306
rect 247144 443278 247434 443306
rect 247788 443278 248170 443306
rect 248524 443278 248998 443306
rect 249352 443278 249734 443306
rect 249996 443278 250470 443306
rect 251284 443292 251312 476342
rect 252374 476232 252430 476241
rect 252374 476167 252376 476176
rect 252428 476167 252430 476176
rect 252376 476138 252428 476144
rect 252008 447024 252060 447030
rect 252008 446966 252060 446972
rect 252020 443292 252048 446966
rect 252480 445754 252508 477391
rect 252558 476640 252614 476649
rect 252558 476575 252560 476584
rect 252612 476575 252614 476584
rect 252652 476604 252704 476610
rect 252560 476546 252612 476552
rect 252652 476546 252704 476552
rect 252664 460934 252692 476546
rect 252664 460906 253152 460934
rect 252480 445726 252600 445754
rect 252572 443306 252600 445726
rect 253124 443306 253152 460906
rect 253860 446282 253888 477391
rect 268014 477320 268070 477329
rect 268014 477255 268070 477264
rect 255410 477048 255466 477057
rect 255410 476983 255466 476992
rect 258078 477048 258134 477057
rect 258078 476983 258080 476992
rect 255320 476468 255372 476474
rect 255320 476410 255372 476416
rect 253940 476196 253992 476202
rect 253940 476138 253992 476144
rect 253952 447030 253980 476138
rect 254032 472728 254084 472734
rect 254032 472670 254084 472676
rect 253940 447024 253992 447030
rect 253940 446966 253992 446972
rect 253848 446276 253900 446282
rect 253848 446218 253900 446224
rect 254044 443306 254072 472670
rect 255332 460934 255360 476410
rect 255424 476270 255452 476983
rect 258132 476983 258134 476992
rect 262220 477012 262272 477018
rect 258080 476954 258132 476960
rect 262220 476954 262272 476960
rect 258078 476776 258134 476785
rect 258078 476711 258080 476720
rect 258132 476711 258134 476720
rect 258262 476776 258318 476785
rect 258262 476711 258318 476720
rect 258724 476740 258776 476746
rect 258080 476682 258132 476688
rect 255962 476368 256018 476377
rect 255962 476303 256018 476312
rect 256792 476332 256844 476338
rect 255412 476264 255464 476270
rect 255412 476206 255464 476212
rect 255332 460906 255544 460934
rect 254860 447024 254912 447030
rect 254860 446966 254912 446972
rect 254872 443306 254900 446966
rect 255516 443306 255544 460906
rect 255976 447098 256004 476303
rect 256792 476274 256844 476280
rect 256606 476232 256662 476241
rect 256606 476167 256662 476176
rect 255964 447092 256016 447098
rect 255964 447034 256016 447040
rect 256620 447030 256648 476167
rect 256804 460934 256832 476274
rect 258172 476264 258224 476270
rect 258172 476206 258224 476212
rect 258184 460934 258212 476206
rect 258276 476134 258304 476711
rect 258724 476682 258776 476688
rect 258264 476128 258316 476134
rect 258264 476070 258316 476076
rect 256804 460906 257016 460934
rect 258184 460906 258672 460934
rect 256608 447024 256660 447030
rect 256608 446966 256660 446972
rect 256700 446276 256752 446282
rect 256700 446218 256752 446224
rect 252572 443278 252862 443306
rect 253124 443278 253598 443306
rect 254044 443278 254426 443306
rect 254872 443278 255162 443306
rect 255516 443278 255898 443306
rect 256712 443292 256740 446218
rect 256988 443306 257016 460906
rect 258264 447092 258316 447098
rect 258264 447034 258316 447040
rect 256988 443278 257462 443306
rect 258276 443292 258304 447034
rect 258644 443306 258672 460906
rect 258736 446282 258764 476682
rect 260838 476640 260894 476649
rect 260838 476575 260894 476584
rect 260852 476542 260880 476575
rect 260840 476536 260892 476542
rect 260840 476478 260892 476484
rect 260932 476536 260984 476542
rect 260932 476478 260984 476484
rect 260746 476232 260802 476241
rect 259552 476196 259604 476202
rect 260746 476167 260802 476176
rect 259552 476138 259604 476144
rect 259564 460934 259592 476138
rect 259564 460906 260144 460934
rect 259736 447024 259788 447030
rect 259736 446966 259788 446972
rect 258724 446276 258776 446282
rect 258724 446218 258776 446224
rect 258644 443278 259026 443306
rect 259748 443292 259776 446966
rect 260116 443306 260144 460906
rect 260760 446622 260788 476167
rect 260944 460934 260972 476478
rect 261482 476368 261538 476377
rect 261482 476303 261538 476312
rect 260944 460906 261432 460934
rect 260748 446616 260800 446622
rect 260748 446558 260800 446564
rect 261404 446434 261432 460906
rect 261496 447030 261524 476303
rect 262232 460934 262260 476954
rect 263598 476640 263654 476649
rect 263598 476575 263654 476584
rect 264978 476640 265034 476649
rect 264978 476575 264980 476584
rect 263612 476406 263640 476575
rect 265032 476575 265034 476584
rect 264980 476546 265032 476552
rect 264242 476504 264298 476513
rect 268028 476474 268056 477255
rect 270498 477048 270554 477057
rect 270498 476983 270554 476992
rect 304998 477048 305054 477057
rect 304998 476983 305054 476992
rect 307758 477048 307814 477057
rect 307758 476983 307814 476992
rect 264242 476439 264298 476448
rect 268016 476468 268068 476474
rect 263600 476400 263652 476406
rect 263600 476342 263652 476348
rect 262862 476232 262918 476241
rect 262862 476167 262918 476176
rect 262232 460906 262536 460934
rect 261484 447024 261536 447030
rect 261484 446966 261536 446972
rect 261404 446406 261800 446434
rect 261300 446276 261352 446282
rect 261300 446218 261352 446224
rect 260116 443278 260590 443306
rect 261312 443292 261340 446218
rect 261772 443306 261800 446406
rect 262508 443306 262536 460906
rect 262876 447098 262904 476167
rect 263692 461644 263744 461650
rect 263692 461586 263744 461592
rect 262864 447092 262916 447098
rect 262864 447034 262916 447040
rect 261772 443278 262154 443306
rect 262508 443278 262890 443306
rect 263704 443292 263732 461586
rect 264256 446962 264284 476439
rect 268016 476410 268068 476416
rect 265622 476368 265678 476377
rect 265622 476303 265678 476312
rect 267554 476368 267610 476377
rect 270512 476338 270540 476983
rect 302238 476912 302294 476921
rect 302238 476847 302294 476856
rect 291200 476740 291252 476746
rect 291200 476682 291252 476688
rect 278780 476672 278832 476678
rect 277950 476640 278006 476649
rect 278780 476614 278832 476620
rect 277950 476575 278006 476584
rect 277964 476542 277992 476575
rect 277952 476536 278004 476542
rect 273258 476504 273314 476513
rect 277952 476478 278004 476484
rect 273258 476439 273314 476448
rect 267554 476303 267610 476312
rect 270500 476332 270552 476338
rect 265164 450628 265216 450634
rect 265164 450570 265216 450576
rect 264244 446956 264296 446962
rect 264244 446898 264296 446904
rect 264428 446616 264480 446622
rect 264428 446558 264480 446564
rect 264440 443292 264468 446558
rect 265176 443292 265204 450570
rect 265636 446486 265664 476303
rect 266266 476232 266322 476241
rect 266266 476167 266322 476176
rect 266280 451926 266308 476167
rect 267568 475386 267596 476303
rect 270500 476274 270552 476280
rect 273272 476270 273300 476439
rect 274454 476368 274510 476377
rect 274454 476303 274510 476312
rect 276018 476368 276074 476377
rect 276018 476303 276074 476312
rect 273260 476264 273312 476270
rect 267646 476232 267702 476241
rect 267646 476167 267702 476176
rect 269026 476232 269082 476241
rect 269026 476167 269082 476176
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 271786 476232 271842 476241
rect 271786 476167 271842 476176
rect 273166 476232 273222 476241
rect 273260 476206 273312 476212
rect 273166 476167 273222 476176
rect 267556 475380 267608 475386
rect 267556 475322 267608 475328
rect 266452 468580 266504 468586
rect 266452 468522 266504 468528
rect 266268 451920 266320 451926
rect 266268 451862 266320 451868
rect 265992 447024 266044 447030
rect 265992 446966 266044 446972
rect 265624 446480 265676 446486
rect 265624 446422 265676 446428
rect 266004 443292 266032 446966
rect 266464 443306 266492 468522
rect 267660 453354 267688 476167
rect 267740 469940 267792 469946
rect 267740 469882 267792 469888
rect 267752 460934 267780 469882
rect 267752 460906 267872 460934
rect 267648 453348 267700 453354
rect 267648 453290 267700 453296
rect 267556 447092 267608 447098
rect 267556 447034 267608 447040
rect 266464 443278 266754 443306
rect 267568 443292 267596 447034
rect 267844 443306 267872 460906
rect 269040 455394 269068 476167
rect 269212 472728 269264 472734
rect 269212 472670 269264 472676
rect 269224 460934 269252 472670
rect 269224 460906 269528 460934
rect 269028 455388 269080 455394
rect 269028 455330 269080 455336
rect 269120 446956 269172 446962
rect 269120 446898 269172 446904
rect 267844 443278 268318 443306
rect 269132 443292 269160 446898
rect 269500 443306 269528 460906
rect 270420 451994 270448 476167
rect 270960 456136 271012 456142
rect 270960 456078 271012 456084
rect 270408 451988 270460 451994
rect 270408 451930 270460 451936
rect 270592 446480 270644 446486
rect 270592 446422 270644 446428
rect 269500 443278 269882 443306
rect 270604 443292 270632 446422
rect 270972 443306 271000 456078
rect 271800 452810 271828 476167
rect 271880 463004 271932 463010
rect 271880 462946 271932 462952
rect 271788 452804 271840 452810
rect 271788 452746 271840 452752
rect 271892 447030 271920 462946
rect 273180 461786 273208 476167
rect 273168 461780 273220 461786
rect 273168 461722 273220 461728
rect 274468 454782 274496 476303
rect 274546 476232 274602 476241
rect 274546 476167 274602 476176
rect 275926 476232 275982 476241
rect 276032 476202 276060 476303
rect 277306 476232 277362 476241
rect 275926 476167 275982 476176
rect 276020 476196 276072 476202
rect 274456 454776 274508 454782
rect 274456 454718 274508 454724
rect 274088 453416 274140 453422
rect 274088 453358 274140 453364
rect 273260 453348 273312 453354
rect 273260 453290 273312 453296
rect 271972 451920 272024 451926
rect 271972 451862 272024 451868
rect 271880 447024 271932 447030
rect 271880 446966 271932 446972
rect 271984 443306 272012 451862
rect 272708 447024 272760 447030
rect 272708 446966 272760 446972
rect 272720 443306 272748 446966
rect 273272 443306 273300 453290
rect 274100 443306 274128 453358
rect 274560 451926 274588 476167
rect 274640 475380 274692 475386
rect 274640 475322 274692 475328
rect 274652 460934 274680 475322
rect 274652 460906 274864 460934
rect 274548 451920 274600 451926
rect 274548 451862 274600 451868
rect 274836 443306 274864 460906
rect 275940 453354 275968 476167
rect 277306 476167 277362 476176
rect 278686 476232 278742 476241
rect 278686 476167 278742 476176
rect 276020 476138 276072 476144
rect 276020 474088 276072 474094
rect 276020 474030 276072 474036
rect 275928 453348 275980 453354
rect 275928 453290 275980 453296
rect 270972 443278 271446 443306
rect 271984 443278 272182 443306
rect 272720 443278 273010 443306
rect 273272 443278 273746 443306
rect 274100 443278 274482 443306
rect 274836 443278 275310 443306
rect 276032 443292 276060 474030
rect 277320 461718 277348 476167
rect 277584 476128 277636 476134
rect 277584 476070 277636 476076
rect 277308 461712 277360 461718
rect 277308 461654 277360 461660
rect 276480 455388 276532 455394
rect 276480 455330 276532 455336
rect 276492 443306 276520 455330
rect 277492 451988 277544 451994
rect 277492 451930 277544 451936
rect 277504 447030 277532 451930
rect 277492 447024 277544 447030
rect 277492 446966 277544 446972
rect 276492 443278 276874 443306
rect 277596 443292 277624 476070
rect 278700 454714 278728 476167
rect 278688 454708 278740 454714
rect 278688 454650 278740 454656
rect 278044 447024 278096 447030
rect 278044 446966 278096 446972
rect 278056 443306 278084 446966
rect 278792 443306 278820 476614
rect 280160 476604 280212 476610
rect 280160 476546 280212 476552
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 279424 452804 279476 452810
rect 279424 452746 279476 452752
rect 279436 443306 279464 452746
rect 280080 451994 280108 476167
rect 280172 460934 280200 476546
rect 281540 476536 281592 476542
rect 281540 476478 281592 476484
rect 280250 476232 280306 476241
rect 280250 476167 280306 476176
rect 280264 461650 280292 476167
rect 280344 461780 280396 461786
rect 280344 461722 280396 461728
rect 280252 461644 280304 461650
rect 280252 461586 280304 461592
rect 280356 460934 280384 461722
rect 281552 460934 281580 476478
rect 282920 476468 282972 476474
rect 282920 476410 282972 476416
rect 280172 460906 280292 460934
rect 280356 460906 281120 460934
rect 281552 460906 281856 460934
rect 280068 451988 280120 451994
rect 280068 451930 280120 451936
rect 280264 445754 280292 460906
rect 280264 445726 280384 445754
rect 280356 443306 280384 445726
rect 281092 443306 281120 460906
rect 281828 443306 281856 460906
rect 282932 447030 282960 476410
rect 284300 476400 284352 476406
rect 284300 476342 284352 476348
rect 283102 476232 283158 476241
rect 283102 476167 283158 476176
rect 283012 454776 283064 454782
rect 283012 454718 283064 454724
rect 282920 447024 282972 447030
rect 282920 446966 282972 446972
rect 278056 443278 278438 443306
rect 278792 443278 279174 443306
rect 279436 443278 279910 443306
rect 280356 443278 280738 443306
rect 281092 443278 281474 443306
rect 281828 443278 282302 443306
rect 283024 443292 283052 454718
rect 283116 450634 283144 476167
rect 283104 450628 283156 450634
rect 283104 450570 283156 450576
rect 284312 447030 284340 476342
rect 285680 476332 285732 476338
rect 285680 476274 285732 476280
rect 284392 451920 284444 451926
rect 284392 451862 284444 451868
rect 283380 447024 283432 447030
rect 283380 446966 283432 446972
rect 284300 447024 284352 447030
rect 284300 446966 284352 446972
rect 283392 443306 283420 446966
rect 284404 443306 284432 451862
rect 285692 447030 285720 476274
rect 288440 476264 288492 476270
rect 285770 476232 285826 476241
rect 285770 476167 285826 476176
rect 287058 476232 287114 476241
rect 288440 476206 288492 476212
rect 289910 476232 289966 476241
rect 287058 476167 287114 476176
rect 285784 468586 285812 476167
rect 287072 469946 287100 476167
rect 287060 469940 287112 469946
rect 287060 469882 287112 469888
rect 285772 468580 285824 468586
rect 285772 468522 285824 468528
rect 287060 461712 287112 461718
rect 287060 461654 287112 461660
rect 287072 460934 287100 461654
rect 287072 460906 287376 460934
rect 285772 453348 285824 453354
rect 285772 453290 285824 453296
rect 285036 447024 285088 447030
rect 285036 446966 285088 446972
rect 285680 447024 285732 447030
rect 285680 446966 285732 446972
rect 285048 443306 285076 446966
rect 285784 443306 285812 453290
rect 286508 447024 286560 447030
rect 286508 446966 286560 446972
rect 286520 443306 286548 446966
rect 287348 443306 287376 460906
rect 283392 443278 283774 443306
rect 284404 443278 284602 443306
rect 285048 443278 285338 443306
rect 285784 443278 286166 443306
rect 286520 443278 286902 443306
rect 287348 443278 287730 443306
rect 288452 443292 288480 476206
rect 289820 476196 289872 476202
rect 289910 476167 289966 476176
rect 289820 476138 289872 476144
rect 288808 454708 288860 454714
rect 288808 454650 288860 454656
rect 288820 443306 288848 454650
rect 289832 443306 289860 476138
rect 289924 472734 289952 476167
rect 289912 472728 289964 472734
rect 289912 472670 289964 472676
rect 290280 451988 290332 451994
rect 290280 451930 290332 451936
rect 290292 443306 290320 451930
rect 291212 443306 291240 476682
rect 292578 476232 292634 476241
rect 292578 476167 292634 476176
rect 295430 476232 295486 476241
rect 295430 476167 295486 476176
rect 298190 476232 298246 476241
rect 298190 476167 298246 476176
rect 300858 476232 300914 476241
rect 300858 476167 300914 476176
rect 292592 456142 292620 476167
rect 295340 467220 295392 467226
rect 295340 467162 295392 467168
rect 295352 460934 295380 467162
rect 295444 463010 295472 476167
rect 298100 471368 298152 471374
rect 298100 471310 298152 471316
rect 295432 463004 295484 463010
rect 295432 462946 295484 462952
rect 295352 460906 295840 460934
rect 292580 456136 292632 456142
rect 292580 456078 292632 456084
rect 294144 451920 294196 451926
rect 294144 451862 294196 451868
rect 293132 446208 293184 446214
rect 293132 446150 293184 446156
rect 292304 446140 292356 446146
rect 292304 446082 292356 446088
rect 288820 443278 289202 443306
rect 289832 443278 290030 443306
rect 290292 443278 290766 443306
rect 291212 443278 291594 443306
rect 292316 443292 292344 446082
rect 293144 443292 293172 446150
rect 293868 445800 293920 445806
rect 293868 445742 293920 445748
rect 293880 443292 293908 445742
rect 294156 443306 294184 451862
rect 295432 444780 295484 444786
rect 295432 444722 295484 444728
rect 294156 443278 294630 443306
rect 295444 443292 295472 444722
rect 295812 443306 295840 460906
rect 296720 453348 296772 453354
rect 296720 453290 296772 453296
rect 296732 443306 296760 453290
rect 298112 443306 298140 471310
rect 298204 453422 298232 476167
rect 300872 474094 300900 476167
rect 302252 476134 302280 476847
rect 305012 476678 305040 476983
rect 305000 476672 305052 476678
rect 305000 476614 305052 476620
rect 307772 476610 307800 476983
rect 307760 476604 307812 476610
rect 307760 476546 307812 476552
rect 302240 476128 302292 476134
rect 302240 476070 302292 476076
rect 301044 475380 301096 475386
rect 301044 475322 301096 475328
rect 300860 474088 300912 474094
rect 300860 474030 300912 474036
rect 300952 456136 301004 456142
rect 300952 456078 301004 456084
rect 298928 454708 298980 454714
rect 298928 454650 298980 454656
rect 298192 453416 298244 453422
rect 298192 453358 298244 453364
rect 298940 443306 298968 454650
rect 300964 447030 300992 456078
rect 300952 447024 301004 447030
rect 300952 446966 301004 446972
rect 300032 444848 300084 444854
rect 300032 444790 300084 444796
rect 295812 443278 296194 443306
rect 296732 443278 297022 443306
rect 298112 443278 298494 443306
rect 298940 443278 299322 443306
rect 300044 443292 300072 444790
rect 301056 443306 301084 475322
rect 305000 464432 305052 464438
rect 305000 464374 305052 464380
rect 305012 460934 305040 464374
rect 309152 460934 309180 478178
rect 314752 478168 314804 478174
rect 314752 478110 314804 478116
rect 310518 476912 310574 476921
rect 310518 476847 310574 476856
rect 310532 476542 310560 476847
rect 310520 476536 310572 476542
rect 310520 476478 310572 476484
rect 313278 476504 313334 476513
rect 313278 476439 313280 476448
rect 313332 476439 313334 476448
rect 314658 476504 314714 476513
rect 314658 476439 314714 476448
rect 313280 476410 313332 476416
rect 314672 476406 314700 476439
rect 314660 476400 314712 476406
rect 314660 476342 314712 476348
rect 314764 470594 314792 478110
rect 322938 476912 322994 476921
rect 322938 476847 322994 476856
rect 325790 476912 325846 476921
rect 325790 476847 325846 476856
rect 317418 476368 317474 476377
rect 317418 476303 317420 476312
rect 317472 476303 317474 476312
rect 320178 476368 320234 476377
rect 320178 476303 320234 476312
rect 317420 476274 317472 476280
rect 320192 476270 320220 476303
rect 320180 476264 320232 476270
rect 320180 476206 320232 476212
rect 322952 476202 322980 476847
rect 325804 476746 325832 476847
rect 325792 476740 325844 476746
rect 325792 476682 325844 476688
rect 322940 476196 322992 476202
rect 322940 476138 322992 476144
rect 331220 474768 331272 474774
rect 331220 474710 331272 474716
rect 320180 474088 320232 474094
rect 320180 474030 320232 474036
rect 314672 470566 314792 470594
rect 305012 460906 305960 460934
rect 309152 460906 309824 460934
rect 303620 457564 303672 457570
rect 303620 457506 303672 457512
rect 303160 449404 303212 449410
rect 303160 449346 303212 449352
rect 301228 447024 301280 447030
rect 301228 446966 301280 446972
rect 300886 443278 301084 443306
rect 301240 443306 301268 446966
rect 302424 446616 302476 446622
rect 302424 446558 302476 446564
rect 301240 443278 301622 443306
rect 302436 443292 302464 446558
rect 303172 443292 303200 449346
rect 303632 443306 303660 457506
rect 305460 449540 305512 449546
rect 305460 449482 305512 449488
rect 304724 446276 304776 446282
rect 304724 446218 304776 446224
rect 303632 443278 303922 443306
rect 304736 443292 304764 446218
rect 305472 443292 305500 449482
rect 305932 443306 305960 460906
rect 308128 458924 308180 458930
rect 308128 458866 308180 458872
rect 307852 449676 307904 449682
rect 307852 449618 307904 449624
rect 307024 446344 307076 446350
rect 307024 446286 307076 446292
rect 305932 443278 306314 443306
rect 307036 443292 307064 446286
rect 307864 443292 307892 449618
rect 308140 443306 308168 458866
rect 309324 443692 309376 443698
rect 309324 443634 309376 443640
rect 308140 443278 308614 443306
rect 309336 443292 309364 443634
rect 309796 443306 309824 460906
rect 313188 446684 313240 446690
rect 313188 446626 313240 446632
rect 312452 446548 312504 446554
rect 312452 446490 312504 446496
rect 310888 446480 310940 446486
rect 310888 446422 310940 446428
rect 309796 443278 310178 443306
rect 310900 443292 310928 446422
rect 311716 446412 311768 446418
rect 311716 446354 311768 446360
rect 311728 443292 311756 446354
rect 312464 443292 312492 446490
rect 313200 443292 313228 446626
rect 314016 444440 314068 444446
rect 314016 444382 314068 444388
rect 314028 443292 314056 444382
rect 314672 443306 314700 470566
rect 314752 465724 314804 465730
rect 314752 465666 314804 465672
rect 314764 460934 314792 465666
rect 317420 461644 317472 461650
rect 317420 461586 317472 461592
rect 317432 460934 317460 461586
rect 320192 460934 320220 474030
rect 328460 471300 328512 471306
rect 328460 471242 328512 471248
rect 327080 469872 327132 469878
rect 327080 469814 327132 469820
rect 324320 468512 324372 468518
rect 324320 468454 324372 468460
rect 321560 467152 321612 467158
rect 321560 467094 321612 467100
rect 321572 460934 321600 467094
rect 324332 460934 324360 468454
rect 314764 460906 315160 460934
rect 317432 460906 318288 460934
rect 320192 460906 320680 460934
rect 321572 460906 322152 460934
rect 324332 460906 324544 460934
rect 315132 443306 315160 460906
rect 317144 449608 317196 449614
rect 317144 449550 317196 449556
rect 316316 443624 316368 443630
rect 316316 443566 316368 443572
rect 314672 443278 314778 443306
rect 315132 443278 315606 443306
rect 316328 443292 316356 443566
rect 317156 443292 317184 449550
rect 317880 447976 317932 447982
rect 317880 447918 317932 447924
rect 317892 443292 317920 447918
rect 318260 443306 318288 460906
rect 319444 449472 319496 449478
rect 319444 449414 319496 449420
rect 318260 443278 318642 443306
rect 319456 443292 319484 449414
rect 320180 447908 320232 447914
rect 320180 447850 320232 447856
rect 320192 443292 320220 447850
rect 320652 443306 320680 460906
rect 321744 449336 321796 449342
rect 321744 449278 321796 449284
rect 320652 443278 321034 443306
rect 321756 443292 321784 449278
rect 322124 443306 322152 460906
rect 322940 460284 322992 460290
rect 322940 460226 322992 460232
rect 322952 443306 322980 460226
rect 323584 456068 323636 456074
rect 323584 456010 323636 456016
rect 323596 443306 323624 456010
rect 324516 443306 324544 460906
rect 325608 450628 325660 450634
rect 325608 450570 325660 450576
rect 322124 443278 322506 443306
rect 322952 443278 323334 443306
rect 323596 443278 324070 443306
rect 324516 443278 324898 443306
rect 325620 443292 325648 450570
rect 326436 449268 326488 449274
rect 326436 449210 326488 449216
rect 326448 443292 326476 449210
rect 327092 443306 327120 469814
rect 327172 465724 327224 465730
rect 327172 465666 327224 465672
rect 327184 460934 327212 465666
rect 328472 460934 328500 471242
rect 329840 468512 329892 468518
rect 329840 468454 329892 468460
rect 327184 460906 327488 460934
rect 328472 460906 329144 460934
rect 327460 443306 327488 460906
rect 328736 449200 328788 449206
rect 328736 449142 328788 449148
rect 327092 443278 327198 443306
rect 327460 443278 327934 443306
rect 328748 443292 328776 449142
rect 329116 443306 329144 460906
rect 329852 443306 329880 468454
rect 331232 460934 331260 474710
rect 347872 474020 347924 474026
rect 347872 473962 347924 473968
rect 346492 472660 346544 472666
rect 346492 472602 346544 472608
rect 334072 469872 334124 469878
rect 334072 469814 334124 469820
rect 332600 463004 332652 463010
rect 332600 462946 332652 462952
rect 331232 460906 331536 460934
rect 331036 450560 331088 450566
rect 331036 450502 331088 450508
rect 329116 443278 329498 443306
rect 329852 443278 330326 443306
rect 331048 443292 331076 450502
rect 331508 443306 331536 460906
rect 331508 443278 331890 443306
rect 332612 443292 332640 462946
rect 332692 462392 332744 462398
rect 332692 462334 332744 462340
rect 332704 460934 332732 462334
rect 334084 460934 334112 469814
rect 332704 460906 333008 460934
rect 334084 460906 334480 460934
rect 332980 443306 333008 460906
rect 333980 446616 334032 446622
rect 333980 446558 334032 446564
rect 333992 445058 334020 446558
rect 334164 445188 334216 445194
rect 334164 445130 334216 445136
rect 333980 445052 334032 445058
rect 333980 444994 334032 445000
rect 332980 443278 333362 443306
rect 334176 443292 334204 445130
rect 334452 443306 334480 460906
rect 341892 448112 341944 448118
rect 341892 448054 341944 448060
rect 339592 446684 339644 446690
rect 339592 446626 339644 446632
rect 337200 446616 337252 446622
rect 337200 446558 337252 446564
rect 336464 445256 336516 445262
rect 336464 445198 336516 445204
rect 335544 443488 335596 443494
rect 335544 443430 335596 443436
rect 335556 443306 335584 443430
rect 334452 443278 334926 443306
rect 335556 443278 335754 443306
rect 336476 443292 336504 445198
rect 337212 443292 337240 446558
rect 338028 446004 338080 446010
rect 338028 445946 338080 445952
rect 338040 443292 338068 445946
rect 338764 445120 338816 445126
rect 338764 445062 338816 445068
rect 338776 443292 338804 445062
rect 339604 443292 339632 446626
rect 341156 444984 341208 444990
rect 341156 444926 341208 444932
rect 340052 443352 340104 443358
rect 340104 443300 340354 443306
rect 340052 443294 340354 443300
rect 340064 443278 340354 443294
rect 341168 443292 341196 444926
rect 341904 443292 341932 448054
rect 344192 448044 344244 448050
rect 344192 447986 344244 447992
rect 343456 444712 343508 444718
rect 343456 444654 343508 444660
rect 342260 443420 342312 443426
rect 342260 443362 342312 443368
rect 342272 443306 342300 443362
rect 342272 443278 342654 443306
rect 343468 443292 343496 444654
rect 344204 443292 344232 447986
rect 345020 446072 345072 446078
rect 345020 446014 345072 446020
rect 345032 443292 345060 446014
rect 345756 444644 345808 444650
rect 345756 444586 345808 444592
rect 345768 443292 345796 444586
rect 346504 443306 346532 472602
rect 347884 460934 347912 473962
rect 351920 464364 351972 464370
rect 351920 464306 351972 464312
rect 347884 460906 348464 460934
rect 347320 445936 347372 445942
rect 347320 445878 347372 445884
rect 346504 443278 346610 443306
rect 347332 443292 347360 445878
rect 348056 444576 348108 444582
rect 348056 444518 348108 444524
rect 348068 443292 348096 444518
rect 348436 443306 348464 460906
rect 350080 460216 350132 460222
rect 350080 460158 350132 460164
rect 349620 445868 349672 445874
rect 349620 445810 349672 445816
rect 348436 443278 348910 443306
rect 349632 443292 349660 445810
rect 350092 443306 350120 460158
rect 350816 458856 350868 458862
rect 350816 458798 350868 458804
rect 350828 443306 350856 458798
rect 350092 443278 350474 443306
rect 350828 443278 351210 443306
rect 351932 443292 351960 464306
rect 352288 457496 352340 457502
rect 352288 457438 352340 457444
rect 352300 443306 352328 457438
rect 353484 447840 353536 447846
rect 353484 447782 353536 447788
rect 352300 443278 352774 443306
rect 353496 443292 353524 447782
rect 357452 446690 357480 700266
rect 357440 446684 357492 446690
rect 357440 446626 357492 446632
rect 357544 446486 357572 700402
rect 357636 478242 357664 700538
rect 358820 700528 358872 700534
rect 358820 700470 358872 700476
rect 357624 478236 357676 478242
rect 357624 478178 357676 478184
rect 358832 446622 358860 700470
rect 358912 700392 358964 700398
rect 358912 700334 358964 700340
rect 358820 446616 358872 446622
rect 358820 446558 358872 446564
rect 358924 446554 358952 700334
rect 359464 700324 359516 700330
rect 359464 700266 359516 700272
rect 359476 469878 359504 700266
rect 360844 670744 360896 670750
rect 360844 670686 360896 670692
rect 359464 469872 359516 469878
rect 359464 469814 359516 469820
rect 360856 454714 360884 670686
rect 363604 590708 363656 590714
rect 363604 590650 363656 590656
rect 363616 460290 363644 590650
rect 363604 460284 363656 460290
rect 363604 460226 363656 460232
rect 364352 458930 364380 702406
rect 397472 700330 397500 703520
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 371884 696992 371936 696998
rect 371884 696934 371936 696940
rect 367744 643136 367796 643142
rect 367744 643078 367796 643084
rect 364340 458924 364392 458930
rect 364340 458866 364392 458872
rect 360844 454708 360896 454714
rect 360844 454650 360896 454656
rect 367756 450634 367784 643078
rect 369124 576904 369176 576910
rect 369124 576846 369176 576852
rect 369136 467226 369164 576846
rect 369124 467220 369176 467226
rect 369124 467162 369176 467168
rect 371896 465730 371924 696934
rect 373264 630692 373316 630698
rect 373264 630634 373316 630640
rect 373276 471374 373304 630634
rect 378784 616888 378836 616894
rect 378784 616830 378836 616836
rect 373264 471368 373316 471374
rect 373264 471310 373316 471316
rect 371884 465724 371936 465730
rect 371884 465666 371936 465672
rect 378796 453354 378824 616830
rect 381544 563100 381596 563106
rect 381544 563042 381596 563048
rect 378784 453348 378836 453354
rect 378784 453290 378836 453296
rect 381556 451926 381584 563042
rect 381544 451920 381596 451926
rect 381544 451862 381596 451868
rect 367744 450628 367796 450634
rect 367744 450570 367796 450576
rect 412652 449682 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 699718 429884 703520
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 464438 428504 699654
rect 428464 464432 428516 464438
rect 428464 464374 428516 464380
rect 462332 463010 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 467104 700324 467156 700330
rect 467104 700266 467156 700272
rect 467116 468518 467144 700266
rect 467104 468512 467156 468518
rect 467104 468454 467156 468460
rect 462320 463004 462372 463010
rect 462320 462946 462372 462952
rect 412640 449676 412692 449682
rect 412640 449618 412692 449624
rect 477512 449546 477540 702406
rect 480904 484424 480956 484430
rect 480904 484366 480956 484372
rect 480916 461650 480944 484366
rect 480904 461644 480956 461650
rect 480904 461586 480956 461592
rect 494072 457570 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 527824 700324 527876 700330
rect 527824 700266 527876 700272
rect 498844 536852 498896 536858
rect 498844 536794 498896 536800
rect 498856 474094 498884 536794
rect 498844 474088 498896 474094
rect 498844 474030 498896 474036
rect 494060 457564 494112 457570
rect 494060 457506 494112 457512
rect 527836 456142 527864 700266
rect 527824 456136 527876 456142
rect 527824 456078 527876 456084
rect 477500 449540 477552 449546
rect 477500 449482 477552 449488
rect 542372 449410 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 475386 580304 683839
rect 580264 475380 580316 475386
rect 580264 475322 580316 475328
rect 542360 449404 542412 449410
rect 542360 449346 542412 449352
rect 358912 446548 358964 446554
rect 358912 446490 358964 446496
rect 357532 446480 357584 446486
rect 357532 446422 357584 446428
rect 362224 446412 362276 446418
rect 362224 446354 362276 446360
rect 361028 446208 361080 446214
rect 361028 446150 361080 446156
rect 355876 444916 355928 444922
rect 355876 444858 355928 444864
rect 354048 443290 354338 443306
rect 355888 443292 355916 444858
rect 358176 444508 358228 444514
rect 358176 444450 358228 444456
rect 358188 443292 358216 444450
rect 354036 443284 354338 443290
rect 354088 443278 354338 443284
rect 354036 443226 354088 443232
rect 354772 443216 354824 443222
rect 354824 443164 355074 443170
rect 354772 443158 355074 443164
rect 354784 443142 355074 443158
rect 356256 443154 356638 443170
rect 356244 443148 356638 443154
rect 356296 443142 356638 443148
rect 356244 443090 356296 443096
rect 356980 443080 357032 443086
rect 298006 443048 298062 443057
rect 297758 443006 298006 443034
rect 357032 443028 357374 443034
rect 356980 443022 357374 443028
rect 356992 443006 357374 443022
rect 358832 443018 358938 443034
rect 358820 443012 358938 443018
rect 298006 442983 298062 442992
rect 358872 443006 358938 443012
rect 358820 442954 358872 442960
rect 359462 442776 359518 442785
rect 359518 442734 359766 442762
rect 360502 442734 360976 442762
rect 359462 442711 359518 442720
rect 229836 442264 229888 442270
rect 229836 442206 229888 442212
rect 229744 440904 229796 440910
rect 229744 440846 229796 440852
rect 228640 398812 228692 398818
rect 228640 398754 228692 398760
rect 228548 372564 228600 372570
rect 228548 372506 228600 372512
rect 230124 307086 230152 310420
rect 230112 307080 230164 307086
rect 230112 307022 230164 307028
rect 230308 296714 230336 310420
rect 230492 304298 230520 310420
rect 230664 306332 230716 306338
rect 230664 306274 230716 306280
rect 230480 304292 230532 304298
rect 230480 304234 230532 304240
rect 229204 296686 230336 296714
rect 228456 293956 228508 293962
rect 228456 293898 228508 293904
rect 229204 249082 229232 296686
rect 230676 273970 230704 306274
rect 230768 306270 230796 310420
rect 230952 306610 230980 310420
rect 230940 306604 230992 306610
rect 230940 306546 230992 306552
rect 231136 306490 231164 310420
rect 230860 306462 231164 306490
rect 230756 306264 230808 306270
rect 230756 306206 230808 306212
rect 230756 306128 230808 306134
rect 230756 306070 230808 306076
rect 230768 287706 230796 306070
rect 230756 287700 230808 287706
rect 230756 287642 230808 287648
rect 230664 273964 230716 273970
rect 230664 273906 230716 273912
rect 229192 249076 229244 249082
rect 229192 249018 229244 249024
rect 228364 247716 228416 247722
rect 228364 247658 228416 247664
rect 230860 246362 230888 306462
rect 230940 306400 230992 306406
rect 230940 306342 230992 306348
rect 230952 262886 230980 306342
rect 231032 306264 231084 306270
rect 231032 306206 231084 306212
rect 231044 298790 231072 306206
rect 231412 302938 231440 310420
rect 231596 306338 231624 310420
rect 231584 306332 231636 306338
rect 231584 306274 231636 306280
rect 231780 306134 231808 310420
rect 232056 308786 232084 310420
rect 232044 308780 232096 308786
rect 232044 308722 232096 308728
rect 232044 306400 232096 306406
rect 232044 306342 232096 306348
rect 231952 306332 232004 306338
rect 231952 306274 232004 306280
rect 231768 306128 231820 306134
rect 231768 306070 231820 306076
rect 231400 302932 231452 302938
rect 231400 302874 231452 302880
rect 231032 298784 231084 298790
rect 231032 298726 231084 298732
rect 230940 262880 230992 262886
rect 230940 262822 230992 262828
rect 231964 260166 231992 306274
rect 232056 283626 232084 306342
rect 232240 302234 232268 310420
rect 232148 302206 232268 302234
rect 232148 289134 232176 302206
rect 232424 296714 232452 310420
rect 232516 310406 232714 310434
rect 232516 306338 232544 310406
rect 232884 308922 232912 310420
rect 232976 310406 233174 310434
rect 232872 308916 232924 308922
rect 232872 308858 232924 308864
rect 232976 306406 233004 310406
rect 232964 306400 233016 306406
rect 232964 306342 233016 306348
rect 232504 306332 232556 306338
rect 232504 306274 232556 306280
rect 232240 296686 232452 296714
rect 232136 289128 232188 289134
rect 232136 289070 232188 289076
rect 232044 283620 232096 283626
rect 232044 283562 232096 283568
rect 231952 260160 232004 260166
rect 231952 260102 232004 260108
rect 232240 251870 232268 296686
rect 232228 251864 232280 251870
rect 232228 251806 232280 251812
rect 230848 246356 230900 246362
rect 230848 246298 230900 246304
rect 233344 244934 233372 310420
rect 233528 308650 233556 310420
rect 233804 308854 233832 310420
rect 233792 308848 233844 308854
rect 233792 308790 233844 308796
rect 233516 308644 233568 308650
rect 233516 308586 233568 308592
rect 233988 306354 234016 310420
rect 233436 306326 234016 306354
rect 233436 282198 233464 306326
rect 234172 305130 234200 310420
rect 234448 308310 234476 310420
rect 234632 308990 234660 310420
rect 234830 310406 234936 310434
rect 234620 308984 234672 308990
rect 234620 308926 234672 308932
rect 234712 308508 234764 308514
rect 234712 308450 234764 308456
rect 234436 308304 234488 308310
rect 234436 308246 234488 308252
rect 234252 308168 234304 308174
rect 234252 308110 234304 308116
rect 233528 305102 234200 305130
rect 233424 282192 233476 282198
rect 233424 282134 233476 282140
rect 233528 245002 233556 305102
rect 234264 302234 234292 308110
rect 233896 302206 234292 302234
rect 233896 282266 233924 302206
rect 233884 282260 233936 282266
rect 233884 282202 233936 282208
rect 234724 261526 234752 308450
rect 234804 308372 234856 308378
rect 234804 308314 234856 308320
rect 234816 279478 234844 308314
rect 234908 280838 234936 310406
rect 234988 308440 235040 308446
rect 234988 308382 235040 308388
rect 235000 291854 235028 308382
rect 234988 291848 235040 291854
rect 234988 291790 235040 291796
rect 234896 280832 234948 280838
rect 234896 280774 234948 280780
rect 234804 279472 234856 279478
rect 234804 279414 234856 279420
rect 234712 261520 234764 261526
rect 234712 261462 234764 261468
rect 235092 253230 235120 310420
rect 235276 308582 235304 310420
rect 235264 308576 235316 308582
rect 235264 308518 235316 308524
rect 235460 308378 235488 310420
rect 235552 310406 235750 310434
rect 235552 308446 235580 310406
rect 235920 308514 235948 310420
rect 235908 308508 235960 308514
rect 235908 308450 235960 308456
rect 235540 308440 235592 308446
rect 235540 308382 235592 308388
rect 236092 308440 236144 308446
rect 236092 308382 236144 308388
rect 235448 308372 235500 308378
rect 235448 308314 235500 308320
rect 236104 276690 236132 308382
rect 236196 278050 236224 310420
rect 236380 308394 236408 310420
rect 236564 308718 236592 310420
rect 236656 310406 236854 310434
rect 236552 308712 236604 308718
rect 236552 308654 236604 308660
rect 236656 308446 236684 310406
rect 236288 308366 236408 308394
rect 236644 308440 236696 308446
rect 236644 308382 236696 308388
rect 236288 284986 236316 308366
rect 237024 308258 237052 310420
rect 237208 309126 237236 310420
rect 237392 310406 237498 310434
rect 237196 309120 237248 309126
rect 237196 309062 237248 309068
rect 237104 308576 237156 308582
rect 237104 308518 237156 308524
rect 236380 308230 237052 308258
rect 236276 284980 236328 284986
rect 236276 284922 236328 284928
rect 236184 278044 236236 278050
rect 236184 277986 236236 277992
rect 236092 276684 236144 276690
rect 236092 276626 236144 276632
rect 235080 253224 235132 253230
rect 235080 253166 235132 253172
rect 236380 250510 236408 308230
rect 237116 307834 237144 308518
rect 236644 307828 236696 307834
rect 236644 307770 236696 307776
rect 237104 307828 237156 307834
rect 237104 307770 237156 307776
rect 236656 258738 236684 307770
rect 237392 300150 237420 310406
rect 237564 308440 237616 308446
rect 237564 308382 237616 308388
rect 237668 308394 237696 310420
rect 237472 308372 237524 308378
rect 237472 308314 237524 308320
rect 237380 300144 237432 300150
rect 237380 300086 237432 300092
rect 236644 258732 236696 258738
rect 236644 258674 236696 258680
rect 236368 250504 236420 250510
rect 236368 250446 236420 250452
rect 233516 244996 233568 245002
rect 233516 244938 233568 244944
rect 233332 244928 233384 244934
rect 233332 244870 233384 244876
rect 99286 168056 99342 168065
rect 99286 167991 99342 168000
rect 97908 159928 97960 159934
rect 97908 159870 97960 159876
rect 160926 159896 160982 159905
rect 160926 159831 160982 159840
rect 163502 159896 163558 159905
rect 163502 159831 163558 159840
rect 165986 159896 166042 159905
rect 165986 159831 166042 159840
rect 203430 159896 203486 159905
rect 203430 159831 203486 159840
rect 97816 159724 97868 159730
rect 97816 159666 97868 159672
rect 160940 158982 160968 159831
rect 163516 159186 163544 159831
rect 163504 159180 163556 159186
rect 163504 159122 163556 159128
rect 166000 159050 166028 159831
rect 200118 159352 200174 159361
rect 200118 159287 200174 159296
rect 165988 159044 166040 159050
rect 165988 158986 166040 158992
rect 160928 158976 160980 158982
rect 160928 158918 160980 158924
rect 158536 158908 158588 158914
rect 158536 158850 158588 158856
rect 119712 158704 119764 158710
rect 116858 158672 116914 158681
rect 116858 158607 116914 158616
rect 119710 158672 119712 158681
rect 158548 158681 158576 158850
rect 168288 158840 168340 158846
rect 168288 158782 168340 158788
rect 168300 158681 168328 158782
rect 119764 158672 119766 158681
rect 119710 158607 119766 158616
rect 121182 158672 121238 158681
rect 121182 158607 121238 158616
rect 122102 158672 122158 158681
rect 122102 158607 122158 158616
rect 123206 158672 123262 158681
rect 123206 158607 123262 158616
rect 125322 158672 125378 158681
rect 125322 158607 125378 158616
rect 126518 158672 126574 158681
rect 126518 158607 126574 158616
rect 127622 158672 127678 158681
rect 127622 158607 127678 158616
rect 128726 158672 128782 158681
rect 128726 158607 128782 158616
rect 130198 158672 130254 158681
rect 130198 158607 130254 158616
rect 131302 158672 131358 158681
rect 131302 158607 131304 158616
rect 97632 157684 97684 157690
rect 97632 157626 97684 157632
rect 116872 156330 116900 158607
rect 121196 158438 121224 158607
rect 121184 158432 121236 158438
rect 121184 158374 121236 158380
rect 122116 158302 122144 158607
rect 122104 158296 122156 158302
rect 117226 158264 117282 158273
rect 117282 158222 117360 158250
rect 122104 158238 122156 158244
rect 117226 158199 117282 158208
rect 117332 156398 117360 158222
rect 118238 157448 118294 157457
rect 118238 157383 118294 157392
rect 117320 156392 117372 156398
rect 117320 156334 117372 156340
rect 116860 156324 116912 156330
rect 116860 156266 116912 156272
rect 118252 153814 118280 157383
rect 123220 157214 123248 158607
rect 125336 157282 125364 158607
rect 125414 157992 125470 158001
rect 125414 157927 125470 157936
rect 125324 157276 125376 157282
rect 125324 157218 125376 157224
rect 123208 157208 123260 157214
rect 123208 157150 123260 157156
rect 125428 155922 125456 157927
rect 126532 157622 126560 158607
rect 127636 158098 127664 158607
rect 127624 158092 127676 158098
rect 127624 158034 127676 158040
rect 128740 157758 128768 158607
rect 130212 158574 130240 158607
rect 131356 158607 131358 158616
rect 132406 158672 132462 158681
rect 132406 158607 132462 158616
rect 133510 158672 133566 158681
rect 133510 158607 133566 158616
rect 134890 158672 134946 158681
rect 134890 158607 134946 158616
rect 158166 158672 158222 158681
rect 158166 158607 158222 158616
rect 158534 158672 158590 158681
rect 158534 158607 158590 158616
rect 159822 158672 159878 158681
rect 159822 158607 159878 158616
rect 168286 158672 168342 158681
rect 168286 158607 168342 158616
rect 191102 158672 191158 158681
rect 191102 158607 191158 158616
rect 131304 158578 131356 158584
rect 130200 158568 130252 158574
rect 130200 158510 130252 158516
rect 128728 157752 128780 157758
rect 128728 157694 128780 157700
rect 126520 157616 126572 157622
rect 126520 157558 126572 157564
rect 132420 157554 132448 158607
rect 133524 158166 133552 158607
rect 133512 158160 133564 158166
rect 133512 158102 133564 158108
rect 132408 157548 132460 157554
rect 132408 157490 132460 157496
rect 134904 157078 134932 158607
rect 135902 158536 135958 158545
rect 135902 158471 135958 158480
rect 137006 158536 137062 158545
rect 137006 158471 137062 158480
rect 139214 158536 139270 158545
rect 139214 158471 139270 158480
rect 140686 158536 140742 158545
rect 140686 158471 140742 158480
rect 134892 157072 134944 157078
rect 134892 157014 134944 157020
rect 135916 157010 135944 158471
rect 136086 157448 136142 157457
rect 136086 157383 136142 157392
rect 135904 157004 135956 157010
rect 135904 156946 135956 156952
rect 125598 156632 125654 156641
rect 125598 156567 125654 156576
rect 125416 155916 125468 155922
rect 125416 155858 125468 155864
rect 118240 153808 118292 153814
rect 118240 153750 118292 153756
rect 114560 138712 114612 138718
rect 114560 138654 114612 138660
rect 110420 137284 110472 137290
rect 110420 137226 110472 137232
rect 103520 135924 103572 135930
rect 103520 135866 103572 135872
rect 100760 127628 100812 127634
rect 100760 127570 100812 127576
rect 99380 91792 99432 91798
rect 99380 91734 99432 91740
rect 99392 16574 99420 91734
rect 99392 16546 99880 16574
rect 98644 3732 98696 3738
rect 98644 3674 98696 3680
rect 97448 3664 97500 3670
rect 97448 3606 97500 3612
rect 96252 3596 96304 3602
rect 96252 3538 96304 3544
rect 97264 3596 97316 3602
rect 97264 3538 97316 3544
rect 95148 3392 95200 3398
rect 95148 3334 95200 3340
rect 95160 480 95188 3334
rect 96264 480 96292 3538
rect 97460 480 97488 3606
rect 98656 480 98684 3674
rect 99852 480 99880 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100772 354 100800 127570
rect 103532 16574 103560 135866
rect 107660 129056 107712 129062
rect 107660 128998 107712 129004
rect 106280 104168 106332 104174
rect 106280 104110 106332 104116
rect 104900 64184 104952 64190
rect 104900 64126 104952 64132
rect 104912 16574 104940 64126
rect 106292 16574 106320 104110
rect 107672 16574 107700 128998
rect 109040 94512 109092 94518
rect 109040 94454 109092 94460
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102140 11756 102192 11762
rect 102140 11698 102192 11704
rect 102152 3602 102180 11698
rect 102232 3800 102284 3806
rect 102232 3742 102284 3748
rect 102140 3596 102192 3602
rect 102140 3538 102192 3544
rect 102244 480 102272 3742
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103428 3596 103480 3602
rect 103428 3538 103480 3544
rect 103348 480 103376 3538
rect 103440 3398 103468 3538
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 94454
rect 110432 3398 110460 137226
rect 111800 102808 111852 102814
rect 111800 102750 111852 102756
rect 111812 16574 111840 102750
rect 113824 90364 113876 90370
rect 113824 90306 113876 90312
rect 111812 16546 112392 16574
rect 110512 3936 110564 3942
rect 110512 3878 110564 3884
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 3878
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113836 3942 113864 90306
rect 114572 16574 114600 138654
rect 118700 130416 118752 130422
rect 118700 130358 118752 130364
rect 115940 93152 115992 93158
rect 115940 93094 115992 93100
rect 115952 16574 115980 93094
rect 117964 25560 118016 25566
rect 117964 25502 118016 25508
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 113824 3936 113876 3942
rect 113824 3878 113876 3884
rect 114008 3188 114060 3194
rect 114008 3130 114060 3136
rect 114020 480 114048 3130
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117596 3868 117648 3874
rect 117596 3810 117648 3816
rect 117608 480 117636 3810
rect 117976 3194 118004 25502
rect 118712 16574 118740 130358
rect 121460 97300 121512 97306
rect 121460 97242 121512 97248
rect 120080 86284 120132 86290
rect 120080 86226 120132 86232
rect 120092 16574 120120 86226
rect 121472 16574 121500 97242
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 117964 3188 118016 3194
rect 117964 3130 118016 3136
rect 118804 480 118832 16546
rect 119896 6180 119948 6186
rect 119896 6122 119948 6128
rect 119908 480 119936 6122
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 123484 8968 123536 8974
rect 123484 8910 123536 8916
rect 123496 480 123524 8910
rect 124680 3936 124732 3942
rect 124680 3878 124732 3884
rect 124692 480 124720 3878
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 156567
rect 133880 153876 133932 153882
rect 133880 153818 133932 153824
rect 132500 148368 132552 148374
rect 132500 148310 132552 148316
rect 128360 146940 128412 146946
rect 128360 146882 128412 146888
rect 126980 140072 127032 140078
rect 126980 140014 127032 140020
rect 126992 480 127020 140014
rect 127072 116612 127124 116618
rect 127072 116554 127124 116560
rect 127084 16574 127112 116554
rect 128372 16574 128400 146882
rect 129740 141432 129792 141438
rect 129740 141374 129792 141380
rect 129752 16574 129780 141374
rect 131120 106956 131172 106962
rect 131120 106898 131172 106904
rect 131132 16574 131160 106898
rect 132512 16574 132540 148310
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 153818
rect 136100 153202 136128 157383
rect 137020 156942 137048 158471
rect 138938 157448 138994 157457
rect 138938 157383 138994 157392
rect 137008 156936 137060 156942
rect 137008 156878 137060 156884
rect 136088 153196 136140 153202
rect 136088 153138 136140 153144
rect 138952 153134 138980 157383
rect 139228 156874 139256 158471
rect 140594 157992 140650 158001
rect 140594 157927 140650 157936
rect 139216 156868 139268 156874
rect 139216 156810 139268 156816
rect 140608 155718 140636 157927
rect 140700 156806 140728 158471
rect 150254 158400 150310 158409
rect 150254 158335 150310 158344
rect 141422 158264 141478 158273
rect 141422 158199 141478 158208
rect 141790 158264 141846 158273
rect 141790 158199 141846 158208
rect 146022 158264 146078 158273
rect 146022 158199 146078 158208
rect 146390 158264 146446 158273
rect 146390 158199 146446 158208
rect 140688 156800 140740 156806
rect 140688 156742 140740 156748
rect 140596 155712 140648 155718
rect 140596 155654 140648 155660
rect 138940 153128 138992 153134
rect 138940 153070 138992 153076
rect 141436 153066 141464 158199
rect 141804 155786 141832 158199
rect 144274 157856 144330 157865
rect 144274 157791 144330 157800
rect 145286 157856 145342 157865
rect 145286 157791 145342 157800
rect 143078 157584 143134 157593
rect 143078 157519 143134 157528
rect 141792 155780 141844 155786
rect 141792 155722 141844 155728
rect 143092 154902 143120 157519
rect 144288 155582 144316 157791
rect 144366 157448 144422 157457
rect 144366 157383 144422 157392
rect 144276 155576 144328 155582
rect 144276 155518 144328 155524
rect 143080 154896 143132 154902
rect 143080 154838 143132 154844
rect 141424 153060 141476 153066
rect 141424 153002 141476 153008
rect 144380 152998 144408 157383
rect 145300 155650 145328 157791
rect 145288 155644 145340 155650
rect 145288 155586 145340 155592
rect 144368 152992 144420 152998
rect 144368 152934 144420 152940
rect 146036 152930 146064 158199
rect 146404 155446 146432 158199
rect 148782 157856 148838 157865
rect 148782 157791 148838 157800
rect 147770 157584 147826 157593
rect 147770 157519 147826 157528
rect 146392 155440 146444 155446
rect 146392 155382 146444 155388
rect 147784 154970 147812 157519
rect 148414 157448 148470 157457
rect 148414 157383 148470 157392
rect 147772 154964 147824 154970
rect 147772 154906 147824 154912
rect 146024 152924 146076 152930
rect 146024 152866 146076 152872
rect 148428 152862 148456 157383
rect 148796 155378 148824 157791
rect 150268 156738 150296 158335
rect 150990 158264 151046 158273
rect 150990 158199 151046 158208
rect 150256 156732 150308 156738
rect 150256 156674 150308 156680
rect 148784 155372 148836 155378
rect 148784 155314 148836 155320
rect 148416 152856 148468 152862
rect 148416 152798 148468 152804
rect 151004 152794 151032 158199
rect 158180 157894 158208 158607
rect 159836 157962 159864 158607
rect 178958 158400 179014 158409
rect 178958 158335 179014 158344
rect 181718 158400 181774 158409
rect 181718 158335 181774 158344
rect 159824 157956 159876 157962
rect 159824 157898 159876 157904
rect 158168 157888 158220 157894
rect 158168 157830 158220 157836
rect 151358 157448 151414 157457
rect 151358 157383 151414 157392
rect 152646 157448 152702 157457
rect 152646 157383 152702 157392
rect 153934 157448 153990 157457
rect 153934 157383 153990 157392
rect 154486 157448 154542 157457
rect 154486 157383 154542 157392
rect 155774 157448 155830 157457
rect 155774 157383 155830 157392
rect 157062 157448 157118 157457
rect 157062 157383 157118 157392
rect 151372 154222 151400 157383
rect 152660 154494 152688 157383
rect 152648 154488 152700 154494
rect 152648 154430 152700 154436
rect 151360 154216 151412 154222
rect 151360 154158 151412 154164
rect 153948 153746 153976 157383
rect 154500 154358 154528 157383
rect 154488 154352 154540 154358
rect 154488 154294 154540 154300
rect 155788 154290 155816 157383
rect 155776 154284 155828 154290
rect 155776 154226 155828 154232
rect 157076 154154 157104 157383
rect 178038 156768 178094 156777
rect 178038 156703 178094 156712
rect 160098 155272 160154 155281
rect 160098 155207 160154 155216
rect 157064 154148 157116 154154
rect 157064 154090 157116 154096
rect 153936 153740 153988 153746
rect 153936 153682 153988 153688
rect 150992 152788 151044 152794
rect 150992 152730 151044 152736
rect 135260 152516 135312 152522
rect 135260 152458 135312 152464
rect 135272 4010 135300 152458
rect 146300 151088 146352 151094
rect 146300 151030 146352 151036
rect 139400 142860 139452 142866
rect 139400 142802 139452 142808
rect 138020 124908 138072 124914
rect 138020 124850 138072 124856
rect 136640 122120 136692 122126
rect 136640 122062 136692 122068
rect 135352 17332 135404 17338
rect 135352 17274 135404 17280
rect 135260 4004 135312 4010
rect 135260 3946 135312 3952
rect 135364 3482 135392 17274
rect 136652 16574 136680 122062
rect 138032 16574 138060 124850
rect 139412 16574 139440 142802
rect 143540 141500 143592 141506
rect 143540 141442 143592 141448
rect 140780 120760 140832 120766
rect 140780 120702 140832 120708
rect 140792 16574 140820 120702
rect 142160 101448 142212 101454
rect 142160 101390 142212 101396
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 4004 136508 4010
rect 136456 3946 136508 3952
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3946
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 101390
rect 143552 480 143580 141442
rect 143632 119400 143684 119406
rect 143632 119342 143684 119348
rect 143644 16574 143672 119342
rect 144920 22772 144972 22778
rect 144920 22714 144972 22720
rect 144932 16574 144960 22714
rect 146312 16574 146340 151030
rect 153200 149728 153252 149734
rect 153200 149670 153252 149676
rect 150440 144220 150492 144226
rect 150440 144162 150492 144168
rect 147680 134564 147732 134570
rect 147680 134506 147732 134512
rect 147692 16574 147720 134506
rect 149060 100020 149112 100026
rect 149060 99962 149112 99968
rect 149072 16574 149100 99962
rect 150452 16574 150480 144162
rect 151820 117972 151872 117978
rect 151820 117914 151872 117920
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 117914
rect 151912 24132 151964 24138
rect 151912 24074 151964 24080
rect 151924 16574 151952 24074
rect 153212 16574 153240 149670
rect 157340 145580 157392 145586
rect 157340 145522 157392 145528
rect 154580 144288 154632 144294
rect 154580 144230 154632 144236
rect 154592 16574 154620 144230
rect 155960 126268 156012 126274
rect 155960 126210 156012 126216
rect 155972 16574 156000 126210
rect 157352 16574 157380 145522
rect 158720 133204 158772 133210
rect 158720 133146 158772 133152
rect 158732 16574 158760 133146
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11830 160140 155207
rect 168380 153944 168432 153950
rect 168380 153886 168432 153892
rect 161480 138780 161532 138786
rect 161480 138722 161532 138728
rect 160192 98660 160244 98666
rect 160192 98602 160244 98608
rect 160100 11824 160152 11830
rect 160100 11766 160152 11772
rect 160204 6914 160232 98602
rect 161492 16574 161520 138722
rect 165620 137352 165672 137358
rect 165620 137294 165672 137300
rect 162860 115252 162912 115258
rect 162860 115194 162912 115200
rect 162872 16574 162900 115194
rect 165632 16574 165660 137294
rect 167000 112464 167052 112470
rect 167000 112406 167052 112412
rect 167012 16574 167040 112406
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11824 161348 11830
rect 161296 11766 161348 11772
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11766
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 164884 4004 164936 4010
rect 164884 3946 164936 3952
rect 164896 480 164924 3946
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 153886
rect 171140 152584 171192 152590
rect 171140 152526 171192 152532
rect 168472 135992 168524 135998
rect 168472 135934 168524 135940
rect 168484 16574 168512 135934
rect 169760 113824 169812 113830
rect 169760 113766 169812 113772
rect 169772 16574 169800 113766
rect 171152 16574 171180 152526
rect 175280 151156 175332 151162
rect 175280 151098 175332 151104
rect 172520 134632 172572 134638
rect 172520 134574 172572 134580
rect 172532 16574 172560 134574
rect 173900 123480 173952 123486
rect 173900 123422 173952 123428
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 169588 480 169616 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 123422
rect 175292 16574 175320 151098
rect 176660 147008 176712 147014
rect 176660 146950 176712 146956
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 480 176700 146950
rect 178052 16574 178080 156703
rect 178972 156670 179000 158335
rect 178960 156664 179012 156670
rect 178960 156606 179012 156612
rect 181732 156602 181760 158335
rect 185950 158128 186006 158137
rect 185950 158063 186006 158072
rect 181720 156596 181772 156602
rect 181720 156538 181772 156544
rect 185964 155961 185992 158063
rect 191116 157826 191144 158607
rect 195886 158400 195942 158409
rect 195886 158335 195942 158344
rect 198462 158400 198518 158409
rect 198462 158335 198518 158344
rect 193954 157856 194010 157865
rect 191104 157820 191156 157826
rect 193954 157791 194010 157800
rect 191104 157762 191156 157768
rect 185950 155952 186006 155961
rect 185950 155887 186006 155896
rect 182178 155408 182234 155417
rect 182178 155343 182234 155352
rect 179420 133272 179472 133278
rect 179420 133214 179472 133220
rect 179432 16574 179460 133214
rect 180800 111104 180852 111110
rect 180800 111046 180852 111052
rect 180812 16574 180840 111046
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 4820 177908 4826
rect 177856 4762 177908 4768
rect 177868 480 177896 4762
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 155343
rect 193968 155310 193996 157791
rect 193956 155304 194008 155310
rect 193956 155246 194008 155252
rect 195900 155242 195928 158335
rect 198476 156534 198504 158335
rect 198464 156528 198516 156534
rect 198464 156470 198516 156476
rect 195888 155236 195940 155242
rect 195888 155178 195940 155184
rect 193220 154012 193272 154018
rect 193220 153954 193272 153960
rect 184940 149796 184992 149802
rect 184940 149738 184992 149744
rect 183560 131776 183612 131782
rect 183560 131718 183612 131724
rect 183572 16574 183600 131718
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 149738
rect 189080 148436 189132 148442
rect 189080 148378 189132 148384
rect 186320 130484 186372 130490
rect 186320 130426 186372 130432
rect 185032 109744 185084 109750
rect 185032 109686 185084 109692
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 185044 6914 185072 109686
rect 186332 16574 186360 130426
rect 187700 108316 187752 108322
rect 187700 108258 187752 108264
rect 187712 16574 187740 108258
rect 189092 16574 189120 148378
rect 191840 131844 191892 131850
rect 191840 131786 191892 131792
rect 190460 129124 190512 129130
rect 190460 129066 190512 129072
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 129066
rect 191852 16574 191880 131786
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 153954
rect 195980 145648 196032 145654
rect 195980 145590 196032 145596
rect 193312 142928 193364 142934
rect 193312 142870 193364 142876
rect 193324 16574 193352 142870
rect 194600 18624 194652 18630
rect 194600 18566 194652 18572
rect 194612 16574 194640 18566
rect 195992 16574 196020 145590
rect 197360 140140 197412 140146
rect 197360 140082 197412 140088
rect 197372 16574 197400 140082
rect 198740 105596 198792 105602
rect 198740 105538 198792 105544
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 105538
rect 200132 16574 200160 159287
rect 203444 159118 203472 159831
rect 213918 159488 213974 159497
rect 213918 159423 213974 159432
rect 203432 159112 203484 159118
rect 203432 159054 203484 159060
rect 201038 157584 201094 157593
rect 201038 157519 201094 157528
rect 206282 157584 206338 157593
rect 206282 157519 206338 157528
rect 201052 155174 201080 157519
rect 202878 156904 202934 156913
rect 202878 156839 202934 156848
rect 201040 155168 201092 155174
rect 201040 155110 201092 155116
rect 201500 148504 201552 148510
rect 201500 148446 201552 148452
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 148446
rect 201592 19984 201644 19990
rect 201592 19926 201644 19932
rect 201604 16574 201632 19926
rect 202892 16574 202920 156839
rect 206296 155106 206324 157519
rect 206284 155100 206336 155106
rect 206284 155042 206336 155048
rect 207020 152652 207072 152658
rect 207020 152594 207072 152600
rect 205640 130552 205692 130558
rect 205640 130494 205692 130500
rect 204260 127696 204312 127702
rect 204260 127638 204312 127644
rect 204272 16574 204300 127638
rect 205652 16574 205680 130494
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 152594
rect 209780 151224 209832 151230
rect 209780 151166 209832 151172
rect 208400 138848 208452 138854
rect 208400 138790 208452 138796
rect 208412 16574 208440 138790
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 151166
rect 211160 126336 211212 126342
rect 211160 126278 211212 126284
rect 209872 104236 209924 104242
rect 209872 104178 209924 104184
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 104178
rect 211172 16574 211200 126278
rect 212540 21412 212592 21418
rect 212540 21354 212592 21360
rect 212552 16574 212580 21354
rect 213932 16574 213960 159423
rect 234620 159384 234672 159390
rect 234620 159326 234672 159332
rect 231860 156460 231912 156466
rect 231860 156402 231912 156408
rect 220818 155544 220874 155553
rect 220818 155479 220874 155488
rect 218060 149864 218112 149870
rect 218060 149806 218112 149812
rect 216680 147076 216732 147082
rect 216680 147018 216732 147024
rect 215300 137420 215352 137426
rect 215300 137362 215352 137368
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 137362
rect 216692 16574 216720 147018
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 149806
rect 218152 124976 218204 124982
rect 218152 124918 218204 124924
rect 218164 16574 218192 124918
rect 219440 102876 219492 102882
rect 219440 102818 219492 102824
rect 219452 16574 219480 102818
rect 220832 16574 220860 155479
rect 227720 154080 227772 154086
rect 227720 154022 227772 154028
rect 224960 144356 225012 144362
rect 224960 144298 225012 144304
rect 223580 141568 223632 141574
rect 223580 141510 223632 141516
rect 222200 136060 222252 136066
rect 222200 136002 222252 136008
rect 222212 16574 222240 136002
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 141510
rect 224972 16574 225000 144298
rect 226340 123548 226392 123554
rect 226340 123490 226392 123496
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 123490
rect 227732 16574 227760 154022
rect 229100 145716 229152 145722
rect 229100 145658 229152 145664
rect 229112 16574 229140 145658
rect 230480 129192 230532 129198
rect 230480 129134 230532 129140
rect 230492 16574 230520 129134
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227536 7608 227588 7614
rect 227536 7550 227588 7556
rect 227548 480 227576 7550
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 156402
rect 233240 155032 233292 155038
rect 233240 154974 233292 154980
rect 233252 16574 233280 154974
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11830 234660 159326
rect 236000 152720 236052 152726
rect 236000 152662 236052 152668
rect 234712 122188 234764 122194
rect 234712 122130 234764 122136
rect 234620 11824 234672 11830
rect 234620 11766 234672 11772
rect 234724 6914 234752 122130
rect 236012 16574 236040 152662
rect 237484 33794 237512 308314
rect 237576 275330 237604 308382
rect 237668 308366 237788 308394
rect 237656 308304 237708 308310
rect 237656 308246 237708 308252
rect 237668 286346 237696 308246
rect 237760 290494 237788 308366
rect 237748 290488 237800 290494
rect 237748 290430 237800 290436
rect 237656 286340 237708 286346
rect 237656 286282 237708 286288
rect 237564 275324 237616 275330
rect 237564 275266 237616 275272
rect 237472 33788 237524 33794
rect 237472 33730 237524 33736
rect 236012 16546 236592 16574
rect 235816 11824 235868 11830
rect 235816 11766 235868 11772
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11766
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237852 14482 237880 310420
rect 237944 310406 238142 310434
rect 237944 308446 237972 310406
rect 238116 308508 238168 308514
rect 238116 308450 238168 308456
rect 237932 308440 237984 308446
rect 237932 308382 237984 308388
rect 238022 308408 238078 308417
rect 238022 308343 238078 308352
rect 238036 159089 238064 308343
rect 238022 159080 238078 159089
rect 238128 159050 238156 308450
rect 238312 308310 238340 310420
rect 238404 310406 238602 310434
rect 238404 308378 238432 310406
rect 238772 308446 238800 310420
rect 238970 310406 239076 310434
rect 238944 308576 238996 308582
rect 238944 308518 238996 308524
rect 238760 308440 238812 308446
rect 238760 308382 238812 308388
rect 238392 308372 238444 308378
rect 238392 308314 238444 308320
rect 238852 308372 238904 308378
rect 238852 308314 238904 308320
rect 238300 308304 238352 308310
rect 238300 308246 238352 308252
rect 238760 308236 238812 308242
rect 238760 308178 238812 308184
rect 238772 298858 238800 308178
rect 238864 300218 238892 308314
rect 238852 300212 238904 300218
rect 238852 300154 238904 300160
rect 238760 298852 238812 298858
rect 238760 298794 238812 298800
rect 238956 271182 238984 308518
rect 239048 272542 239076 310406
rect 239128 308440 239180 308446
rect 239128 308382 239180 308388
rect 239232 308394 239260 310420
rect 239140 301510 239168 308382
rect 239232 308366 239352 308394
rect 239416 308378 239444 310420
rect 239600 308582 239628 310420
rect 239692 310406 239890 310434
rect 239588 308576 239640 308582
rect 239588 308518 239640 308524
rect 239220 308304 239272 308310
rect 239220 308246 239272 308252
rect 239128 301504 239180 301510
rect 239128 301446 239180 301452
rect 239036 272536 239088 272542
rect 239036 272478 239088 272484
rect 238944 271176 238996 271182
rect 238944 271118 238996 271124
rect 238208 265872 238260 265878
rect 238208 265814 238260 265820
rect 238022 159015 238078 159024
rect 238116 159044 238168 159050
rect 238116 158986 238168 158992
rect 238220 158273 238248 265814
rect 238392 250640 238444 250646
rect 238392 250582 238444 250588
rect 238300 170400 238352 170406
rect 238300 170342 238352 170348
rect 238312 159594 238340 170342
rect 238300 159588 238352 159594
rect 238300 159530 238352 159536
rect 238206 158264 238262 158273
rect 238206 158199 238262 158208
rect 238404 158137 238432 250582
rect 238484 167680 238536 167686
rect 238484 167622 238536 167628
rect 238496 159662 238524 167622
rect 238484 159656 238536 159662
rect 238484 159598 238536 159604
rect 238390 158128 238446 158137
rect 238390 158063 238446 158072
rect 237840 14476 237892 14482
rect 237840 14418 237892 14424
rect 237656 10396 237708 10402
rect 237656 10338 237708 10344
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 10338
rect 239232 10334 239260 308246
rect 239324 89010 239352 308366
rect 239404 308372 239456 308378
rect 239404 308314 239456 308320
rect 239692 308310 239720 310406
rect 239680 308304 239732 308310
rect 239680 308246 239732 308252
rect 240060 308242 240088 310420
rect 240048 308236 240100 308242
rect 240048 308178 240100 308184
rect 239404 298784 239456 298790
rect 239404 298726 239456 298732
rect 239312 89004 239364 89010
rect 239312 88946 239364 88952
rect 239220 10328 239272 10334
rect 239220 10270 239272 10276
rect 239312 4072 239364 4078
rect 239312 4014 239364 4020
rect 239324 480 239352 4014
rect 239416 3874 239444 298726
rect 240244 269822 240272 310420
rect 240428 310406 240534 310434
rect 240324 308440 240376 308446
rect 240324 308382 240376 308388
rect 240336 283694 240364 308382
rect 240428 289202 240456 310406
rect 240704 307154 240732 310420
rect 240692 307148 240744 307154
rect 240692 307090 240744 307096
rect 240888 307034 240916 310420
rect 240980 310406 241178 310434
rect 240980 308446 241008 310406
rect 240968 308440 241020 308446
rect 240968 308382 241020 308388
rect 240520 307006 240916 307034
rect 240416 289196 240468 289202
rect 240416 289138 240468 289144
rect 240324 283688 240376 283694
rect 240324 283630 240376 283636
rect 240232 269816 240284 269822
rect 240232 269758 240284 269764
rect 240520 268394 240548 307006
rect 241348 297498 241376 310420
rect 241532 310406 241638 310434
rect 241532 306474 241560 310406
rect 241808 308650 241836 310420
rect 241796 308644 241848 308650
rect 241796 308586 241848 308592
rect 241992 308394 242020 310420
rect 241716 308366 242020 308394
rect 242084 310406 242282 310434
rect 241612 308304 241664 308310
rect 241612 308246 241664 308252
rect 241520 306468 241572 306474
rect 241520 306410 241572 306416
rect 241336 297492 241388 297498
rect 241336 297434 241388 297440
rect 241624 294642 241652 308246
rect 241716 296002 241744 308366
rect 242084 307816 242112 310406
rect 242452 309074 242480 310420
rect 241900 307788 242112 307816
rect 242176 309046 242480 309074
rect 241796 306468 241848 306474
rect 241796 306410 241848 306416
rect 241808 297430 241836 306410
rect 241796 297424 241848 297430
rect 241796 297366 241848 297372
rect 241704 295996 241756 296002
rect 241704 295938 241756 295944
rect 241612 294636 241664 294642
rect 241612 294578 241664 294584
rect 240508 268388 240560 268394
rect 240508 268330 240560 268336
rect 241900 265674 241928 307788
rect 242176 307714 242204 309046
rect 242256 308984 242308 308990
rect 242256 308926 242308 308932
rect 241992 307686 242204 307714
rect 241992 305658 242020 307686
rect 242164 307624 242216 307630
rect 242164 307566 242216 307572
rect 241980 305652 242032 305658
rect 241980 305594 242032 305600
rect 241888 265668 241940 265674
rect 241888 265610 241940 265616
rect 242176 13122 242204 307566
rect 242268 86290 242296 308926
rect 242636 308310 242664 310420
rect 242912 308446 242940 310420
rect 242900 308440 242952 308446
rect 242900 308382 242952 308388
rect 243096 308394 243124 310420
rect 242992 308372 243044 308378
rect 243096 308366 243216 308394
rect 242992 308314 243044 308320
rect 242624 308304 242676 308310
rect 242624 308246 242676 308252
rect 242532 308100 242584 308106
rect 242532 308042 242584 308048
rect 242544 296714 242572 308042
rect 243004 304366 243032 308314
rect 243084 308304 243136 308310
rect 243084 308246 243136 308252
rect 242992 304360 243044 304366
rect 242992 304302 243044 304308
rect 242360 296686 242572 296714
rect 242360 129062 242388 296686
rect 243096 290562 243124 308246
rect 243188 308174 243216 308366
rect 243176 308168 243228 308174
rect 243176 308110 243228 308116
rect 243280 307816 243308 310420
rect 243188 307788 243308 307816
rect 243372 310406 243570 310434
rect 243188 291922 243216 307788
rect 243268 307692 243320 307698
rect 243268 307634 243320 307640
rect 243176 291916 243228 291922
rect 243176 291858 243228 291864
rect 243084 290556 243136 290562
rect 243084 290498 243136 290504
rect 243280 262954 243308 307634
rect 243372 264246 243400 310406
rect 243544 308644 243596 308650
rect 243544 308586 243596 308592
rect 243452 308440 243504 308446
rect 243452 308382 243504 308388
rect 243464 296070 243492 308382
rect 243452 296064 243504 296070
rect 243452 296006 243504 296012
rect 243360 264240 243412 264246
rect 243360 264182 243412 264188
rect 243268 262948 243320 262954
rect 243268 262890 243320 262896
rect 242348 129056 242400 129062
rect 242348 128998 242400 129004
rect 242256 86284 242308 86290
rect 242256 86226 242308 86232
rect 242900 15904 242952 15910
rect 242900 15846 242952 15852
rect 242164 13116 242216 13122
rect 242164 13058 242216 13064
rect 241704 9036 241756 9042
rect 241704 8978 241756 8984
rect 240508 7676 240560 7682
rect 240508 7618 240560 7624
rect 239404 3868 239456 3874
rect 239404 3810 239456 3816
rect 240520 480 240548 7618
rect 241716 480 241744 8978
rect 242912 480 242940 15846
rect 243556 8974 243584 308586
rect 243740 308378 243768 310420
rect 243832 310406 244030 310434
rect 243728 308372 243780 308378
rect 243728 308314 243780 308320
rect 243832 308310 243860 310406
rect 243820 308304 243872 308310
rect 243820 308246 243872 308252
rect 243728 308032 243780 308038
rect 243728 307974 243780 307980
rect 243636 290488 243688 290494
rect 243636 290430 243688 290436
rect 243544 8968 243596 8974
rect 243544 8910 243596 8916
rect 243648 3942 243676 290430
rect 243740 135930 243768 307974
rect 244200 307698 244228 310420
rect 244188 307692 244240 307698
rect 244188 307634 244240 307640
rect 244384 303074 244412 310420
rect 244568 310406 244674 310434
rect 244464 306332 244516 306338
rect 244464 306274 244516 306280
rect 244372 303068 244424 303074
rect 244372 303010 244424 303016
rect 244372 302932 244424 302938
rect 244372 302874 244424 302880
rect 243728 135924 243780 135930
rect 243728 135866 243780 135872
rect 244096 4888 244148 4894
rect 244096 4830 244148 4836
rect 243636 3936 243688 3942
rect 243636 3878 243688 3884
rect 244108 480 244136 4830
rect 244384 3534 244412 302874
rect 244476 261594 244504 306274
rect 244464 261588 244516 261594
rect 244464 261530 244516 261536
rect 244372 3528 244424 3534
rect 244372 3470 244424 3476
rect 244568 3466 244596 310406
rect 244844 307222 244872 310420
rect 244924 307964 244976 307970
rect 244924 307906 244976 307912
rect 244832 307216 244884 307222
rect 244832 307158 244884 307164
rect 244936 137290 244964 307906
rect 245028 307834 245056 310420
rect 245120 310406 245318 310434
rect 245016 307828 245068 307834
rect 245016 307770 245068 307776
rect 245120 302938 245148 310406
rect 245488 306338 245516 310420
rect 245686 310406 245884 310434
rect 245856 306882 245884 310406
rect 245844 306876 245896 306882
rect 245844 306818 245896 306824
rect 245948 306762 245976 310420
rect 245672 306734 245976 306762
rect 245476 306332 245528 306338
rect 245476 306274 245528 306280
rect 245672 303142 245700 306734
rect 245844 306604 245896 306610
rect 245844 306546 245896 306552
rect 245752 306468 245804 306474
rect 245752 306410 245804 306416
rect 245660 303136 245712 303142
rect 245660 303078 245712 303084
rect 245108 302932 245160 302938
rect 245108 302874 245160 302880
rect 245764 279546 245792 306410
rect 245856 280906 245884 306546
rect 245936 306536 245988 306542
rect 245936 306478 245988 306484
rect 245948 286414 245976 306478
rect 246132 306354 246160 310420
rect 246316 306474 246344 310420
rect 246408 310406 246606 310434
rect 246408 306542 246436 310406
rect 246488 307896 246540 307902
rect 246488 307838 246540 307844
rect 246396 306536 246448 306542
rect 246396 306478 246448 306484
rect 246304 306468 246356 306474
rect 246304 306410 246356 306416
rect 246040 306326 246160 306354
rect 246040 293282 246068 306326
rect 246120 306264 246172 306270
rect 246500 306218 246528 307838
rect 246776 306270 246804 310420
rect 246856 307828 246908 307834
rect 246856 307770 246908 307776
rect 246120 306206 246172 306212
rect 246028 293276 246080 293282
rect 246028 293218 246080 293224
rect 245936 286408 245988 286414
rect 245936 286350 245988 286356
rect 245844 280900 245896 280906
rect 245844 280842 245896 280848
rect 245752 279540 245804 279546
rect 245752 279482 245804 279488
rect 246132 260234 246160 306206
rect 246316 306190 246528 306218
rect 246764 306264 246816 306270
rect 246764 306206 246816 306212
rect 246120 260228 246172 260234
rect 246120 260170 246172 260176
rect 244924 137284 244976 137290
rect 244924 137226 244976 137232
rect 246316 11762 246344 306190
rect 246868 302234 246896 307770
rect 247052 306338 247080 310420
rect 247236 306354 247264 310420
rect 247434 310406 247540 310434
rect 247316 306468 247368 306474
rect 247316 306410 247368 306416
rect 247040 306332 247092 306338
rect 247040 306274 247092 306280
rect 247144 306326 247264 306354
rect 246408 302206 246896 302234
rect 246408 127634 246436 302206
rect 247144 301578 247172 306326
rect 247224 306264 247276 306270
rect 247224 306206 247276 306212
rect 247132 301572 247184 301578
rect 247132 301514 247184 301520
rect 246396 127628 246448 127634
rect 246396 127570 246448 127576
rect 246304 11756 246356 11762
rect 246304 11698 246356 11704
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 244556 3460 244608 3466
rect 244556 3402 244608 3408
rect 245212 480 245240 3810
rect 247236 3670 247264 306206
rect 247328 91798 247356 306410
rect 247408 306400 247460 306406
rect 247408 306342 247460 306348
rect 247316 91792 247368 91798
rect 247316 91734 247368 91740
rect 247420 3738 247448 306342
rect 247408 3732 247460 3738
rect 247408 3674 247460 3680
rect 247224 3664 247276 3670
rect 247224 3606 247276 3612
rect 247512 3602 247540 310406
rect 247696 309058 247724 310420
rect 247684 309052 247736 309058
rect 247684 308994 247736 309000
rect 247774 308544 247830 308553
rect 247774 308479 247830 308488
rect 247684 308440 247736 308446
rect 247684 308382 247736 308388
rect 247592 306332 247644 306338
rect 247592 306274 247644 306280
rect 247604 301646 247632 306274
rect 247592 301640 247644 301646
rect 247592 301582 247644 301588
rect 247696 145586 247724 308382
rect 247788 159225 247816 308479
rect 247880 306270 247908 310420
rect 248064 306406 248092 310420
rect 248156 310406 248354 310434
rect 248156 306474 248184 310406
rect 248524 307834 248552 310420
rect 248512 307828 248564 307834
rect 248512 307770 248564 307776
rect 248144 306468 248196 306474
rect 248144 306410 248196 306416
rect 248052 306400 248104 306406
rect 248052 306342 248104 306348
rect 248512 306400 248564 306406
rect 248512 306342 248564 306348
rect 247868 306264 247920 306270
rect 247868 306206 247920 306212
rect 247774 159216 247830 159225
rect 247774 159151 247830 159160
rect 247684 145580 247736 145586
rect 247684 145522 247736 145528
rect 248524 64190 248552 306342
rect 248604 306332 248656 306338
rect 248604 306274 248656 306280
rect 248616 104174 248644 306274
rect 248604 104168 248656 104174
rect 248604 104110 248656 104116
rect 248512 64184 248564 64190
rect 248512 64126 248564 64132
rect 247592 6248 247644 6254
rect 247592 6190 247644 6196
rect 247500 3596 247552 3602
rect 247500 3538 247552 3544
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246408 480 246436 3402
rect 247604 480 247632 6190
rect 248708 3806 248736 310420
rect 248984 307902 249012 310420
rect 249168 308038 249196 310420
rect 249260 310406 249458 310434
rect 249156 308032 249208 308038
rect 249156 307974 249208 307980
rect 248972 307896 249024 307902
rect 248972 307838 249024 307844
rect 249064 307828 249116 307834
rect 249064 307770 249116 307776
rect 249076 93158 249104 307770
rect 249260 306406 249288 310406
rect 249340 308848 249392 308854
rect 249340 308790 249392 308796
rect 249248 306400 249300 306406
rect 249248 306342 249300 306348
rect 249352 296714 249380 308790
rect 249628 306338 249656 310420
rect 249812 308106 249840 310420
rect 249996 310406 250102 310434
rect 249800 308100 249852 308106
rect 249800 308042 249852 308048
rect 249892 306468 249944 306474
rect 249892 306410 249944 306416
rect 249616 306332 249668 306338
rect 249616 306274 249668 306280
rect 249168 296686 249380 296714
rect 249168 149734 249196 296686
rect 249156 149728 249208 149734
rect 249156 149670 249208 149676
rect 249064 93152 249116 93158
rect 249064 93094 249116 93100
rect 249904 90370 249932 306410
rect 249996 94518 250024 310406
rect 250076 306536 250128 306542
rect 250076 306478 250128 306484
rect 250088 102814 250116 306478
rect 250272 306474 250300 310420
rect 250456 307970 250484 310420
rect 250548 310406 250746 310434
rect 250444 307964 250496 307970
rect 250444 307906 250496 307912
rect 250548 306542 250576 310406
rect 250536 306536 250588 306542
rect 250536 306478 250588 306484
rect 250260 306468 250312 306474
rect 250260 306410 250312 306416
rect 250916 306354 250944 310420
rect 250996 308236 251048 308242
rect 250996 308178 251048 308184
rect 250272 306326 250944 306354
rect 250168 303748 250220 303754
rect 250168 303690 250220 303696
rect 250180 138718 250208 303690
rect 250168 138712 250220 138718
rect 250168 138654 250220 138660
rect 250076 102808 250128 102814
rect 250076 102750 250128 102756
rect 249984 94512 250036 94518
rect 249984 94454 250036 94460
rect 249892 90364 249944 90370
rect 249892 90306 249944 90312
rect 250272 25566 250300 306326
rect 251008 302234 251036 308178
rect 251100 303754 251128 310420
rect 251376 307834 251404 310420
rect 251560 309134 251588 310420
rect 251560 309106 251680 309134
rect 251364 307828 251416 307834
rect 251364 307770 251416 307776
rect 251180 307080 251232 307086
rect 251180 307022 251232 307028
rect 251088 303748 251140 303754
rect 251088 303690 251140 303696
rect 250548 302206 251036 302234
rect 250548 296714 250576 302206
rect 250456 296686 250576 296714
rect 250456 158914 250484 296686
rect 250444 158908 250496 158914
rect 250444 158850 250496 158856
rect 250260 25560 250312 25566
rect 250260 25502 250312 25508
rect 248788 8968 248840 8974
rect 248788 8910 248840 8916
rect 248696 3800 248748 3806
rect 248696 3742 248748 3748
rect 248800 480 248828 8910
rect 249984 3596 250036 3602
rect 249984 3538 250036 3544
rect 249996 480 250024 3538
rect 251192 3534 251220 307022
rect 251456 304292 251508 304298
rect 251456 304234 251508 304240
rect 251364 303136 251416 303142
rect 251364 303078 251416 303084
rect 251272 302728 251324 302734
rect 251272 302670 251324 302676
rect 251284 6186 251312 302670
rect 251376 97306 251404 303078
rect 251468 130422 251496 304234
rect 251652 299474 251680 309106
rect 251744 304298 251772 310420
rect 251836 310406 252034 310434
rect 251732 304292 251784 304298
rect 251732 304234 251784 304240
rect 251836 302734 251864 310406
rect 252204 308990 252232 310420
rect 252296 310406 252494 310434
rect 252192 308984 252244 308990
rect 252192 308926 252244 308932
rect 252008 308780 252060 308786
rect 252008 308722 252060 308728
rect 251916 308372 251968 308378
rect 251916 308314 251968 308320
rect 251824 302728 251876 302734
rect 251824 302670 251876 302676
rect 251928 302234 251956 308314
rect 251560 299446 251680 299474
rect 251836 302206 251956 302234
rect 251560 298790 251588 299446
rect 251548 298784 251600 298790
rect 251548 298726 251600 298732
rect 251836 148374 251864 302206
rect 252020 296714 252048 308722
rect 252296 303142 252324 310406
rect 252664 308718 252692 310420
rect 252862 310406 252968 310434
rect 252652 308712 252704 308718
rect 252652 308654 252704 308660
rect 252744 308712 252796 308718
rect 252744 308654 252796 308660
rect 252652 306400 252704 306406
rect 252652 306342 252704 306348
rect 252284 303136 252336 303142
rect 252284 303078 252336 303084
rect 251928 296686 252048 296714
rect 251928 158982 251956 296686
rect 251916 158976 251968 158982
rect 251916 158918 251968 158924
rect 251824 148368 251876 148374
rect 251824 148310 251876 148316
rect 252664 140078 252692 306342
rect 252756 146946 252784 308654
rect 252836 306332 252888 306338
rect 252836 306274 252888 306280
rect 252848 156641 252876 306274
rect 252940 290494 252968 310406
rect 253032 310406 253138 310434
rect 253032 306338 253060 310406
rect 253308 306406 253336 310420
rect 253296 306400 253348 306406
rect 253296 306342 253348 306348
rect 253020 306332 253072 306338
rect 253020 306274 253072 306280
rect 253492 305266 253520 310420
rect 253584 310406 253782 310434
rect 253584 308718 253612 310406
rect 253572 308712 253624 308718
rect 253572 308654 253624 308660
rect 253756 308644 253808 308650
rect 253756 308586 253808 308592
rect 253572 308576 253624 308582
rect 253572 308518 253624 308524
rect 253032 305238 253520 305266
rect 252928 290488 252980 290494
rect 252928 290430 252980 290436
rect 252834 156632 252890 156641
rect 252834 156567 252890 156576
rect 252744 146940 252796 146946
rect 252744 146882 252796 146888
rect 252652 140072 252704 140078
rect 252652 140014 252704 140020
rect 251456 130416 251508 130422
rect 251456 130358 251508 130364
rect 253032 116618 253060 305238
rect 253584 302234 253612 308518
rect 253768 308378 253796 308586
rect 253756 308372 253808 308378
rect 253756 308314 253808 308320
rect 253952 306338 253980 310420
rect 253940 306332 253992 306338
rect 253940 306274 253992 306280
rect 254136 306184 254164 310420
rect 254412 308650 254440 310420
rect 254400 308644 254452 308650
rect 254400 308586 254452 308592
rect 254216 306332 254268 306338
rect 254216 306274 254268 306280
rect 254308 306332 254360 306338
rect 254308 306274 254360 306280
rect 253216 302206 253612 302234
rect 254044 306156 254164 306184
rect 253216 151162 253244 302206
rect 253204 151156 253256 151162
rect 253204 151098 253256 151104
rect 253204 146940 253256 146946
rect 253204 146882 253256 146888
rect 253020 116612 253072 116618
rect 253020 116554 253072 116560
rect 251364 97300 251416 97306
rect 251364 97242 251416 97248
rect 251272 6180 251324 6186
rect 251272 6122 251324 6128
rect 253216 4078 253244 146882
rect 254044 106962 254072 306156
rect 254124 306060 254176 306066
rect 254124 306002 254176 306008
rect 254136 122126 254164 306002
rect 254228 141438 254256 306274
rect 254320 152522 254348 306274
rect 254596 302234 254624 310420
rect 254412 302206 254624 302234
rect 254688 310406 254886 310434
rect 254412 153882 254440 302206
rect 254688 296714 254716 310406
rect 255056 306338 255084 310420
rect 255044 306332 255096 306338
rect 255044 306274 255096 306280
rect 255240 306066 255268 310420
rect 255412 306400 255464 306406
rect 255412 306342 255464 306348
rect 255320 306332 255372 306338
rect 255320 306274 255372 306280
rect 255228 306060 255280 306066
rect 255228 306002 255280 306008
rect 254504 296686 254716 296714
rect 254400 153876 254452 153882
rect 254400 153818 254452 153824
rect 254308 152516 254360 152522
rect 254308 152458 254360 152464
rect 254216 141432 254268 141438
rect 254216 141374 254268 141380
rect 254124 122120 254176 122126
rect 254124 122062 254176 122068
rect 254032 106956 254084 106962
rect 254032 106898 254084 106904
rect 254504 17338 254532 296686
rect 255332 101454 255360 306274
rect 255424 119406 255452 306342
rect 255516 306320 255544 310420
rect 255700 306320 255728 310420
rect 255516 306292 255636 306320
rect 255700 306292 255820 306320
rect 255504 306196 255556 306202
rect 255504 306138 255556 306144
rect 255516 120766 255544 306138
rect 255608 124914 255636 306292
rect 255688 306128 255740 306134
rect 255688 306070 255740 306076
rect 255700 141506 255728 306070
rect 255792 142866 255820 306292
rect 255884 306202 255912 310420
rect 255976 310406 256174 310434
rect 255976 306338 256004 310406
rect 256056 308644 256108 308650
rect 256056 308586 256108 308592
rect 255964 306332 256016 306338
rect 255964 306274 256016 306280
rect 255872 306196 255924 306202
rect 255872 306138 255924 306144
rect 256068 296714 256096 308586
rect 256344 306134 256372 310420
rect 256528 306406 256556 310420
rect 256712 310406 256818 310434
rect 256516 306400 256568 306406
rect 256516 306342 256568 306348
rect 256332 306128 256384 306134
rect 256332 306070 256384 306076
rect 255976 296686 256096 296714
rect 255976 156777 256004 296686
rect 255962 156768 256018 156777
rect 255962 156703 256018 156712
rect 255780 142860 255832 142866
rect 255780 142802 255832 142808
rect 255688 141500 255740 141506
rect 255688 141442 255740 141448
rect 255596 124908 255648 124914
rect 255596 124850 255648 124856
rect 255504 120760 255556 120766
rect 255504 120702 255556 120708
rect 255964 120760 256016 120766
rect 255964 120702 256016 120708
rect 255412 119400 255464 119406
rect 255412 119342 255464 119348
rect 255320 101448 255372 101454
rect 255320 101390 255372 101396
rect 254492 17332 254544 17338
rect 254492 17274 254544 17280
rect 254032 17264 254084 17270
rect 254032 17206 254084 17212
rect 254044 16574 254072 17206
rect 254044 16546 254256 16574
rect 253204 4072 253256 4078
rect 253204 4014 253256 4020
rect 251272 3664 251324 3670
rect 251272 3606 251324 3612
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 251284 1850 251312 3606
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 253480 3528 253532 3534
rect 253480 3470 253532 3476
rect 251192 1822 251312 1850
rect 251192 480 251220 1822
rect 252388 480 252416 3470
rect 253492 480 253520 3470
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255872 13184 255924 13190
rect 255872 13126 255924 13132
rect 255884 480 255912 13126
rect 255976 3874 256004 120702
rect 256712 22778 256740 310406
rect 256988 306649 257016 310420
rect 256974 306640 257030 306649
rect 256974 306575 257030 306584
rect 257172 306474 257200 310420
rect 257264 310406 257462 310434
rect 256976 306468 257028 306474
rect 256976 306410 257028 306416
rect 257160 306468 257212 306474
rect 257160 306410 257212 306416
rect 256884 306400 256936 306406
rect 256884 306342 256936 306348
rect 256792 306332 256844 306338
rect 256792 306274 256844 306280
rect 256804 100026 256832 306274
rect 256896 117978 256924 306342
rect 256988 134570 257016 306410
rect 257158 306368 257214 306377
rect 257264 306338 257292 310406
rect 257344 307828 257396 307834
rect 257344 307770 257396 307776
rect 257158 306303 257214 306312
rect 257252 306332 257304 306338
rect 257068 306128 257120 306134
rect 257068 306070 257120 306076
rect 257080 144226 257108 306070
rect 257172 151094 257200 306303
rect 257252 306274 257304 306280
rect 257160 151088 257212 151094
rect 257160 151030 257212 151036
rect 257068 144220 257120 144226
rect 257068 144162 257120 144168
rect 256976 134564 257028 134570
rect 256976 134506 257028 134512
rect 256884 117972 256936 117978
rect 256884 117914 256936 117920
rect 256792 100020 256844 100026
rect 256792 99962 256844 99968
rect 257356 24138 257384 307770
rect 257632 306134 257660 310420
rect 257724 310406 257922 310434
rect 257724 306406 257752 310406
rect 258092 307834 258120 310420
rect 258276 308854 258304 310420
rect 258368 310406 258566 310434
rect 258264 308848 258316 308854
rect 258264 308790 258316 308796
rect 258080 307828 258132 307834
rect 258080 307770 258132 307776
rect 257712 306400 257764 306406
rect 257712 306342 257764 306348
rect 258264 306400 258316 306406
rect 258264 306342 258316 306348
rect 258172 306332 258224 306338
rect 258172 306274 258224 306280
rect 257620 306128 257672 306134
rect 257620 306070 257672 306076
rect 258184 126274 258212 306274
rect 258276 133210 258304 306342
rect 258368 144294 258396 310406
rect 258736 306338 258764 310420
rect 258920 308446 258948 310420
rect 259012 310406 259210 310434
rect 258908 308440 258960 308446
rect 258908 308382 258960 308388
rect 259012 306406 259040 310406
rect 259000 306400 259052 306406
rect 259000 306342 259052 306348
rect 258724 306332 258776 306338
rect 258724 306274 258776 306280
rect 259380 296714 259408 310420
rect 259460 306332 259512 306338
rect 259460 306274 259512 306280
rect 258460 296686 259408 296714
rect 258356 144288 258408 144294
rect 258356 144230 258408 144236
rect 258264 133204 258316 133210
rect 258264 133146 258316 133152
rect 258172 126268 258224 126274
rect 258172 126210 258224 126216
rect 258460 98666 258488 296686
rect 258448 98660 258500 98666
rect 258448 98602 258500 98608
rect 257344 24132 257396 24138
rect 257344 24074 257396 24080
rect 256700 22772 256752 22778
rect 256700 22714 256752 22720
rect 257068 6180 257120 6186
rect 257068 6122 257120 6128
rect 255964 3868 256016 3874
rect 255964 3810 256016 3816
rect 257080 480 257108 6122
rect 259472 4010 259500 306274
rect 259564 306270 259592 310420
rect 259748 310406 259854 310434
rect 259644 306400 259696 306406
rect 259644 306342 259696 306348
rect 259552 306264 259604 306270
rect 259552 306206 259604 306212
rect 259552 306128 259604 306134
rect 259552 306070 259604 306076
rect 259564 112470 259592 306070
rect 259656 115258 259684 306342
rect 259748 306252 259776 310406
rect 260024 306406 260052 310420
rect 260116 310406 260314 310434
rect 260012 306400 260064 306406
rect 260012 306342 260064 306348
rect 260116 306338 260144 310406
rect 260196 308440 260248 308446
rect 260196 308382 260248 308388
rect 260104 306332 260156 306338
rect 260104 306274 260156 306280
rect 259920 306264 259972 306270
rect 259748 306224 259868 306252
rect 259736 306060 259788 306066
rect 259736 306002 259788 306008
rect 259748 137358 259776 306002
rect 259840 138786 259868 306224
rect 259920 306206 259972 306212
rect 259932 155281 259960 306206
rect 260208 296714 260236 308382
rect 260484 306066 260512 310420
rect 260668 306134 260696 310420
rect 260840 306468 260892 306474
rect 260840 306410 260892 306416
rect 260656 306128 260708 306134
rect 260656 306070 260708 306076
rect 260472 306060 260524 306066
rect 260472 306002 260524 306008
rect 260116 296686 260236 296714
rect 259918 155272 259974 155281
rect 259918 155207 259974 155216
rect 259828 138780 259880 138786
rect 259828 138722 259880 138728
rect 259736 137352 259788 137358
rect 259736 137294 259788 137300
rect 259644 115252 259696 115258
rect 259644 115194 259696 115200
rect 259552 112464 259604 112470
rect 259552 112406 259604 112412
rect 260012 13116 260064 13122
rect 260012 13058 260064 13064
rect 259460 4004 259512 4010
rect 259460 3946 259512 3952
rect 259460 3732 259512 3738
rect 259460 3674 259512 3680
rect 258264 3596 258316 3602
rect 258264 3538 258316 3544
rect 258276 480 258304 3538
rect 259472 480 259500 3674
rect 260024 3482 260052 13058
rect 260116 4826 260144 296686
rect 260194 160712 260250 160721
rect 260194 160647 260250 160656
rect 260104 4820 260156 4826
rect 260104 4762 260156 4768
rect 260208 3602 260236 160647
rect 260852 113830 260880 306410
rect 260944 306202 260972 310420
rect 261024 306332 261076 306338
rect 261024 306274 261076 306280
rect 260932 306196 260984 306202
rect 260932 306138 260984 306144
rect 260932 306060 260984 306066
rect 260932 306002 260984 306008
rect 260944 123486 260972 306002
rect 261036 134638 261064 306274
rect 261128 135998 261156 310420
rect 261312 306474 261340 310420
rect 261404 310406 261602 310434
rect 261300 306468 261352 306474
rect 261300 306410 261352 306416
rect 261404 306320 261432 310406
rect 261772 306338 261800 310420
rect 261312 306292 261432 306320
rect 261760 306332 261812 306338
rect 261208 162172 261260 162178
rect 261208 162114 261260 162120
rect 261116 135992 261168 135998
rect 261116 135934 261168 135940
rect 261024 134632 261076 134638
rect 261024 134574 261076 134580
rect 260932 123480 260984 123486
rect 260932 123422 260984 123428
rect 260840 113824 260892 113830
rect 260840 113766 260892 113772
rect 261220 16574 261248 162114
rect 261312 152590 261340 306292
rect 261760 306274 261812 306280
rect 261392 306196 261444 306202
rect 261392 306138 261444 306144
rect 261404 153950 261432 306138
rect 261956 306066 261984 310420
rect 262232 308582 262260 310420
rect 262220 308576 262272 308582
rect 262220 308518 262272 308524
rect 262312 308372 262364 308378
rect 262312 308314 262364 308320
rect 261944 306060 261996 306066
rect 261944 306002 261996 306008
rect 261392 153944 261444 153950
rect 261392 153886 261444 153892
rect 261300 152584 261352 152590
rect 261300 152526 261352 152532
rect 261484 134564 261536 134570
rect 261484 134506 261536 134512
rect 261220 16546 261432 16574
rect 260196 3596 260248 3602
rect 260196 3538 260248 3544
rect 261404 3482 261432 16546
rect 261496 3874 261524 134506
rect 262324 133278 262352 308314
rect 262416 147014 262444 310420
rect 262496 308576 262548 308582
rect 262496 308518 262548 308524
rect 262508 308242 262536 308518
rect 262600 308446 262628 310420
rect 262876 308650 262904 310420
rect 262864 308644 262916 308650
rect 262864 308586 262916 308592
rect 262588 308440 262640 308446
rect 262588 308382 262640 308388
rect 263060 308378 263088 310420
rect 263152 310406 263350 310434
rect 263048 308372 263100 308378
rect 263048 308314 263100 308320
rect 263152 308258 263180 310406
rect 262496 308236 262548 308242
rect 262496 308178 262548 308184
rect 262600 308230 263180 308258
rect 262496 306332 262548 306338
rect 262496 306274 262548 306280
rect 262508 155417 262536 306274
rect 262494 155408 262550 155417
rect 262494 155343 262550 155352
rect 262404 147008 262456 147014
rect 262404 146950 262456 146956
rect 262312 133272 262364 133278
rect 262312 133214 262364 133220
rect 262600 111110 262628 308230
rect 262864 308168 262916 308174
rect 262864 308110 262916 308116
rect 262588 111104 262640 111110
rect 262588 111046 262640 111052
rect 262876 8974 262904 308110
rect 263520 306338 263548 310420
rect 263718 310406 263916 310434
rect 263888 306610 263916 310406
rect 263876 306604 263928 306610
rect 263876 306546 263928 306552
rect 263980 306490 264008 310420
rect 263704 306462 264008 306490
rect 263508 306332 263560 306338
rect 263508 306274 263560 306280
rect 263600 306332 263652 306338
rect 263600 306274 263652 306280
rect 263612 108322 263640 306274
rect 263704 109750 263732 306462
rect 263876 306400 263928 306406
rect 263876 306342 263928 306348
rect 263784 306264 263836 306270
rect 263784 306206 263836 306212
rect 263796 130490 263824 306206
rect 263888 131782 263916 306342
rect 263968 306196 264020 306202
rect 263968 306138 264020 306144
rect 263980 148442 264008 306138
rect 264164 296714 264192 310420
rect 264244 308712 264296 308718
rect 264244 308654 264296 308660
rect 264072 296686 264192 296714
rect 264072 149802 264100 296686
rect 264060 149796 264112 149802
rect 264060 149738 264112 149744
rect 263968 148436 264020 148442
rect 263968 148378 264020 148384
rect 263876 131776 263928 131782
rect 263876 131718 263928 131724
rect 263784 130484 263836 130490
rect 263784 130426 263836 130432
rect 263692 109744 263744 109750
rect 263692 109686 263744 109692
rect 263600 108316 263652 108322
rect 263600 108258 263652 108264
rect 264256 13190 264284 308654
rect 264348 306270 264376 310420
rect 264440 310406 264638 310434
rect 264440 306338 264468 310406
rect 264428 306332 264480 306338
rect 264428 306274 264480 306280
rect 264336 306264 264388 306270
rect 264336 306206 264388 306212
rect 264808 306202 264836 310420
rect 265006 310406 265112 310434
rect 264980 306264 265032 306270
rect 264980 306206 265032 306212
rect 264796 306196 264848 306202
rect 264796 306138 264848 306144
rect 264336 148368 264388 148374
rect 264336 148310 264388 148316
rect 264244 13184 264296 13190
rect 264244 13126 264296 13132
rect 262864 8968 262916 8974
rect 262864 8910 262916 8916
rect 264152 4820 264204 4826
rect 264152 4762 264204 4768
rect 261484 3868 261536 3874
rect 261484 3810 261536 3816
rect 260024 3454 260696 3482
rect 261404 3454 261800 3482
rect 260668 480 260696 3454
rect 261772 480 261800 3454
rect 262956 3324 263008 3330
rect 262956 3266 263008 3272
rect 262968 480 262996 3266
rect 264164 480 264192 4762
rect 264348 3806 264376 148310
rect 264428 108316 264480 108322
rect 264428 108258 264480 108264
rect 264336 3800 264388 3806
rect 264336 3742 264388 3748
rect 264440 3330 264468 108258
rect 264992 18630 265020 306206
rect 265084 129130 265112 310406
rect 265176 310406 265282 310434
rect 265176 131850 265204 310406
rect 265348 306400 265400 306406
rect 265348 306342 265400 306348
rect 265256 306332 265308 306338
rect 265256 306274 265308 306280
rect 265268 142934 265296 306274
rect 265360 145654 265388 306342
rect 265452 154018 265480 310420
rect 265544 310406 265742 310434
rect 265544 306338 265572 310406
rect 265624 307828 265676 307834
rect 265624 307770 265676 307776
rect 265532 306332 265584 306338
rect 265532 306274 265584 306280
rect 265636 159361 265664 307770
rect 265912 306270 265940 310420
rect 266096 306406 266124 310420
rect 266372 306814 266400 310420
rect 266556 309134 266584 310420
rect 266464 309106 266584 309134
rect 266360 306808 266412 306814
rect 266360 306750 266412 306756
rect 266084 306400 266136 306406
rect 266084 306342 266136 306348
rect 265900 306264 265952 306270
rect 265900 306206 265952 306212
rect 265622 159352 265678 159361
rect 265622 159287 265678 159296
rect 265440 154012 265492 154018
rect 265440 153954 265492 153960
rect 265624 153876 265676 153882
rect 265624 153818 265676 153824
rect 265348 145648 265400 145654
rect 265348 145590 265400 145596
rect 265256 142928 265308 142934
rect 265256 142870 265308 142876
rect 265348 142860 265400 142866
rect 265348 142802 265400 142808
rect 265164 131844 265216 131850
rect 265164 131786 265216 131792
rect 265072 129124 265124 129130
rect 265072 129066 265124 129072
rect 264980 18624 265032 18630
rect 264980 18566 265032 18572
rect 264428 3324 264480 3330
rect 264428 3266 264480 3272
rect 265360 480 265388 142802
rect 265636 3398 265664 153818
rect 266464 105602 266492 309106
rect 266740 307834 266768 310420
rect 266832 310406 267030 310434
rect 266728 307828 266780 307834
rect 266728 307770 266780 307776
rect 266636 306808 266688 306814
rect 266636 306750 266688 306756
rect 266544 306196 266596 306202
rect 266544 306138 266596 306144
rect 266556 127702 266584 306138
rect 266648 140146 266676 306750
rect 266832 306354 266860 310406
rect 266740 306326 266860 306354
rect 266740 148510 266768 306326
rect 266820 306264 266872 306270
rect 266820 306206 266872 306212
rect 266832 156913 266860 306206
rect 267200 296714 267228 310420
rect 267384 306270 267412 310420
rect 267476 310406 267674 310434
rect 267372 306264 267424 306270
rect 267372 306206 267424 306212
rect 267476 306202 267504 310406
rect 267844 306354 267872 310420
rect 268042 310406 268240 310434
rect 268108 306400 268160 306406
rect 267844 306326 267964 306354
rect 268108 306342 268160 306348
rect 267740 306264 267792 306270
rect 267740 306206 267792 306212
rect 267464 306196 267516 306202
rect 267464 306138 267516 306144
rect 266924 296686 267228 296714
rect 266818 156904 266874 156913
rect 266818 156839 266874 156848
rect 266728 148504 266780 148510
rect 266728 148446 266780 148452
rect 266636 140140 266688 140146
rect 266636 140082 266688 140088
rect 266544 127696 266596 127702
rect 266544 127638 266596 127644
rect 266544 106956 266596 106962
rect 266544 106898 266596 106904
rect 266452 105596 266504 105602
rect 266452 105538 266504 105544
rect 265624 3392 265676 3398
rect 265624 3334 265676 3340
rect 266556 480 266584 106898
rect 266924 19990 266952 296686
rect 267752 104242 267780 306206
rect 267832 306196 267884 306202
rect 267832 306138 267884 306144
rect 267844 126342 267872 306138
rect 267936 130558 267964 306326
rect 268016 306332 268068 306338
rect 268016 306274 268068 306280
rect 268028 138854 268056 306274
rect 268120 151230 268148 306342
rect 268212 152658 268240 310406
rect 268304 306338 268332 310420
rect 268384 308780 268436 308786
rect 268384 308722 268436 308728
rect 268396 308174 268424 308722
rect 268384 308168 268436 308174
rect 268384 308110 268436 308116
rect 268292 306332 268344 306338
rect 268292 306274 268344 306280
rect 268488 306270 268516 310420
rect 268580 310406 268778 310434
rect 268580 306406 268608 310406
rect 268568 306400 268620 306406
rect 268568 306342 268620 306348
rect 268476 306264 268528 306270
rect 268476 306206 268528 306212
rect 268948 306202 268976 310420
rect 268936 306196 268988 306202
rect 268936 306138 268988 306144
rect 268476 303544 268528 303550
rect 268476 303486 268528 303492
rect 268384 303272 268436 303278
rect 268384 303214 268436 303220
rect 268396 152862 268424 303214
rect 268488 152930 268516 303486
rect 268568 303476 268620 303482
rect 268568 303418 268620 303424
rect 268580 152998 268608 303418
rect 268658 300520 268714 300529
rect 268658 300455 268714 300464
rect 268568 152992 268620 152998
rect 268568 152934 268620 152940
rect 268476 152924 268528 152930
rect 268476 152866 268528 152872
rect 268384 152856 268436 152862
rect 268384 152798 268436 152804
rect 268672 152794 268700 300455
rect 268660 152788 268712 152794
rect 268660 152730 268712 152736
rect 268200 152652 268252 152658
rect 268200 152594 268252 152600
rect 268108 151224 268160 151230
rect 268108 151166 268160 151172
rect 268200 151088 268252 151094
rect 268200 151030 268252 151036
rect 268016 138848 268068 138854
rect 268016 138790 268068 138796
rect 267924 130552 267976 130558
rect 267924 130494 267976 130500
rect 267832 126336 267884 126342
rect 267832 126278 267884 126284
rect 267924 126268 267976 126274
rect 267924 126210 267976 126216
rect 267740 104236 267792 104242
rect 267740 104178 267792 104184
rect 266912 19984 266964 19990
rect 266912 19926 266964 19932
rect 267936 3602 267964 126210
rect 268212 6914 268240 151030
rect 269132 21418 269160 310420
rect 269316 310406 269422 310434
rect 269212 306332 269264 306338
rect 269212 306274 269264 306280
rect 269224 102882 269252 306274
rect 269316 305046 269344 310406
rect 269592 306354 269620 310420
rect 269408 306326 269620 306354
rect 269304 305040 269356 305046
rect 269304 304982 269356 304988
rect 269304 302388 269356 302394
rect 269304 302330 269356 302336
rect 269316 124982 269344 302330
rect 269408 137426 269436 306326
rect 269776 305266 269804 310420
rect 269500 305238 269804 305266
rect 269868 310406 270066 310434
rect 269500 147082 269528 305238
rect 269868 305130 269896 310406
rect 269592 305102 269896 305130
rect 269592 149870 269620 305102
rect 269672 305040 269724 305046
rect 269672 304982 269724 304988
rect 269684 159497 269712 304982
rect 270236 302394 270264 310420
rect 270420 306338 270448 310420
rect 270696 306474 270724 310420
rect 270684 306468 270736 306474
rect 270684 306410 270736 306416
rect 270500 306400 270552 306406
rect 270880 306354 270908 310420
rect 271064 310406 271170 310434
rect 270960 306468 271012 306474
rect 270960 306410 271012 306416
rect 270500 306342 270552 306348
rect 270408 306332 270460 306338
rect 270408 306274 270460 306280
rect 270224 302388 270276 302394
rect 270224 302330 270276 302336
rect 269670 159488 269726 159497
rect 269670 159423 269726 159432
rect 269762 150376 269818 150385
rect 269762 150311 269818 150320
rect 269580 149864 269632 149870
rect 269580 149806 269632 149812
rect 269488 147076 269540 147082
rect 269488 147018 269540 147024
rect 269396 137420 269448 137426
rect 269396 137362 269448 137368
rect 269304 124976 269356 124982
rect 269304 124918 269356 124924
rect 269212 102876 269264 102882
rect 269212 102818 269264 102824
rect 269120 21412 269172 21418
rect 269120 21354 269172 21360
rect 268028 6886 268240 6914
rect 267924 3596 267976 3602
rect 267924 3538 267976 3544
rect 268028 3482 268056 6886
rect 269776 3738 269804 150311
rect 270512 7614 270540 306342
rect 270592 306332 270644 306338
rect 270592 306274 270644 306280
rect 270696 306326 270908 306354
rect 270604 123554 270632 306274
rect 270696 136066 270724 306326
rect 270776 306264 270828 306270
rect 270776 306206 270828 306212
rect 270788 141574 270816 306206
rect 270868 306196 270920 306202
rect 270868 306138 270920 306144
rect 270880 144362 270908 306138
rect 270972 155553 271000 306410
rect 271064 306270 271092 310406
rect 271144 307828 271196 307834
rect 271144 307770 271196 307776
rect 271052 306264 271104 306270
rect 271052 306206 271104 306212
rect 270958 155544 271014 155553
rect 270958 155479 271014 155488
rect 271156 154086 271184 307770
rect 271340 306202 271368 310420
rect 271524 306338 271552 310420
rect 271616 310406 271814 310434
rect 271616 306406 271644 310406
rect 271984 307834 272012 310420
rect 271972 307828 272024 307834
rect 271972 307770 272024 307776
rect 272168 307018 272196 310420
rect 272260 310406 272458 310434
rect 272156 307012 272208 307018
rect 272156 306954 272208 306960
rect 272064 306808 272116 306814
rect 272064 306750 272116 306756
rect 271604 306400 271656 306406
rect 271604 306342 271656 306348
rect 271512 306332 271564 306338
rect 271512 306274 271564 306280
rect 271328 306196 271380 306202
rect 271328 306138 271380 306144
rect 271972 304292 272024 304298
rect 271972 304234 272024 304240
rect 271236 302864 271288 302870
rect 271236 302806 271288 302812
rect 271144 154080 271196 154086
rect 271144 154022 271196 154028
rect 271248 153066 271276 302806
rect 271420 302796 271472 302802
rect 271420 302738 271472 302744
rect 271328 302728 271380 302734
rect 271328 302670 271380 302676
rect 271340 153202 271368 302670
rect 271328 153196 271380 153202
rect 271328 153138 271380 153144
rect 271432 153134 271460 302738
rect 271420 153128 271472 153134
rect 271420 153070 271472 153076
rect 271236 153060 271288 153066
rect 271236 153002 271288 153008
rect 270868 144356 270920 144362
rect 270868 144298 270920 144304
rect 271144 143812 271196 143818
rect 271144 143754 271196 143760
rect 270776 141568 270828 141574
rect 270776 141510 270828 141516
rect 270684 136060 270736 136066
rect 270684 136002 270736 136008
rect 270592 123548 270644 123554
rect 270592 123490 270644 123496
rect 270776 10532 270828 10538
rect 270776 10474 270828 10480
rect 270500 7608 270552 7614
rect 270500 7550 270552 7556
rect 269764 3732 269816 3738
rect 269764 3674 269816 3680
rect 268476 3596 268528 3602
rect 268476 3538 268528 3544
rect 267752 3454 268056 3482
rect 267752 480 267780 3454
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 3538
rect 270040 3528 270092 3534
rect 270040 3470 270092 3476
rect 270052 480 270080 3470
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 10474
rect 271156 3602 271184 143754
rect 271236 135992 271288 135998
rect 271236 135934 271288 135940
rect 271144 3596 271196 3602
rect 271144 3538 271196 3544
rect 271248 3534 271276 135934
rect 271984 129198 272012 304234
rect 272076 145722 272104 306750
rect 272156 306264 272208 306270
rect 272156 306206 272208 306212
rect 272168 155038 272196 306206
rect 272260 304298 272288 310406
rect 272248 304292 272300 304298
rect 272248 304234 272300 304240
rect 272628 302234 272656 310420
rect 272812 306270 272840 310420
rect 272904 310406 273102 310434
rect 272800 306264 272852 306270
rect 272800 306206 272852 306212
rect 272260 302206 272656 302234
rect 272260 156466 272288 302206
rect 272904 296714 272932 310406
rect 273272 306202 273300 310420
rect 273470 310406 273576 310434
rect 273444 306672 273496 306678
rect 273444 306614 273496 306620
rect 273352 306400 273404 306406
rect 273352 306342 273404 306348
rect 273260 306196 273312 306202
rect 273260 306138 273312 306144
rect 273260 306060 273312 306066
rect 273260 306002 273312 306008
rect 272352 296686 272932 296714
rect 272248 156460 272300 156466
rect 272248 156402 272300 156408
rect 272156 155032 272208 155038
rect 272156 154974 272208 154980
rect 272064 145716 272116 145722
rect 272064 145658 272116 145664
rect 271972 129192 272024 129198
rect 271972 129134 272024 129140
rect 272352 122194 272380 296686
rect 272340 122188 272392 122194
rect 272340 122130 272392 122136
rect 273272 7682 273300 306002
rect 273364 9042 273392 306342
rect 273456 10402 273484 306614
rect 273548 306490 273576 310406
rect 273640 310406 273746 310434
rect 273640 306678 273668 310406
rect 273628 306672 273680 306678
rect 273628 306614 273680 306620
rect 273548 306462 273760 306490
rect 273536 306332 273588 306338
rect 273536 306274 273588 306280
rect 273548 15910 273576 306274
rect 273628 306264 273680 306270
rect 273628 306206 273680 306212
rect 273640 146946 273668 306206
rect 273732 152726 273760 306462
rect 273916 306270 273944 310420
rect 274008 310406 274206 310434
rect 273904 306264 273956 306270
rect 273904 306206 273956 306212
rect 273812 306196 273864 306202
rect 273812 306138 273864 306144
rect 273824 159390 273852 306138
rect 274008 306066 274036 310406
rect 274376 306406 274404 310420
rect 274364 306400 274416 306406
rect 274364 306342 274416 306348
rect 274560 306338 274588 310420
rect 274744 310406 274850 310434
rect 274548 306332 274600 306338
rect 274548 306274 274600 306280
rect 274744 306202 274772 310406
rect 274824 308304 274876 308310
rect 274824 308246 274876 308252
rect 274836 307086 274864 308246
rect 274824 307080 274876 307086
rect 274824 307022 274876 307028
rect 275020 306490 275048 310420
rect 274836 306462 275048 306490
rect 274732 306196 274784 306202
rect 274732 306138 274784 306144
rect 273996 306060 274048 306066
rect 273996 306002 274048 306008
rect 274732 306060 274784 306066
rect 274732 306002 274784 306008
rect 273994 303512 274050 303521
rect 273994 303447 274050 303456
rect 273904 302932 273956 302938
rect 273904 302874 273956 302880
rect 273812 159384 273864 159390
rect 273812 159326 273864 159332
rect 273916 155106 273944 302874
rect 274008 157321 274036 303447
rect 274088 303000 274140 303006
rect 274088 302942 274140 302948
rect 274100 159118 274128 302942
rect 274088 159112 274140 159118
rect 274088 159054 274140 159060
rect 274638 158264 274694 158273
rect 274638 158199 274694 158208
rect 274652 158098 274680 158199
rect 274640 158092 274692 158098
rect 274640 158034 274692 158040
rect 273994 157312 274050 157321
rect 273994 157247 274050 157256
rect 273904 155100 273956 155106
rect 273904 155042 273956 155048
rect 273720 152720 273772 152726
rect 273720 152662 273772 152668
rect 273628 146940 273680 146946
rect 273628 146882 273680 146888
rect 273536 15904 273588 15910
rect 273536 15846 273588 15852
rect 273904 14000 273956 14006
rect 273904 13942 273956 13948
rect 273444 10396 273496 10402
rect 273444 10338 273496 10344
rect 273352 9036 273404 9042
rect 273352 8978 273404 8984
rect 273260 7676 273312 7682
rect 273260 7618 273312 7624
rect 273628 4004 273680 4010
rect 273628 3946 273680 3952
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 272444 480 272472 3470
rect 273640 480 273668 3946
rect 273916 3534 273944 13942
rect 274744 6254 274772 306002
rect 274836 120766 274864 306462
rect 274916 306332 274968 306338
rect 275204 306320 275232 310420
rect 274916 306274 274968 306280
rect 275020 306292 275232 306320
rect 275296 310406 275494 310434
rect 274928 148374 274956 306274
rect 275020 153882 275048 306292
rect 275192 306196 275244 306202
rect 275192 306138 275244 306144
rect 275008 153876 275060 153882
rect 275008 153818 275060 153824
rect 275100 153876 275152 153882
rect 275100 153818 275152 153824
rect 274916 148368 274968 148374
rect 274916 148310 274968 148316
rect 274824 120760 274876 120766
rect 274824 120702 274876 120708
rect 274732 6248 274784 6254
rect 274732 6190 274784 6196
rect 273904 3528 273956 3534
rect 273904 3470 273956 3476
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 354 274906 480
rect 275112 354 275140 153818
rect 275204 4894 275232 306138
rect 275296 306066 275324 310406
rect 275664 308786 275692 310420
rect 275652 308780 275704 308786
rect 275652 308722 275704 308728
rect 275376 307828 275428 307834
rect 275376 307770 275428 307776
rect 275284 306060 275336 306066
rect 275284 306002 275336 306008
rect 275388 296714 275416 307770
rect 275848 306338 275876 310420
rect 275836 306332 275888 306338
rect 275836 306274 275888 306280
rect 275928 306264 275980 306270
rect 275928 306206 275980 306212
rect 275296 296686 275416 296714
rect 275296 17270 275324 296686
rect 275940 158273 275968 306206
rect 276020 158636 276072 158642
rect 276020 158578 276072 158584
rect 276032 158409 276060 158578
rect 276018 158400 276074 158409
rect 276018 158335 276074 158344
rect 275926 158264 275982 158273
rect 275926 158199 275982 158208
rect 276124 134570 276152 310420
rect 276308 308310 276336 310420
rect 276400 310406 276598 310434
rect 276296 308304 276348 308310
rect 276296 308246 276348 308252
rect 276400 306320 276428 310406
rect 276664 307964 276716 307970
rect 276664 307906 276716 307912
rect 276216 306292 276428 306320
rect 276216 143818 276244 306292
rect 276296 306196 276348 306202
rect 276296 306138 276348 306144
rect 276204 143812 276256 143818
rect 276204 143754 276256 143760
rect 276112 134564 276164 134570
rect 276112 134506 276164 134512
rect 275284 17264 275336 17270
rect 275284 17206 275336 17212
rect 276020 7608 276072 7614
rect 276020 7550 276072 7556
rect 275192 4888 275244 4894
rect 275192 4830 275244 4836
rect 276032 480 276060 7550
rect 276308 6186 276336 306138
rect 276676 106962 276704 307906
rect 276768 307834 276796 310420
rect 276952 308718 276980 310420
rect 277044 310406 277242 310434
rect 276940 308712 276992 308718
rect 276940 308654 276992 308660
rect 276756 307828 276808 307834
rect 276756 307770 276808 307776
rect 277044 306202 277072 310406
rect 277412 307873 277440 310420
rect 277596 308009 277624 310420
rect 277688 310406 277886 310434
rect 277582 308000 277638 308009
rect 277582 307935 277638 307944
rect 277398 307864 277454 307873
rect 277124 307828 277176 307834
rect 277398 307799 277454 307808
rect 277124 307770 277176 307776
rect 277032 306196 277084 306202
rect 277032 306138 277084 306144
rect 276940 303204 276992 303210
rect 276940 303146 276992 303152
rect 276848 303136 276900 303142
rect 276848 303078 276900 303084
rect 276756 303068 276808 303074
rect 276756 303010 276808 303016
rect 276768 155174 276796 303010
rect 276860 155242 276888 303078
rect 276952 156534 276980 303146
rect 277136 296714 277164 307770
rect 277688 306592 277716 310406
rect 278056 307834 278084 310420
rect 278136 307896 278188 307902
rect 278136 307838 278188 307844
rect 278044 307828 278096 307834
rect 278044 307770 278096 307776
rect 277504 306564 277716 306592
rect 277308 306060 277360 306066
rect 277308 306002 277360 306008
rect 277216 297900 277268 297906
rect 277216 297842 277268 297848
rect 277044 296686 277164 296714
rect 277044 162178 277072 296686
rect 277032 162172 277084 162178
rect 277032 162114 277084 162120
rect 277228 158030 277256 297842
rect 277320 158409 277348 306002
rect 277306 158400 277362 158409
rect 277306 158335 277362 158344
rect 277216 158024 277268 158030
rect 277216 157966 277268 157972
rect 276940 156528 276992 156534
rect 276940 156470 276992 156476
rect 276848 155236 276900 155242
rect 276848 155178 276900 155184
rect 276756 155168 276808 155174
rect 276756 155110 276808 155116
rect 276664 106956 276716 106962
rect 276664 106898 276716 106904
rect 277504 13122 277532 306564
rect 277584 306468 277636 306474
rect 277584 306410 277636 306416
rect 277596 108322 277624 306410
rect 277768 306332 277820 306338
rect 277768 306274 277820 306280
rect 277676 306196 277728 306202
rect 277676 306138 277728 306144
rect 277688 142866 277716 306138
rect 277676 142860 277728 142866
rect 277676 142802 277728 142808
rect 277584 108316 277636 108322
rect 277584 108258 277636 108264
rect 277492 13116 277544 13122
rect 277492 13058 277544 13064
rect 276296 6180 276348 6186
rect 276296 6122 276348 6128
rect 277780 4826 277808 306274
rect 278148 302234 278176 307838
rect 278240 306474 278268 310420
rect 278332 310406 278530 310434
rect 278228 306468 278280 306474
rect 278228 306410 278280 306416
rect 278332 306338 278360 310406
rect 278320 306332 278372 306338
rect 278320 306274 278372 306280
rect 278700 306202 278728 310420
rect 278780 308032 278832 308038
rect 278780 307974 278832 307980
rect 278688 306196 278740 306202
rect 278688 306138 278740 306144
rect 278688 305652 278740 305658
rect 278688 305594 278740 305600
rect 278056 302206 278176 302234
rect 278056 10538 278084 302206
rect 278594 300656 278650 300665
rect 278594 300591 278650 300600
rect 278412 300212 278464 300218
rect 278412 300154 278464 300160
rect 278320 297832 278372 297838
rect 278320 297774 278372 297780
rect 278332 158098 278360 297774
rect 278320 158092 278372 158098
rect 278320 158034 278372 158040
rect 278424 157146 278452 300154
rect 278504 300144 278556 300150
rect 278504 300086 278556 300092
rect 278136 157140 278188 157146
rect 278136 157082 278188 157088
rect 278412 157140 278464 157146
rect 278412 157082 278464 157088
rect 278148 156806 278176 157082
rect 278136 156800 278188 156806
rect 278136 156742 278188 156748
rect 278516 155718 278544 300086
rect 278504 155712 278556 155718
rect 278504 155654 278556 155660
rect 278608 154986 278636 300591
rect 278700 157894 278728 305594
rect 278688 157888 278740 157894
rect 278688 157830 278740 157836
rect 278700 157593 278728 157830
rect 278686 157584 278742 157593
rect 278686 157519 278742 157528
rect 278688 155712 278740 155718
rect 278688 155654 278740 155660
rect 278700 155106 278728 155654
rect 278688 155100 278740 155106
rect 278688 155042 278740 155048
rect 278608 154958 278728 154986
rect 278700 154562 278728 154958
rect 278688 154556 278740 154562
rect 278688 154498 278740 154504
rect 278700 154222 278728 154498
rect 278688 154216 278740 154222
rect 278688 154158 278740 154164
rect 278136 12504 278188 12510
rect 278136 12446 278188 12452
rect 278044 10532 278096 10538
rect 278044 10474 278096 10480
rect 277768 4820 277820 4826
rect 277768 4762 277820 4768
rect 278148 3194 278176 12446
rect 278792 6914 278820 307974
rect 278884 307970 278912 310420
rect 279068 310406 279174 310434
rect 278872 307964 278924 307970
rect 278872 307906 278924 307912
rect 278964 306400 279016 306406
rect 278964 306342 279016 306348
rect 278872 306332 278924 306338
rect 278872 306274 278924 306280
rect 278884 14006 278912 306274
rect 278976 126274 279004 306342
rect 279068 306134 279096 310406
rect 279344 306406 279372 310420
rect 279436 310406 279634 310434
rect 279332 306400 279384 306406
rect 279332 306342 279384 306348
rect 279436 306218 279464 310406
rect 279804 307902 279832 310420
rect 279792 307896 279844 307902
rect 279792 307838 279844 307844
rect 279516 307828 279568 307834
rect 279516 307770 279568 307776
rect 279252 306190 279464 306218
rect 279056 306128 279108 306134
rect 279056 306070 279108 306076
rect 279252 304314 279280 306190
rect 279332 306128 279384 306134
rect 279528 306082 279556 307770
rect 279988 306338 280016 310420
rect 279976 306332 280028 306338
rect 280264 306320 280292 310420
rect 280264 306292 280384 306320
rect 279976 306274 280028 306280
rect 280252 306196 280304 306202
rect 280252 306138 280304 306144
rect 279332 306070 279384 306076
rect 279068 304286 279280 304314
rect 279068 135998 279096 304286
rect 279344 299474 279372 306070
rect 279160 299446 279372 299474
rect 279436 306054 279556 306082
rect 279160 151094 279188 299446
rect 279148 151088 279200 151094
rect 279148 151030 279200 151036
rect 279056 135992 279108 135998
rect 279056 135934 279108 135940
rect 278964 126268 279016 126274
rect 278964 126210 279016 126216
rect 278872 14000 278924 14006
rect 278872 13942 278924 13948
rect 278792 6886 279096 6914
rect 278320 5568 278372 5574
rect 278320 5510 278372 5516
rect 277124 3188 277176 3194
rect 277124 3130 277176 3136
rect 278136 3188 278188 3194
rect 278136 3130 278188 3136
rect 277136 480 277164 3130
rect 278332 480 278360 5510
rect 274794 326 275140 354
rect 274794 -960 274906 326
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 6886
rect 279436 5574 279464 306054
rect 279608 303408 279660 303414
rect 279608 303350 279660 303356
rect 279516 303340 279568 303346
rect 279516 303282 279568 303288
rect 279528 155310 279556 303282
rect 279620 157826 279648 303350
rect 280066 300792 280122 300801
rect 280066 300727 280122 300736
rect 279976 297696 280028 297702
rect 279976 297638 280028 297644
rect 279608 157820 279660 157826
rect 279608 157762 279660 157768
rect 279516 155304 279568 155310
rect 279516 155246 279568 155252
rect 279988 154154 280016 297638
rect 280080 155718 280108 300727
rect 280068 155712 280120 155718
rect 280068 155654 280120 155660
rect 280080 155582 280108 155654
rect 280068 155576 280120 155582
rect 280068 155518 280120 155524
rect 279976 154148 280028 154154
rect 279976 154090 280028 154096
rect 279516 135244 279568 135250
rect 279516 135186 279568 135192
rect 279424 5568 279476 5574
rect 279424 5510 279476 5516
rect 279528 4010 279556 135186
rect 280264 12510 280292 306138
rect 280356 135250 280384 306292
rect 280448 153882 280476 310420
rect 280632 296714 280660 310420
rect 280724 310406 280922 310434
rect 280724 306202 280752 310406
rect 281092 307834 281120 310420
rect 281172 308916 281224 308922
rect 281172 308858 281224 308864
rect 281080 307828 281132 307834
rect 281080 307770 281132 307776
rect 280712 306196 280764 306202
rect 280712 306138 280764 306144
rect 281080 305992 281132 305998
rect 281080 305934 281132 305940
rect 280988 303612 281040 303618
rect 280988 303554 281040 303560
rect 280540 296686 280660 296714
rect 280436 153876 280488 153882
rect 280436 153818 280488 153824
rect 280344 135244 280396 135250
rect 280344 135186 280396 135192
rect 280252 12504 280304 12510
rect 280252 12446 280304 12452
rect 280540 7614 280568 296686
rect 280896 158636 280948 158642
rect 280896 158578 280948 158584
rect 280908 155378 280936 158578
rect 281000 157350 281028 303554
rect 280988 157344 281040 157350
rect 280988 157286 281040 157292
rect 281092 155786 281120 305934
rect 281184 305810 281212 308858
rect 281276 308038 281304 310420
rect 281448 309052 281500 309058
rect 281448 308994 281500 309000
rect 281356 308984 281408 308990
rect 281356 308926 281408 308932
rect 281264 308032 281316 308038
rect 281264 307974 281316 307980
rect 281184 305782 281304 305810
rect 281172 305720 281224 305726
rect 281172 305662 281224 305668
rect 281184 158642 281212 305662
rect 281172 158636 281224 158642
rect 281172 158578 281224 158584
rect 281172 157344 281224 157350
rect 281172 157286 281224 157292
rect 281184 156738 281212 157286
rect 281276 156806 281304 305782
rect 281368 156942 281396 308926
rect 281460 157010 281488 308994
rect 281552 306474 281580 310420
rect 281540 306468 281592 306474
rect 281540 306410 281592 306416
rect 281736 306320 281764 310420
rect 281552 306292 281764 306320
rect 281828 310406 282026 310434
rect 281448 157004 281500 157010
rect 281448 156946 281500 156952
rect 281356 156936 281408 156942
rect 281356 156878 281408 156884
rect 281264 156800 281316 156806
rect 281264 156742 281316 156748
rect 281172 156732 281224 156738
rect 281172 156674 281224 156680
rect 281080 155780 281132 155786
rect 281080 155722 281132 155728
rect 281448 155780 281500 155786
rect 281448 155722 281500 155728
rect 281460 155514 281488 155722
rect 281448 155508 281500 155514
rect 281448 155450 281500 155456
rect 280896 155372 280948 155378
rect 280896 155314 280948 155320
rect 280712 12504 280764 12510
rect 280712 12446 280764 12452
rect 280528 7608 280580 7614
rect 280528 7550 280580 7556
rect 279516 4004 279568 4010
rect 279516 3946 279568 3952
rect 280724 480 280752 12446
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 306292
rect 281632 306196 281684 306202
rect 281632 306138 281684 306144
rect 281644 3194 281672 306138
rect 281724 306128 281776 306134
rect 281724 306070 281776 306076
rect 281736 4214 281764 306070
rect 281828 8294 281856 310406
rect 281908 306468 281960 306474
rect 281908 306410 281960 306416
rect 281920 12510 281948 306410
rect 282196 306202 282224 310420
rect 282184 306196 282236 306202
rect 282184 306138 282236 306144
rect 282380 306134 282408 310420
rect 282656 308106 282684 310420
rect 282736 308780 282788 308786
rect 282736 308722 282788 308728
rect 282644 308100 282696 308106
rect 282644 308042 282696 308048
rect 282368 306128 282420 306134
rect 282368 306070 282420 306076
rect 282368 305924 282420 305930
rect 282368 305866 282420 305872
rect 282276 305856 282328 305862
rect 282276 305798 282328 305804
rect 282184 305788 282236 305794
rect 282184 305730 282236 305736
rect 282196 156602 282224 305730
rect 282288 156670 282316 305798
rect 282380 158545 282408 305866
rect 282748 302234 282776 308722
rect 282840 307902 282868 310420
rect 282828 307896 282880 307902
rect 282828 307838 282880 307844
rect 283024 306610 283052 310420
rect 283116 310406 283314 310434
rect 283012 306604 283064 306610
rect 283012 306546 283064 306552
rect 283116 306490 283144 310406
rect 282932 306462 283144 306490
rect 282748 302206 282868 302234
rect 282736 300280 282788 300286
rect 282736 300222 282788 300228
rect 282366 158536 282422 158545
rect 282366 158471 282422 158480
rect 282276 156664 282328 156670
rect 282276 156606 282328 156612
rect 282184 156596 282236 156602
rect 282184 156538 282236 156544
rect 282368 155780 282420 155786
rect 282368 155722 282420 155728
rect 282380 155446 282408 155722
rect 282748 155650 282776 300222
rect 282840 155786 282868 302206
rect 282828 155780 282880 155786
rect 282828 155722 282880 155728
rect 282736 155644 282788 155650
rect 282736 155586 282788 155592
rect 282368 155440 282420 155446
rect 282368 155382 282420 155388
rect 281908 12504 281960 12510
rect 281908 12446 281960 12452
rect 281816 8288 281868 8294
rect 281816 8230 281868 8236
rect 282932 4826 282960 306462
rect 283484 306354 283512 310420
rect 283564 308100 283616 308106
rect 283564 308042 283616 308048
rect 283012 306332 283064 306338
rect 283012 306274 283064 306280
rect 283208 306326 283512 306354
rect 283024 7002 283052 306274
rect 283104 306264 283156 306270
rect 283104 306206 283156 306212
rect 283116 9178 283144 306206
rect 283208 138854 283236 306326
rect 283288 306264 283340 306270
rect 283288 306206 283340 306212
rect 283300 149938 283328 306206
rect 283576 155854 283604 308042
rect 283668 306338 283696 310420
rect 283760 310406 283958 310434
rect 283656 306332 283708 306338
rect 283656 306274 283708 306280
rect 283760 306270 283788 310406
rect 283932 308644 283984 308650
rect 283932 308586 283984 308592
rect 283748 306264 283800 306270
rect 283748 306206 283800 306212
rect 283944 305182 283972 308586
rect 284128 307834 284156 310420
rect 284208 308372 284260 308378
rect 284208 308314 284260 308320
rect 284116 307828 284168 307834
rect 284116 307770 284168 307776
rect 284024 305516 284076 305522
rect 284024 305458 284076 305464
rect 283932 305176 283984 305182
rect 283932 305118 283984 305124
rect 283932 300552 283984 300558
rect 283932 300494 283984 300500
rect 283564 155848 283616 155854
rect 283564 155790 283616 155796
rect 283380 155576 283432 155582
rect 283380 155518 283432 155524
rect 283392 154970 283420 155518
rect 283472 155440 283524 155446
rect 283472 155382 283524 155388
rect 283380 154964 283432 154970
rect 283380 154906 283432 154912
rect 283484 154902 283512 155382
rect 283472 154896 283524 154902
rect 283472 154838 283524 154844
rect 283944 153814 283972 300494
rect 284036 155446 284064 305458
rect 284220 305266 284248 308314
rect 284312 307086 284340 310420
rect 284496 310406 284602 310434
rect 284300 307080 284352 307086
rect 284300 307022 284352 307028
rect 284392 306400 284444 306406
rect 284392 306342 284444 306348
rect 284300 306332 284352 306338
rect 284300 306274 284352 306280
rect 284128 305238 284248 305266
rect 284128 156398 284156 305238
rect 284208 305176 284260 305182
rect 284208 305118 284260 305124
rect 284116 156392 284168 156398
rect 284116 156334 284168 156340
rect 284220 155582 284248 305118
rect 284208 155576 284260 155582
rect 284208 155518 284260 155524
rect 284024 155440 284076 155446
rect 284024 155382 284076 155388
rect 283932 153808 283984 153814
rect 283932 153750 283984 153756
rect 283288 149932 283340 149938
rect 283288 149874 283340 149880
rect 283196 138848 283248 138854
rect 283196 138790 283248 138796
rect 283104 9172 283156 9178
rect 283104 9114 283156 9120
rect 283104 8288 283156 8294
rect 283104 8230 283156 8236
rect 283012 6996 283064 7002
rect 283012 6938 283064 6944
rect 282920 4820 282972 4826
rect 282920 4762 282972 4768
rect 281724 4208 281776 4214
rect 281724 4150 281776 4156
rect 281632 3188 281684 3194
rect 281632 3130 281684 3136
rect 283116 480 283144 8230
rect 284312 5234 284340 306274
rect 284404 152658 284432 306342
rect 284496 156942 284524 310406
rect 284772 306338 284800 310420
rect 285048 307834 285076 310420
rect 285128 307896 285180 307902
rect 285128 307838 285180 307844
rect 284944 307828 284996 307834
rect 284944 307770 284996 307776
rect 285036 307828 285088 307834
rect 285036 307770 285088 307776
rect 284760 306332 284812 306338
rect 284760 306274 284812 306280
rect 284852 297764 284904 297770
rect 284852 297706 284904 297712
rect 284760 247648 284812 247654
rect 284760 247590 284812 247596
rect 284772 247081 284800 247590
rect 284758 247072 284814 247081
rect 284758 247007 284814 247016
rect 284864 158545 284892 297706
rect 284666 158536 284722 158545
rect 284666 158471 284722 158480
rect 284850 158536 284906 158545
rect 284850 158471 284906 158480
rect 284576 158160 284628 158166
rect 284574 158128 284576 158137
rect 284628 158128 284630 158137
rect 284574 158063 284630 158072
rect 284680 157962 284708 158471
rect 284668 157956 284720 157962
rect 284668 157898 284720 157904
rect 284484 156936 284536 156942
rect 284484 156878 284536 156884
rect 284392 152652 284444 152658
rect 284392 152594 284444 152600
rect 284956 6458 284984 307770
rect 285140 302234 285168 307838
rect 285232 306406 285260 310420
rect 285416 307873 285444 310420
rect 285496 308304 285548 308310
rect 285496 308246 285548 308252
rect 285402 307864 285458 307873
rect 285402 307799 285458 307808
rect 285220 306400 285272 306406
rect 285220 306342 285272 306348
rect 285048 302206 285168 302234
rect 285048 144090 285076 302206
rect 285312 300348 285364 300354
rect 285312 300290 285364 300296
rect 285128 300008 285180 300014
rect 285128 299950 285180 299956
rect 285140 171086 285168 299950
rect 285220 243636 285272 243642
rect 285220 243578 285272 243584
rect 285128 171080 285180 171086
rect 285128 171022 285180 171028
rect 285140 170406 285168 171022
rect 285128 170400 285180 170406
rect 285128 170342 285180 170348
rect 285232 158982 285260 243578
rect 285220 158976 285272 158982
rect 285220 158918 285272 158924
rect 285324 158137 285352 300290
rect 285402 158808 285458 158817
rect 285402 158743 285458 158752
rect 285310 158128 285366 158137
rect 285310 158063 285366 158072
rect 285036 144084 285088 144090
rect 285036 144026 285088 144032
rect 285416 9042 285444 158743
rect 285508 156330 285536 308246
rect 285692 306374 285720 310420
rect 285876 306626 285904 310420
rect 286060 307902 286088 310420
rect 286152 310406 286350 310434
rect 286048 307896 286100 307902
rect 286048 307838 286100 307844
rect 285876 306598 286088 306626
rect 285692 306346 285996 306374
rect 285772 306264 285824 306270
rect 285772 306206 285824 306212
rect 285680 305244 285732 305250
rect 285680 305186 285732 305192
rect 285588 247920 285640 247926
rect 285588 247862 285640 247868
rect 285600 247217 285628 247862
rect 285586 247208 285642 247217
rect 285586 247143 285642 247152
rect 285586 169824 285642 169833
rect 285586 169759 285642 169768
rect 285496 156324 285548 156330
rect 285496 156266 285548 156272
rect 285404 9036 285456 9042
rect 285404 8978 285456 8984
rect 284944 6452 284996 6458
rect 284944 6394 284996 6400
rect 284300 5228 284352 5234
rect 284300 5170 284352 5176
rect 285404 4208 285456 4214
rect 285404 4150 285456 4156
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 284312 480 284340 3130
rect 285416 480 285444 4150
rect 285600 3466 285628 169759
rect 285588 3460 285640 3466
rect 285588 3402 285640 3408
rect 285692 3398 285720 305186
rect 285784 5166 285812 306206
rect 285968 302234 285996 306346
rect 285876 302206 285996 302234
rect 285876 297498 285904 302206
rect 285864 297492 285916 297498
rect 285864 297434 285916 297440
rect 286060 297378 286088 306598
rect 285876 297350 286088 297378
rect 285876 147082 285904 297350
rect 285956 297288 286008 297294
rect 285956 297230 286008 297236
rect 285968 156738 285996 297230
rect 286152 292574 286180 310406
rect 286324 307828 286376 307834
rect 286324 307770 286376 307776
rect 286060 292546 286180 292574
rect 285956 156732 286008 156738
rect 285956 156674 286008 156680
rect 285956 155848 286008 155854
rect 285956 155790 286008 155796
rect 285864 147076 285916 147082
rect 285864 147018 285916 147024
rect 285968 16574 285996 155790
rect 286060 155174 286088 292546
rect 286336 159594 286364 307770
rect 286520 306270 286548 310420
rect 286508 306264 286560 306270
rect 286508 306206 286560 306212
rect 286704 305250 286732 310420
rect 286980 307873 287008 310420
rect 287178 310406 287376 310434
rect 286966 307864 287022 307873
rect 286966 307799 287022 307808
rect 287244 306400 287296 306406
rect 287244 306342 287296 306348
rect 287152 306332 287204 306338
rect 287152 306274 287204 306280
rect 286692 305244 286744 305250
rect 286692 305186 286744 305192
rect 287060 304292 287112 304298
rect 287060 304234 287112 304240
rect 286784 300688 286836 300694
rect 286784 300630 286836 300636
rect 286600 300484 286652 300490
rect 286600 300426 286652 300432
rect 286324 159588 286376 159594
rect 286324 159530 286376 159536
rect 286140 158704 286192 158710
rect 286140 158646 286192 158652
rect 286152 158166 286180 158646
rect 286612 158370 286640 300426
rect 286692 247512 286744 247518
rect 286692 247454 286744 247460
rect 286704 247081 286732 247454
rect 286690 247072 286746 247081
rect 286690 247007 286746 247016
rect 286692 243568 286744 243574
rect 286692 243510 286744 243516
rect 286600 158364 286652 158370
rect 286600 158306 286652 158312
rect 286140 158160 286192 158166
rect 286140 158102 286192 158108
rect 286324 156936 286376 156942
rect 286324 156878 286376 156884
rect 286140 155780 286192 155786
rect 286140 155722 286192 155728
rect 286152 155378 286180 155722
rect 286140 155372 286192 155378
rect 286140 155314 286192 155320
rect 286048 155168 286100 155174
rect 286048 155110 286100 155116
rect 285968 16546 286272 16574
rect 285772 5160 285824 5166
rect 285772 5102 285824 5108
rect 286244 3482 286272 16546
rect 286336 3602 286364 156878
rect 286600 156800 286652 156806
rect 286600 156742 286652 156748
rect 286612 156330 286640 156742
rect 286600 156324 286652 156330
rect 286600 156266 286652 156272
rect 286704 154290 286732 243510
rect 286796 158166 286824 300630
rect 286876 300416 286928 300422
rect 286876 300358 286928 300364
rect 286784 158160 286836 158166
rect 286784 158102 286836 158108
rect 286888 157078 286916 300358
rect 286968 247580 287020 247586
rect 286968 247522 287020 247528
rect 286980 247081 287008 247522
rect 286966 247072 287022 247081
rect 286966 247007 287022 247016
rect 286966 158808 287022 158817
rect 286966 158743 287022 158752
rect 286876 157072 286928 157078
rect 286876 157014 286928 157020
rect 286692 154284 286744 154290
rect 286692 154226 286744 154232
rect 286980 6186 287008 158743
rect 287072 11762 287100 304234
rect 287164 13122 287192 306274
rect 287256 144294 287284 306342
rect 287348 145654 287376 310406
rect 287440 306338 287468 310420
rect 287428 306332 287480 306338
rect 287428 306274 287480 306280
rect 287428 306060 287480 306066
rect 287428 306002 287480 306008
rect 287440 156602 287468 306002
rect 287624 292574 287652 310420
rect 287704 309052 287756 309058
rect 287704 308994 287756 309000
rect 287532 292546 287652 292574
rect 287532 159526 287560 292546
rect 287520 159520 287572 159526
rect 287520 159462 287572 159468
rect 287716 158846 287744 308994
rect 287808 306406 287836 310420
rect 287900 310406 288098 310434
rect 287796 306400 287848 306406
rect 287796 306342 287848 306348
rect 287900 304298 287928 310406
rect 288268 306066 288296 310420
rect 288452 306338 288480 310420
rect 288544 310406 288742 310434
rect 288440 306332 288492 306338
rect 288440 306274 288492 306280
rect 288256 306060 288308 306066
rect 288256 306002 288308 306008
rect 288440 306060 288492 306066
rect 288440 306002 288492 306008
rect 287888 304292 287940 304298
rect 287888 304234 287940 304240
rect 288256 300076 288308 300082
rect 288256 300018 288308 300024
rect 288164 247988 288216 247994
rect 288164 247930 288216 247936
rect 287980 247852 288032 247858
rect 287980 247794 288032 247800
rect 287888 247784 287940 247790
rect 287888 247726 287940 247732
rect 287900 247081 287928 247726
rect 287992 247217 288020 247794
rect 287978 247208 288034 247217
rect 287978 247143 288034 247152
rect 287886 247072 287942 247081
rect 287886 247007 287942 247016
rect 288070 159080 288126 159089
rect 288070 159015 288126 159024
rect 287978 158944 288034 158953
rect 287978 158879 288034 158888
rect 287704 158840 287756 158846
rect 287704 158782 287756 158788
rect 287886 158808 287942 158817
rect 287886 158743 287942 158752
rect 287428 156596 287480 156602
rect 287428 156538 287480 156544
rect 287336 145648 287388 145654
rect 287336 145590 287388 145596
rect 287244 144288 287296 144294
rect 287244 144230 287296 144236
rect 287336 144084 287388 144090
rect 287336 144026 287388 144032
rect 287152 13116 287204 13122
rect 287152 13058 287204 13064
rect 287060 11756 287112 11762
rect 287060 11698 287112 11704
rect 286968 6180 287020 6186
rect 286968 6122 287020 6128
rect 286324 3596 286376 3602
rect 286324 3538 286376 3544
rect 286244 3454 286640 3482
rect 285680 3392 285732 3398
rect 285680 3334 285732 3340
rect 286612 480 286640 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 144026
rect 287900 6594 287928 158743
rect 287888 6588 287940 6594
rect 287888 6530 287940 6536
rect 287992 6390 288020 158879
rect 288084 8974 288112 159015
rect 288176 158846 288204 247930
rect 288164 158840 288216 158846
rect 288164 158782 288216 158788
rect 288268 158506 288296 300018
rect 288348 245132 288400 245138
rect 288348 245074 288400 245080
rect 288256 158500 288308 158506
rect 288256 158442 288308 158448
rect 288072 8968 288124 8974
rect 288072 8910 288124 8916
rect 287980 6384 288032 6390
rect 287980 6326 288032 6332
rect 288360 3806 288388 245074
rect 288452 17270 288480 306002
rect 288544 130422 288572 310406
rect 288912 307018 288940 310420
rect 288900 307012 288952 307018
rect 288900 306954 288952 306960
rect 288992 306808 289044 306814
rect 288992 306750 289044 306756
rect 288624 306400 288676 306406
rect 288624 306342 288676 306348
rect 288636 141438 288664 306342
rect 288808 306332 288860 306338
rect 288808 306274 288860 306280
rect 288716 301300 288768 301306
rect 288716 301242 288768 301248
rect 288728 142866 288756 301242
rect 288820 149870 288848 306274
rect 288900 306264 288952 306270
rect 288900 306206 288952 306212
rect 288912 155378 288940 306206
rect 289004 159458 289032 306750
rect 289096 301306 289124 310420
rect 289188 310406 289386 310434
rect 289188 306066 289216 310406
rect 289556 306270 289584 310420
rect 289740 306406 289768 310420
rect 289924 310406 290030 310434
rect 289820 306468 289872 306474
rect 289820 306410 289872 306416
rect 289728 306400 289780 306406
rect 289728 306342 289780 306348
rect 289544 306264 289596 306270
rect 289544 306206 289596 306212
rect 289176 306060 289228 306066
rect 289176 306002 289228 306008
rect 289084 301300 289136 301306
rect 289084 301242 289136 301248
rect 289544 300756 289596 300762
rect 289544 300698 289596 300704
rect 289452 300620 289504 300626
rect 289452 300562 289504 300568
rect 289360 248396 289412 248402
rect 289360 248338 289412 248344
rect 289176 247716 289228 247722
rect 289176 247658 289228 247664
rect 289188 247081 289216 247658
rect 289372 247217 289400 248338
rect 289358 247208 289414 247217
rect 289358 247143 289414 247152
rect 289174 247072 289230 247081
rect 289174 247007 289230 247016
rect 288992 159452 289044 159458
rect 288992 159394 289044 159400
rect 289358 158808 289414 158817
rect 289358 158743 289414 158752
rect 288900 155372 288952 155378
rect 288900 155314 288952 155320
rect 288808 149864 288860 149870
rect 288808 149806 288860 149812
rect 288716 142860 288768 142866
rect 288716 142802 288768 142808
rect 288624 141432 288676 141438
rect 288624 141374 288676 141380
rect 288532 130416 288584 130422
rect 288532 130358 288584 130364
rect 288440 17264 288492 17270
rect 288440 17206 288492 17212
rect 289372 9110 289400 158743
rect 289464 158438 289492 300562
rect 289556 158658 289584 300698
rect 289636 246560 289688 246566
rect 289636 246502 289688 246508
rect 289648 158778 289676 246502
rect 289726 158944 289782 158953
rect 289726 158879 289782 158888
rect 289636 158772 289688 158778
rect 289636 158714 289688 158720
rect 289556 158630 289676 158658
rect 289452 158432 289504 158438
rect 289452 158374 289504 158380
rect 289648 158302 289676 158630
rect 289636 158296 289688 158302
rect 289636 158238 289688 158244
rect 289648 158001 289676 158238
rect 289634 157992 289690 158001
rect 289634 157927 289690 157936
rect 289360 9104 289412 9110
rect 289360 9046 289412 9052
rect 288992 6996 289044 7002
rect 288992 6938 289044 6944
rect 288348 3800 288400 3806
rect 288348 3742 288400 3748
rect 289004 480 289032 6938
rect 289740 6526 289768 158879
rect 289832 15910 289860 306410
rect 289924 129062 289952 310406
rect 290200 309097 290228 310420
rect 290186 309088 290242 309097
rect 290186 309023 290242 309032
rect 290476 308961 290504 310420
rect 290556 309120 290608 309126
rect 290556 309062 290608 309068
rect 290462 308952 290518 308961
rect 290462 308887 290518 308896
rect 290096 306400 290148 306406
rect 290096 306342 290148 306348
rect 290004 306332 290056 306338
rect 290004 306274 290056 306280
rect 290016 145586 290044 306274
rect 290108 153882 290136 306342
rect 290568 292574 290596 309062
rect 290660 306474 290688 310420
rect 290648 306468 290700 306474
rect 290648 306410 290700 306416
rect 290844 306406 290872 310420
rect 290936 310406 291134 310434
rect 290832 306400 290884 306406
rect 290832 306342 290884 306348
rect 290936 306338 290964 310406
rect 291016 307964 291068 307970
rect 291016 307906 291068 307912
rect 290924 306332 290976 306338
rect 290924 306274 290976 306280
rect 291028 302234 291056 307906
rect 291304 306354 291332 310420
rect 291502 310406 291700 310434
rect 291672 306610 291700 310406
rect 291660 306604 291712 306610
rect 291660 306546 291712 306552
rect 291764 306490 291792 310420
rect 291844 307896 291896 307902
rect 291844 307838 291896 307844
rect 290476 292546 290596 292574
rect 290844 302206 291056 302234
rect 291212 306326 291332 306354
rect 291396 306462 291792 306490
rect 290476 159186 290504 292546
rect 290740 248056 290792 248062
rect 290740 247998 290792 248004
rect 290648 244724 290700 244730
rect 290648 244666 290700 244672
rect 290660 244361 290688 244666
rect 290646 244352 290702 244361
rect 290646 244287 290702 244296
rect 290464 159180 290516 159186
rect 290464 159122 290516 159128
rect 290752 159118 290780 247998
rect 290740 159112 290792 159118
rect 290740 159054 290792 159060
rect 290646 158808 290702 158817
rect 290646 158743 290702 158752
rect 290096 153876 290148 153882
rect 290096 153818 290148 153824
rect 290004 145580 290056 145586
rect 290004 145522 290056 145528
rect 289912 129056 289964 129062
rect 289912 128998 289964 129004
rect 289820 15904 289872 15910
rect 289820 15846 289872 15852
rect 289728 6520 289780 6526
rect 289728 6462 289780 6468
rect 290660 6322 290688 158743
rect 290844 157214 290872 302206
rect 290924 300824 290976 300830
rect 290924 300766 290976 300772
rect 290936 158710 290964 300766
rect 291108 244996 291160 245002
rect 291108 244938 291160 244944
rect 291016 244928 291068 244934
rect 291016 244870 291068 244876
rect 290924 158704 290976 158710
rect 290924 158646 290976 158652
rect 290832 157208 290884 157214
rect 290832 157150 290884 157156
rect 291028 6662 291056 244870
rect 291120 6730 291148 244938
rect 291212 127634 291240 306326
rect 291292 305584 291344 305590
rect 291292 305526 291344 305532
rect 291304 138718 291332 305526
rect 291396 140078 291424 306462
rect 291660 306332 291712 306338
rect 291660 306274 291712 306280
rect 291568 306264 291620 306270
rect 291568 306206 291620 306212
rect 291476 306060 291528 306066
rect 291476 306002 291528 306008
rect 291488 149802 291516 306002
rect 291580 151094 291608 306206
rect 291672 152590 291700 306274
rect 291752 245472 291804 245478
rect 291752 245414 291804 245420
rect 291764 244361 291792 245414
rect 291750 244352 291806 244361
rect 291750 244287 291806 244296
rect 291660 152584 291712 152590
rect 291660 152526 291712 152532
rect 291568 151088 291620 151094
rect 291568 151030 291620 151036
rect 291476 149796 291528 149802
rect 291476 149738 291528 149744
rect 291384 140072 291436 140078
rect 291384 140014 291436 140020
rect 291384 138848 291436 138854
rect 291384 138790 291436 138796
rect 291292 138712 291344 138718
rect 291292 138654 291344 138660
rect 291200 127628 291252 127634
rect 291200 127570 291252 127576
rect 291108 6724 291160 6730
rect 291108 6666 291160 6672
rect 291016 6656 291068 6662
rect 291016 6598 291068 6604
rect 290648 6316 290700 6322
rect 290648 6258 290700 6264
rect 290188 4820 290240 4826
rect 290188 4762 290240 4768
rect 290200 480 290228 4762
rect 291396 480 291424 138790
rect 291856 14482 291884 307838
rect 291948 306066 291976 310420
rect 292132 306270 292160 310420
rect 292224 310406 292422 310434
rect 292120 306264 292172 306270
rect 292120 306206 292172 306212
rect 291936 306060 291988 306066
rect 291936 306002 291988 306008
rect 292028 306060 292080 306066
rect 292028 306002 292080 306008
rect 292040 305522 292068 306002
rect 292224 305590 292252 310406
rect 292396 306264 292448 306270
rect 292396 306206 292448 306212
rect 292212 305584 292264 305590
rect 292212 305526 292264 305532
rect 292028 305516 292080 305522
rect 292028 305458 292080 305464
rect 292212 299940 292264 299946
rect 292212 299882 292264 299888
rect 292120 245608 292172 245614
rect 292120 245550 292172 245556
rect 292132 244361 292160 245550
rect 292118 244352 292174 244361
rect 292118 244287 292174 244296
rect 292224 158302 292252 299882
rect 292304 248192 292356 248198
rect 292304 248134 292356 248140
rect 292316 159254 292344 248134
rect 292304 159248 292356 159254
rect 292304 159190 292356 159196
rect 292212 158296 292264 158302
rect 292212 158238 292264 158244
rect 292408 157282 292436 306206
rect 292486 158808 292542 158817
rect 292486 158743 292542 158752
rect 292396 157276 292448 157282
rect 292396 157218 292448 157224
rect 291844 14476 291896 14482
rect 291844 14418 291896 14424
rect 292500 6254 292528 158743
rect 292592 126274 292620 310420
rect 292672 306332 292724 306338
rect 292672 306274 292724 306280
rect 292684 137290 292712 306274
rect 292868 305674 292896 310420
rect 292868 305646 292988 305674
rect 292856 305584 292908 305590
rect 292856 305526 292908 305532
rect 292764 302048 292816 302054
rect 292764 301990 292816 301996
rect 292776 144226 292804 301990
rect 292868 149734 292896 305526
rect 292960 155310 292988 305646
rect 293052 302054 293080 310420
rect 293236 307834 293264 310420
rect 293328 310406 293526 310434
rect 293224 307828 293276 307834
rect 293224 307770 293276 307776
rect 293224 307080 293276 307086
rect 293224 307022 293276 307028
rect 293040 302048 293092 302054
rect 293040 301990 293092 301996
rect 292948 155304 293000 155310
rect 292948 155246 293000 155252
rect 292948 149932 293000 149938
rect 292948 149874 293000 149880
rect 292856 149728 292908 149734
rect 292856 149670 292908 149676
rect 292764 144220 292816 144226
rect 292764 144162 292816 144168
rect 292672 137284 292724 137290
rect 292672 137226 292724 137232
rect 292580 126268 292632 126274
rect 292580 126210 292632 126216
rect 292960 12434 292988 149874
rect 293236 16574 293264 307022
rect 293328 305590 293356 310406
rect 293498 309088 293554 309097
rect 293498 309023 293554 309032
rect 293406 308952 293462 308961
rect 293406 308887 293462 308896
rect 293316 305584 293368 305590
rect 293316 305526 293368 305532
rect 293420 296714 293448 308887
rect 293328 296686 293448 296714
rect 293328 147014 293356 296686
rect 293408 245404 293460 245410
rect 293408 245346 293460 245352
rect 293420 244361 293448 245346
rect 293406 244352 293462 244361
rect 293406 244287 293462 244296
rect 293512 156670 293540 309023
rect 293696 306338 293724 310420
rect 293880 307873 293908 310420
rect 294064 310406 294170 310434
rect 293866 307864 293922 307873
rect 293866 307799 293922 307808
rect 293684 306332 293736 306338
rect 293684 306274 293736 306280
rect 293960 306332 294012 306338
rect 293960 306274 294012 306280
rect 293684 248124 293736 248130
rect 293684 248066 293736 248072
rect 293696 197334 293724 248066
rect 293776 245268 293828 245274
rect 293776 245210 293828 245216
rect 293788 244361 293816 245210
rect 293774 244352 293830 244361
rect 293774 244287 293830 244296
rect 293776 243772 293828 243778
rect 293776 243714 293828 243720
rect 293684 197328 293736 197334
rect 293684 197270 293736 197276
rect 293788 159186 293816 243714
rect 293866 196072 293922 196081
rect 293866 196007 293922 196016
rect 293776 159180 293828 159186
rect 293776 159122 293828 159128
rect 293500 156664 293552 156670
rect 293500 156606 293552 156612
rect 293316 147008 293368 147014
rect 293316 146950 293368 146956
rect 293236 16546 293356 16574
rect 292960 12406 293264 12434
rect 292580 9172 292632 9178
rect 292580 9114 292632 9120
rect 292488 6248 292540 6254
rect 292488 6190 292540 6196
rect 292592 480 292620 9114
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 12406
rect 293328 4146 293356 16546
rect 293316 4140 293368 4146
rect 293316 4082 293368 4088
rect 293880 3534 293908 196007
rect 293972 3942 294000 306274
rect 294064 4078 294092 310406
rect 294340 306354 294368 310420
rect 294156 306326 294368 306354
rect 294156 5098 294184 306326
rect 294236 305584 294288 305590
rect 294236 305526 294288 305532
rect 294144 5092 294196 5098
rect 294144 5034 294196 5040
rect 294248 5030 294276 305526
rect 294524 296714 294552 310420
rect 294616 310406 294814 310434
rect 294616 306338 294644 310406
rect 294696 307828 294748 307834
rect 294696 307770 294748 307776
rect 294604 306332 294656 306338
rect 294604 306274 294656 306280
rect 294708 302234 294736 307770
rect 294984 305590 295012 310420
rect 295168 307834 295196 310420
rect 295352 310406 295458 310434
rect 295642 310406 295840 310434
rect 295156 307828 295208 307834
rect 295156 307770 295208 307776
rect 294972 305584 295024 305590
rect 294972 305526 295024 305532
rect 294972 305312 295024 305318
rect 294972 305254 295024 305260
rect 294340 296686 294552 296714
rect 294616 302206 294736 302234
rect 294340 155242 294368 296686
rect 294328 155236 294380 155242
rect 294328 155178 294380 155184
rect 294616 152522 294644 302206
rect 294878 168464 294934 168473
rect 294878 168399 294934 168408
rect 294604 152516 294656 152522
rect 294604 152458 294656 152464
rect 294892 16574 294920 168399
rect 294984 158642 295012 305254
rect 295064 245336 295116 245342
rect 295064 245278 295116 245284
rect 295076 244361 295104 245278
rect 295248 245200 295300 245206
rect 295248 245142 295300 245148
rect 295156 245064 295208 245070
rect 295156 245006 295208 245012
rect 295062 244352 295118 244361
rect 295062 244287 295118 244296
rect 295064 243976 295116 243982
rect 295064 243918 295116 243924
rect 295076 169318 295104 243918
rect 295064 169312 295116 169318
rect 295064 169254 295116 169260
rect 294972 158636 295024 158642
rect 294972 158578 295024 158584
rect 294892 16546 295012 16574
rect 294984 6458 295012 16546
rect 294880 6452 294932 6458
rect 294880 6394 294932 6400
rect 294972 6452 295024 6458
rect 294972 6394 295024 6400
rect 294236 5024 294288 5030
rect 294236 4966 294288 4972
rect 294052 4072 294104 4078
rect 294052 4014 294104 4020
rect 293960 3936 294012 3942
rect 293960 3878 294012 3884
rect 293868 3528 293920 3534
rect 293868 3470 293920 3476
rect 294892 480 294920 6394
rect 295168 3670 295196 245006
rect 295260 3738 295288 245142
rect 295352 4010 295380 310406
rect 295616 306536 295668 306542
rect 295616 306478 295668 306484
rect 295432 306468 295484 306474
rect 295432 306410 295484 306416
rect 295340 4004 295392 4010
rect 295340 3946 295392 3952
rect 295444 3874 295472 306410
rect 295524 306332 295576 306338
rect 295524 306274 295576 306280
rect 295536 6798 295564 306274
rect 295628 18630 295656 306478
rect 295708 306400 295760 306406
rect 295708 306342 295760 306348
rect 295720 146946 295748 306342
rect 295812 148374 295840 310406
rect 295904 306338 295932 310420
rect 295982 307864 296038 307873
rect 295982 307799 296038 307808
rect 295892 306332 295944 306338
rect 295892 306274 295944 306280
rect 295892 158228 295944 158234
rect 295892 158170 295944 158176
rect 295904 157758 295932 158170
rect 295892 157752 295944 157758
rect 295892 157694 295944 157700
rect 295800 148368 295852 148374
rect 295800 148310 295852 148316
rect 295708 146940 295760 146946
rect 295708 146882 295760 146888
rect 295996 24138 296024 307799
rect 296088 306474 296116 310420
rect 296076 306468 296128 306474
rect 296076 306410 296128 306416
rect 296272 306406 296300 310420
rect 296364 310406 296562 310434
rect 296364 306542 296392 310406
rect 296732 309134 296760 310420
rect 296640 309106 296760 309134
rect 296444 307828 296496 307834
rect 296444 307770 296496 307776
rect 296352 306536 296404 306542
rect 296352 306478 296404 306484
rect 296260 306400 296312 306406
rect 296260 306342 296312 306348
rect 296456 305946 296484 307770
rect 296088 305918 296484 305946
rect 296088 124914 296116 305918
rect 296640 305386 296668 309106
rect 296916 305504 296944 310420
rect 297192 307873 297220 310420
rect 297178 307864 297234 307873
rect 297178 307799 297234 307808
rect 296732 305476 296944 305504
rect 296628 305380 296680 305386
rect 296628 305322 296680 305328
rect 296628 305244 296680 305250
rect 296628 305186 296680 305192
rect 296536 248260 296588 248266
rect 296536 248202 296588 248208
rect 296548 159390 296576 248202
rect 296536 159384 296588 159390
rect 296536 159326 296588 159332
rect 296640 158234 296668 305186
rect 296628 158228 296680 158234
rect 296628 158170 296680 158176
rect 296076 124908 296128 124914
rect 296076 124850 296128 124856
rect 295984 24132 296036 24138
rect 295984 24074 296036 24080
rect 295616 18624 295668 18630
rect 295616 18566 295668 18572
rect 295524 6792 295576 6798
rect 295524 6734 295576 6740
rect 296732 4962 296760 305476
rect 296812 305380 296864 305386
rect 296812 305322 296864 305328
rect 296824 245041 296852 305322
rect 297376 296714 297404 310420
rect 297560 308145 297588 310420
rect 297546 308136 297602 308145
rect 297546 308071 297602 308080
rect 297836 307873 297864 310420
rect 298020 308009 298048 310420
rect 298218 310406 298416 310434
rect 298006 308000 298062 308009
rect 298006 307935 298062 307944
rect 297822 307864 297878 307873
rect 297822 307799 297878 307808
rect 298284 306400 298336 306406
rect 298284 306342 298336 306348
rect 298388 306354 298416 310406
rect 298480 307873 298508 310420
rect 298466 307864 298522 307873
rect 298466 307799 298522 307808
rect 298192 306332 298244 306338
rect 298192 306274 298244 306280
rect 298008 298036 298060 298042
rect 298008 297978 298060 297984
rect 297916 297968 297968 297974
rect 297916 297910 297968 297916
rect 296916 296686 297404 296714
rect 296916 245138 296944 296686
rect 297548 254720 297600 254726
rect 297548 254662 297600 254668
rect 297180 253428 297232 253434
rect 297180 253370 297232 253376
rect 296904 245132 296956 245138
rect 296904 245074 296956 245080
rect 296810 245032 296866 245041
rect 296810 244967 296866 244976
rect 297086 245032 297142 245041
rect 297086 244967 297142 244976
rect 297100 244633 297128 244967
rect 297086 244624 297142 244633
rect 297086 244559 297142 244568
rect 297192 244390 297220 253370
rect 297456 252068 297508 252074
rect 297456 252010 297508 252016
rect 297272 246628 297324 246634
rect 297272 246570 297324 246576
rect 297180 244384 297232 244390
rect 297180 244326 297232 244332
rect 297180 197328 297232 197334
rect 297180 197270 297232 197276
rect 297192 158914 297220 197270
rect 297284 196450 297312 246570
rect 297364 244384 297416 244390
rect 297364 244326 297416 244332
rect 297272 196444 297324 196450
rect 297272 196386 297324 196392
rect 297376 195945 297404 244326
rect 297362 195936 297418 195945
rect 297362 195871 297418 195880
rect 297362 193216 297418 193225
rect 297362 193151 297418 193160
rect 297376 192817 297404 193151
rect 297362 192808 297418 192817
rect 297362 192743 297418 192752
rect 297272 169312 297324 169318
rect 297272 169254 297324 169260
rect 297284 159322 297312 169254
rect 297376 159730 297404 192743
rect 297468 191049 297496 252010
rect 297560 193225 297588 254662
rect 297640 253496 297692 253502
rect 297640 253438 297692 253444
rect 297546 193216 297602 193225
rect 297546 193151 297602 193160
rect 297454 191040 297510 191049
rect 297454 190975 297510 190984
rect 297468 159798 297496 190975
rect 297652 190454 297680 253438
rect 297732 244792 297784 244798
rect 297732 244734 297784 244740
rect 297560 190426 297680 190454
rect 297560 189961 297588 190426
rect 297546 189952 297602 189961
rect 297546 189887 297602 189896
rect 297456 159792 297508 159798
rect 297456 159734 297508 159740
rect 297364 159724 297416 159730
rect 297364 159666 297416 159672
rect 297272 159316 297324 159322
rect 297272 159258 297324 159264
rect 297180 158908 297232 158914
rect 297180 158850 297232 158856
rect 297560 157690 297588 189887
rect 297638 188184 297694 188193
rect 297638 188119 297694 188128
rect 297652 159866 297680 188119
rect 297744 168337 297772 244734
rect 297824 244384 297876 244390
rect 297822 244352 297824 244361
rect 297876 244352 297878 244361
rect 297822 244287 297878 244296
rect 297824 243704 297876 243710
rect 297824 243646 297876 243652
rect 297730 168328 297786 168337
rect 297730 168263 297786 168272
rect 297744 167686 297772 168263
rect 297732 167680 297784 167686
rect 297732 167622 297784 167628
rect 297640 159860 297692 159866
rect 297640 159802 297692 159808
rect 297548 157684 297600 157690
rect 297548 157626 297600 157632
rect 297836 154358 297864 243646
rect 297928 154426 297956 297910
rect 298020 186402 298048 297978
rect 298204 244905 298232 306274
rect 298190 244896 298246 244905
rect 298190 244831 298246 244840
rect 298296 244497 298324 306342
rect 298388 306326 298508 306354
rect 298664 306338 298692 310420
rect 298940 308009 298968 310420
rect 298926 308000 298982 308009
rect 298926 307935 298982 307944
rect 298376 305584 298428 305590
rect 298376 305526 298428 305532
rect 298282 244488 298338 244497
rect 298282 244423 298338 244432
rect 298388 244361 298416 305526
rect 298374 244352 298430 244361
rect 298374 244287 298430 244296
rect 298020 186374 298140 186402
rect 298112 180794 298140 186374
rect 298112 180766 298232 180794
rect 298008 171080 298060 171086
rect 298008 171022 298060 171028
rect 298020 169969 298048 171022
rect 298006 169960 298062 169969
rect 298006 169895 298062 169904
rect 298006 167104 298062 167113
rect 298006 167039 298062 167048
rect 297916 154420 297968 154426
rect 297916 154362 297968 154368
rect 297824 154352 297876 154358
rect 297824 154294 297876 154300
rect 296720 4956 296772 4962
rect 296720 4898 296772 4904
rect 296076 4140 296128 4146
rect 296076 4082 296128 4088
rect 295432 3868 295484 3874
rect 295432 3810 295484 3816
rect 295248 3732 295300 3738
rect 295248 3674 295300 3680
rect 295156 3664 295208 3670
rect 295156 3606 295208 3612
rect 296088 480 296116 4082
rect 298020 3602 298048 167039
rect 298204 153746 298232 180766
rect 298192 153740 298244 153746
rect 298192 153682 298244 153688
rect 298480 16574 298508 306326
rect 298652 306332 298704 306338
rect 298652 306274 298704 306280
rect 299124 305590 299152 310420
rect 299308 306406 299336 310420
rect 299480 306740 299532 306746
rect 299480 306682 299532 306688
rect 299296 306400 299348 306406
rect 299296 306342 299348 306348
rect 299492 306252 299520 306682
rect 299584 306354 299612 310420
rect 299768 306626 299796 310420
rect 299952 306746 299980 310420
rect 299940 306740 299992 306746
rect 299940 306682 299992 306688
rect 299768 306598 299980 306626
rect 299584 306326 299796 306354
rect 299492 306224 299704 306252
rect 299112 305584 299164 305590
rect 299112 305526 299164 305532
rect 299572 305516 299624 305522
rect 299572 305458 299624 305464
rect 299204 305380 299256 305386
rect 299204 305322 299256 305328
rect 298652 248328 298704 248334
rect 298652 248270 298704 248276
rect 298664 243438 298692 248270
rect 299110 245576 299166 245585
rect 299110 245511 299166 245520
rect 298928 244860 298980 244866
rect 298928 244802 298980 244808
rect 298836 244656 298888 244662
rect 298742 244624 298798 244633
rect 298836 244598 298888 244604
rect 298742 244559 298798 244568
rect 298652 243432 298704 243438
rect 298652 243374 298704 243380
rect 298664 196897 298692 243374
rect 298650 196888 298706 196897
rect 298650 196823 298706 196832
rect 298560 196444 298612 196450
rect 298560 196386 298612 196392
rect 298572 159050 298600 196386
rect 298560 159044 298612 159050
rect 298560 158986 298612 158992
rect 298480 16546 298600 16574
rect 298468 5228 298520 5234
rect 298468 5170 298520 5176
rect 298284 4072 298336 4078
rect 298204 4020 298284 4026
rect 298204 4014 298336 4020
rect 298204 3998 298324 4014
rect 298204 3942 298232 3998
rect 298192 3936 298244 3942
rect 298192 3878 298244 3884
rect 297272 3596 297324 3602
rect 297272 3538 297324 3544
rect 298008 3596 298060 3602
rect 298008 3538 298060 3544
rect 297284 480 297312 3538
rect 298480 480 298508 5170
rect 298572 4894 298600 16546
rect 298560 4888 298612 4894
rect 298560 4830 298612 4836
rect 298756 3942 298784 244559
rect 298848 193769 298876 244598
rect 298834 193760 298890 193769
rect 298834 193695 298890 193704
rect 298848 159934 298876 193695
rect 298940 188193 298968 244802
rect 299124 244322 299152 245511
rect 299112 244316 299164 244322
rect 299112 244258 299164 244264
rect 299020 243908 299072 243914
rect 299020 243850 299072 243856
rect 298926 188184 298982 188193
rect 298926 188119 298982 188128
rect 298836 159928 298888 159934
rect 298836 159870 298888 159876
rect 298928 159656 298980 159662
rect 298928 159598 298980 159604
rect 298940 155922 298968 159598
rect 299032 158574 299060 243850
rect 299112 243840 299164 243846
rect 299112 243782 299164 243788
rect 299124 158681 299152 243782
rect 299110 158672 299166 158681
rect 299110 158607 299166 158616
rect 299020 158568 299072 158574
rect 299020 158510 299072 158516
rect 299124 157554 299152 158607
rect 299216 157622 299244 305322
rect 299480 305176 299532 305182
rect 299480 305118 299532 305124
rect 299296 305108 299348 305114
rect 299296 305050 299348 305056
rect 299308 159662 299336 305050
rect 299388 254788 299440 254794
rect 299388 254730 299440 254736
rect 299400 168065 299428 254730
rect 299492 244769 299520 305118
rect 299584 245206 299612 305458
rect 299572 245200 299624 245206
rect 299572 245142 299624 245148
rect 299676 245041 299704 306224
rect 299662 245032 299718 245041
rect 299768 245002 299796 306326
rect 299848 306332 299900 306338
rect 299848 306274 299900 306280
rect 299860 247489 299888 306274
rect 299952 248169 299980 306598
rect 300124 305584 300176 305590
rect 300124 305526 300176 305532
rect 300136 305318 300164 305526
rect 300124 305312 300176 305318
rect 300124 305254 300176 305260
rect 300228 305182 300256 310420
rect 300412 306338 300440 310420
rect 300400 306332 300452 306338
rect 300400 306274 300452 306280
rect 300596 305522 300624 310420
rect 300584 305516 300636 305522
rect 300584 305458 300636 305464
rect 300216 305176 300268 305182
rect 300216 305118 300268 305124
rect 299938 248160 299994 248169
rect 299938 248095 299994 248104
rect 299846 247480 299902 247489
rect 299846 247415 299902 247424
rect 300768 246696 300820 246702
rect 300768 246638 300820 246644
rect 299662 244967 299718 244976
rect 299756 244996 299808 245002
rect 299756 244938 299808 244944
rect 299478 244760 299534 244769
rect 299478 244695 299534 244704
rect 300780 243982 300808 246638
rect 300872 244934 300900 310420
rect 301070 310406 301176 310434
rect 301044 306400 301096 306406
rect 301044 306342 301096 306348
rect 300952 306332 301004 306338
rect 300952 306274 301004 306280
rect 300860 244928 300912 244934
rect 300860 244870 300912 244876
rect 300964 244361 300992 306274
rect 301056 245177 301084 306342
rect 301148 248305 301176 310406
rect 301332 308281 301360 310420
rect 301318 308272 301374 308281
rect 301318 308207 301374 308216
rect 301516 306338 301544 310420
rect 301504 306332 301556 306338
rect 301504 306274 301556 306280
rect 301596 306332 301648 306338
rect 301596 306274 301648 306280
rect 301608 305250 301636 306274
rect 301596 305244 301648 305250
rect 301596 305186 301648 305192
rect 301700 296714 301728 310420
rect 301976 308961 302004 310420
rect 301962 308952 302018 308961
rect 301962 308887 302018 308896
rect 302160 306406 302188 310420
rect 302358 310406 302464 310434
rect 302240 306468 302292 306474
rect 302240 306410 302292 306416
rect 302148 306400 302200 306406
rect 302148 306342 302200 306348
rect 301240 296686 301728 296714
rect 301134 248296 301190 248305
rect 301134 248231 301190 248240
rect 301240 248033 301268 296686
rect 301226 248024 301282 248033
rect 301226 247959 301282 247968
rect 302252 245313 302280 306410
rect 302436 306082 302464 310406
rect 302528 310406 302634 310434
rect 302528 306474 302556 310406
rect 302516 306468 302568 306474
rect 302516 306410 302568 306416
rect 302436 306054 302556 306082
rect 302332 305380 302384 305386
rect 302332 305322 302384 305328
rect 302344 245614 302372 305322
rect 302424 305244 302476 305250
rect 302424 305186 302476 305192
rect 302332 245608 302384 245614
rect 302332 245550 302384 245556
rect 302238 245304 302294 245313
rect 302436 245274 302464 305186
rect 302528 247897 302556 306054
rect 302804 305386 302832 310420
rect 302792 305380 302844 305386
rect 302792 305322 302844 305328
rect 302608 305312 302660 305318
rect 302608 305254 302660 305260
rect 302514 247888 302570 247897
rect 302514 247823 302570 247832
rect 302620 247761 302648 305254
rect 302988 296714 303016 310420
rect 303080 310406 303278 310434
rect 303080 305250 303108 310406
rect 303448 305318 303476 310420
rect 303436 305312 303488 305318
rect 303436 305254 303488 305260
rect 303068 305244 303120 305250
rect 303068 305186 303120 305192
rect 303632 304366 303660 310420
rect 303724 310406 303922 310434
rect 303620 304360 303672 304366
rect 303620 304302 303672 304308
rect 303620 304224 303672 304230
rect 303620 304166 303672 304172
rect 302712 296686 303016 296714
rect 302606 247752 302662 247761
rect 302606 247687 302662 247696
rect 302712 247625 302740 296686
rect 302698 247616 302754 247625
rect 302698 247551 302754 247560
rect 302238 245239 302294 245248
rect 302424 245268 302476 245274
rect 302424 245210 302476 245216
rect 301042 245168 301098 245177
rect 301042 245103 301098 245112
rect 303632 244390 303660 304166
rect 303724 245070 303752 310406
rect 304092 306354 304120 310420
rect 303816 306326 304120 306354
rect 304184 310406 304382 310434
rect 303816 248402 303844 306326
rect 304184 306218 304212 310406
rect 303908 306190 304212 306218
rect 303804 248396 303856 248402
rect 303804 248338 303856 248344
rect 303908 247586 303936 306190
rect 304552 304570 304580 310420
rect 304540 304564 304592 304570
rect 304540 304506 304592 304512
rect 304736 304450 304764 310420
rect 305012 308961 305040 310420
rect 304998 308952 305054 308961
rect 304998 308887 305054 308896
rect 305196 306354 305224 310420
rect 304000 304422 304764 304450
rect 305012 306326 305224 306354
rect 304000 247790 304028 304422
rect 304080 304360 304132 304366
rect 304080 304302 304132 304308
rect 304092 247926 304120 304302
rect 304080 247920 304132 247926
rect 304080 247862 304132 247868
rect 303988 247784 304040 247790
rect 303988 247726 304040 247732
rect 303896 247580 303948 247586
rect 303896 247522 303948 247528
rect 305012 245410 305040 306326
rect 305092 305108 305144 305114
rect 305092 305050 305144 305056
rect 305000 245404 305052 245410
rect 305000 245346 305052 245352
rect 305104 245342 305132 305050
rect 305380 304314 305408 310420
rect 305184 304292 305236 304298
rect 305184 304234 305236 304240
rect 305288 304286 305408 304314
rect 305472 310406 305670 310434
rect 305472 304298 305500 310406
rect 305840 305114 305868 310420
rect 305828 305108 305880 305114
rect 305828 305050 305880 305056
rect 305460 304292 305512 304298
rect 305196 247654 305224 304234
rect 305288 247722 305316 304286
rect 305460 304234 305512 304240
rect 306024 302234 306052 310420
rect 305380 302206 306052 302234
rect 306116 310406 306314 310434
rect 305380 247858 305408 302206
rect 306116 296714 306144 310406
rect 306484 306490 306512 310420
rect 306392 306462 306512 306490
rect 306576 310406 306774 310434
rect 306392 305386 306420 306462
rect 306576 306354 306604 310406
rect 306484 306326 306604 306354
rect 306656 306400 306708 306406
rect 306944 306354 306972 310420
rect 307128 306406 307156 310420
rect 307220 310406 307418 310434
rect 306656 306342 306708 306348
rect 306380 305380 306432 305386
rect 306380 305322 306432 305328
rect 306380 305244 306432 305250
rect 306380 305186 306432 305192
rect 305472 296686 306144 296714
rect 305368 247852 305420 247858
rect 305368 247794 305420 247800
rect 305276 247716 305328 247722
rect 305276 247658 305328 247664
rect 305184 247648 305236 247654
rect 305184 247590 305236 247596
rect 305472 247518 305500 296686
rect 305460 247512 305512 247518
rect 305460 247454 305512 247460
rect 305092 245336 305144 245342
rect 305092 245278 305144 245284
rect 303712 245064 303764 245070
rect 303712 245006 303764 245012
rect 306392 245002 306420 305186
rect 306484 245206 306512 306326
rect 306564 305312 306616 305318
rect 306564 305254 306616 305260
rect 306472 245200 306524 245206
rect 306472 245142 306524 245148
rect 306576 245070 306604 305254
rect 306668 245478 306696 306342
rect 306760 306326 306972 306354
rect 307116 306400 307168 306406
rect 307116 306342 307168 306348
rect 306656 245472 306708 245478
rect 306656 245414 306708 245420
rect 306760 245274 306788 306326
rect 306840 305380 306892 305386
rect 306840 305322 306892 305328
rect 306748 245268 306800 245274
rect 306748 245210 306800 245216
rect 306564 245064 306616 245070
rect 306564 245006 306616 245012
rect 306380 244996 306432 245002
rect 306380 244938 306432 244944
rect 306852 244730 306880 305322
rect 307220 305250 307248 310406
rect 307588 305318 307616 310420
rect 307786 310406 307892 310434
rect 307760 306536 307812 306542
rect 307760 306478 307812 306484
rect 307576 305312 307628 305318
rect 307576 305254 307628 305260
rect 307208 305244 307260 305250
rect 307208 305186 307260 305192
rect 307772 245138 307800 306478
rect 307864 245410 307892 310406
rect 308048 307970 308076 310420
rect 308036 307964 308088 307970
rect 308036 307906 308088 307912
rect 308036 306468 308088 306474
rect 308036 306410 308088 306416
rect 307944 305380 307996 305386
rect 307944 305322 307996 305328
rect 307956 245546 307984 305322
rect 307944 245540 307996 245546
rect 307944 245482 307996 245488
rect 307852 245404 307904 245410
rect 307852 245346 307904 245352
rect 308048 245342 308076 306410
rect 308128 306400 308180 306406
rect 308128 306342 308180 306348
rect 308140 247858 308168 306342
rect 308232 247926 308260 310420
rect 308416 306542 308444 310420
rect 308508 310406 308706 310434
rect 308404 306536 308456 306542
rect 308404 306478 308456 306484
rect 308508 306474 308536 310406
rect 308496 306468 308548 306474
rect 308496 306410 308548 306416
rect 308876 306406 308904 310420
rect 308864 306400 308916 306406
rect 308864 306342 308916 306348
rect 309060 305386 309088 310420
rect 309152 310406 309350 310434
rect 309048 305380 309100 305386
rect 309048 305322 309100 305328
rect 308220 247920 308272 247926
rect 308220 247862 308272 247868
rect 308128 247852 308180 247858
rect 308128 247794 308180 247800
rect 308036 245336 308088 245342
rect 308036 245278 308088 245284
rect 309152 245177 309180 310406
rect 309520 309134 309548 310420
rect 309428 309106 309548 309134
rect 309612 310406 309810 310434
rect 309324 306400 309376 306406
rect 309324 306342 309376 306348
rect 309232 304292 309284 304298
rect 309232 304234 309284 304240
rect 309244 245478 309272 304234
rect 309232 245472 309284 245478
rect 309232 245414 309284 245420
rect 309138 245168 309194 245177
rect 307760 245132 307812 245138
rect 309138 245103 309194 245112
rect 307760 245074 307812 245080
rect 309336 245041 309364 306342
rect 309428 247625 309456 309106
rect 309612 304298 309640 310406
rect 309980 306406 310008 310420
rect 309968 306400 310020 306406
rect 309968 306342 310020 306348
rect 309600 304292 309652 304298
rect 309600 304234 309652 304240
rect 310164 302234 310192 310420
rect 309520 302206 310192 302234
rect 310256 310406 310454 310434
rect 309520 253366 309548 302206
rect 310256 296714 310284 310406
rect 310520 306468 310572 306474
rect 310520 306410 310572 306416
rect 309612 296686 310284 296714
rect 309612 275233 309640 296686
rect 309598 275224 309654 275233
rect 309598 275159 309654 275168
rect 309508 253360 309560 253366
rect 309508 253302 309560 253308
rect 310532 250578 310560 306410
rect 310624 305386 310652 310420
rect 310822 310406 310928 310434
rect 310704 306400 310756 306406
rect 310704 306342 310756 306348
rect 310612 305380 310664 305386
rect 310612 305322 310664 305328
rect 310612 305244 310664 305250
rect 310612 305186 310664 305192
rect 310624 274106 310652 305186
rect 310716 283762 310744 306342
rect 310900 305538 310928 310406
rect 310900 305510 311020 305538
rect 310888 305380 310940 305386
rect 310888 305322 310940 305328
rect 310796 304292 310848 304298
rect 310796 304234 310848 304240
rect 310808 285122 310836 304234
rect 310900 287745 310928 305322
rect 310992 289270 311020 305510
rect 311084 304298 311112 310420
rect 311268 306474 311296 310420
rect 311256 306468 311308 306474
rect 311256 306410 311308 306416
rect 311452 306406 311480 310420
rect 311544 310406 311742 310434
rect 311926 310406 312032 310434
rect 311440 306400 311492 306406
rect 311440 306342 311492 306348
rect 311544 305250 311572 310406
rect 311900 308100 311952 308106
rect 311900 308042 311952 308048
rect 311532 305244 311584 305250
rect 311532 305186 311584 305192
rect 311072 304292 311124 304298
rect 311072 304234 311124 304240
rect 310980 289264 311032 289270
rect 310980 289206 311032 289212
rect 310886 287736 310942 287745
rect 310886 287671 310942 287680
rect 310796 285116 310848 285122
rect 310796 285058 310848 285064
rect 310704 283756 310756 283762
rect 310704 283698 310756 283704
rect 310612 274100 310664 274106
rect 310612 274042 310664 274048
rect 310520 250572 310572 250578
rect 310520 250514 310572 250520
rect 309414 247616 309470 247625
rect 309414 247551 309470 247560
rect 311912 246498 311940 308042
rect 312004 260302 312032 310406
rect 312084 308440 312136 308446
rect 312084 308382 312136 308388
rect 312096 271318 312124 308382
rect 312188 308174 312216 310420
rect 312372 308394 312400 310420
rect 312280 308366 312400 308394
rect 312176 308168 312228 308174
rect 312176 308110 312228 308116
rect 312176 308032 312228 308038
rect 312176 307974 312228 307980
rect 312188 280974 312216 307974
rect 312280 286550 312308 308366
rect 312360 308168 312412 308174
rect 312360 308110 312412 308116
rect 312372 303249 312400 308110
rect 312556 308106 312584 310420
rect 312832 308281 312860 310420
rect 313016 308446 313044 310420
rect 313004 308440 313056 308446
rect 313004 308382 313056 308388
rect 312818 308272 312874 308281
rect 312818 308207 312874 308216
rect 312544 308100 312596 308106
rect 312544 308042 312596 308048
rect 313200 308038 313228 310420
rect 313372 308440 313424 308446
rect 313372 308382 313424 308388
rect 313280 308100 313332 308106
rect 313280 308042 313332 308048
rect 313188 308032 313240 308038
rect 313188 307974 313240 307980
rect 312358 303240 312414 303249
rect 312358 303175 312414 303184
rect 312268 286544 312320 286550
rect 312268 286486 312320 286492
rect 312176 280968 312228 280974
rect 312176 280910 312228 280916
rect 312084 271312 312136 271318
rect 312084 271254 312136 271260
rect 311992 260296 312044 260302
rect 311992 260238 312044 260244
rect 313292 249150 313320 308042
rect 313384 269958 313412 308382
rect 313476 282334 313504 310420
rect 313660 308446 313688 310420
rect 313648 308440 313700 308446
rect 313648 308382 313700 308388
rect 313556 308168 313608 308174
rect 313556 308110 313608 308116
rect 313568 283694 313596 308110
rect 313844 296714 313872 310420
rect 313922 308272 313978 308281
rect 313922 308207 313978 308216
rect 313660 296686 313872 296714
rect 313660 286414 313688 296686
rect 313936 287774 313964 308207
rect 314120 308009 314148 310420
rect 314304 308174 314332 310420
rect 314292 308168 314344 308174
rect 314292 308110 314344 308116
rect 314488 308106 314516 310420
rect 314660 308440 314712 308446
rect 314660 308382 314712 308388
rect 314476 308100 314528 308106
rect 314476 308042 314528 308048
rect 314106 308000 314162 308009
rect 314106 307935 314162 307944
rect 313924 287768 313976 287774
rect 313924 287710 313976 287716
rect 313648 286408 313700 286414
rect 313648 286350 313700 286356
rect 313556 283688 313608 283694
rect 313556 283630 313608 283636
rect 313464 282328 313516 282334
rect 313464 282270 313516 282276
rect 313372 269952 313424 269958
rect 313372 269894 313424 269900
rect 314672 258874 314700 308382
rect 314764 308174 314792 310420
rect 314948 308394 314976 310420
rect 314856 308366 314976 308394
rect 315040 310406 315238 310434
rect 314752 308168 314804 308174
rect 314752 308110 314804 308116
rect 314752 308032 314804 308038
rect 314752 307974 314804 307980
rect 314764 267238 314792 307974
rect 314856 268530 314884 308366
rect 314936 308168 314988 308174
rect 314936 308110 314988 308116
rect 314948 279614 314976 308110
rect 314936 279608 314988 279614
rect 314936 279550 314988 279556
rect 315040 279546 315068 310406
rect 315408 304502 315436 310420
rect 315592 308038 315620 310420
rect 315684 310406 315882 310434
rect 315684 308446 315712 310406
rect 315672 308440 315724 308446
rect 315672 308382 315724 308388
rect 315764 308440 315816 308446
rect 315764 308382 315816 308388
rect 315580 308032 315632 308038
rect 315580 307974 315632 307980
rect 315776 307970 315804 308382
rect 315764 307964 315816 307970
rect 315764 307906 315816 307912
rect 315396 304496 315448 304502
rect 315396 304438 315448 304444
rect 315028 279540 315080 279546
rect 315028 279482 315080 279488
rect 314844 268524 314896 268530
rect 314844 268466 314896 268472
rect 314752 267232 314804 267238
rect 314752 267174 314804 267180
rect 314660 258868 314712 258874
rect 314660 258810 314712 258816
rect 316052 254658 316080 310420
rect 316250 310406 316356 310434
rect 316328 308258 316356 310406
rect 316512 308394 316540 310420
rect 316512 308366 316632 308394
rect 316328 308230 316540 308258
rect 316316 308168 316368 308174
rect 316316 308110 316368 308116
rect 316224 308100 316276 308106
rect 316224 308042 316276 308048
rect 316132 308032 316184 308038
rect 316132 307974 316184 307980
rect 316040 254652 316092 254658
rect 316040 254594 316092 254600
rect 316144 254590 316172 307974
rect 316236 297566 316264 308042
rect 316328 300393 316356 308110
rect 316512 307222 316540 308230
rect 316500 307216 316552 307222
rect 316500 307158 316552 307164
rect 316604 301646 316632 308366
rect 316696 308281 316724 310420
rect 316682 308272 316738 308281
rect 316682 308207 316738 308216
rect 316880 308174 316908 310420
rect 316972 310406 317170 310434
rect 316868 308168 316920 308174
rect 316868 308110 316920 308116
rect 316972 308106 317000 310406
rect 316960 308100 317012 308106
rect 316960 308042 317012 308048
rect 317340 308038 317368 310420
rect 317616 308394 317644 310420
rect 317616 308366 317736 308394
rect 317604 308168 317656 308174
rect 317604 308110 317656 308116
rect 317512 308100 317564 308106
rect 317512 308042 317564 308048
rect 317328 308032 317380 308038
rect 317328 307974 317380 307980
rect 317420 308032 317472 308038
rect 317420 307974 317472 307980
rect 316592 301640 316644 301646
rect 316592 301582 316644 301588
rect 316314 300384 316370 300393
rect 316314 300319 316370 300328
rect 316224 297560 316276 297566
rect 316224 297502 316276 297508
rect 317432 264314 317460 307974
rect 317524 265810 317552 308042
rect 317616 276758 317644 308110
rect 317708 282266 317736 308366
rect 317800 308174 317828 310420
rect 317788 308168 317840 308174
rect 317788 308110 317840 308116
rect 317984 297634 318012 310420
rect 318062 308000 318118 308009
rect 318062 307935 318118 307944
rect 317972 297628 318024 297634
rect 317972 297570 318024 297576
rect 318076 286482 318104 307935
rect 318260 307154 318288 310420
rect 318444 308106 318472 310420
rect 318432 308100 318484 308106
rect 318432 308042 318484 308048
rect 318628 308038 318656 310420
rect 318812 310406 318918 310434
rect 318812 308038 318840 310406
rect 319088 308394 319116 310420
rect 318904 308366 319116 308394
rect 318616 308032 318668 308038
rect 318616 307974 318668 307980
rect 318800 308032 318852 308038
rect 318800 307974 318852 307980
rect 318800 307896 318852 307902
rect 318800 307838 318852 307844
rect 318248 307148 318300 307154
rect 318248 307090 318300 307096
rect 318064 286476 318116 286482
rect 318064 286418 318116 286424
rect 317696 282260 317748 282266
rect 317696 282202 317748 282208
rect 317604 276752 317656 276758
rect 317604 276694 317656 276700
rect 317512 265804 317564 265810
rect 317512 265746 317564 265752
rect 317420 264308 317472 264314
rect 317420 264250 317472 264256
rect 318812 262954 318840 307838
rect 318904 264246 318932 308366
rect 319272 308258 319300 310420
rect 318996 308230 319300 308258
rect 319364 310406 319562 310434
rect 318996 278118 319024 308230
rect 319076 308168 319128 308174
rect 319364 308156 319392 310406
rect 319442 308272 319498 308281
rect 319442 308207 319498 308216
rect 319076 308110 319128 308116
rect 319180 308128 319392 308156
rect 319088 280906 319116 308110
rect 319180 303113 319208 308128
rect 319260 308032 319312 308038
rect 319260 307974 319312 307980
rect 319272 304434 319300 307974
rect 319260 304428 319312 304434
rect 319260 304370 319312 304376
rect 319166 303104 319222 303113
rect 319166 303039 319222 303048
rect 319076 280900 319128 280906
rect 319076 280842 319128 280848
rect 318984 278112 319036 278118
rect 318984 278054 319036 278060
rect 318892 264240 318944 264246
rect 318892 264182 318944 264188
rect 318800 262948 318852 262954
rect 318800 262890 318852 262896
rect 319456 258806 319484 308207
rect 319732 308174 319760 310420
rect 319720 308168 319772 308174
rect 319720 308110 319772 308116
rect 319916 307902 319944 310420
rect 319904 307896 319956 307902
rect 319904 307838 319956 307844
rect 320192 306746 320220 310420
rect 320390 310406 320496 310434
rect 320272 308168 320324 308174
rect 320272 308110 320324 308116
rect 320180 306740 320232 306746
rect 320180 306682 320232 306688
rect 320180 306604 320232 306610
rect 320180 306546 320232 306552
rect 320192 261594 320220 306546
rect 320284 262886 320312 308110
rect 320364 307692 320416 307698
rect 320364 307634 320416 307640
rect 320376 275398 320404 307634
rect 320468 279478 320496 310406
rect 320560 310406 320666 310434
rect 320560 307698 320588 310406
rect 320836 308394 320864 310420
rect 320652 308366 320864 308394
rect 320548 307692 320600 307698
rect 320548 307634 320600 307640
rect 320548 307556 320600 307562
rect 320548 307498 320600 307504
rect 320560 300257 320588 307498
rect 320652 301578 320680 308366
rect 321020 308174 321048 310420
rect 321112 310406 321310 310434
rect 321008 308168 321060 308174
rect 321008 308110 321060 308116
rect 320732 306740 320784 306746
rect 320732 306682 320784 306688
rect 320744 306105 320772 306682
rect 321112 306610 321140 310406
rect 321480 307562 321508 310420
rect 321678 310406 321876 310434
rect 321468 307556 321520 307562
rect 321468 307498 321520 307504
rect 321100 306604 321152 306610
rect 321100 306546 321152 306552
rect 320730 306096 320786 306105
rect 320730 306031 320786 306040
rect 321652 305380 321704 305386
rect 321652 305322 321704 305328
rect 321560 305244 321612 305250
rect 321560 305186 321612 305192
rect 320640 301572 320692 301578
rect 320640 301514 320692 301520
rect 320546 300248 320602 300257
rect 320546 300183 320602 300192
rect 320456 279472 320508 279478
rect 320456 279414 320508 279420
rect 320364 275392 320416 275398
rect 320364 275334 320416 275340
rect 320272 262880 320324 262886
rect 320272 262822 320324 262828
rect 320180 261588 320232 261594
rect 320180 261530 320232 261536
rect 319444 258800 319496 258806
rect 319444 258742 319496 258748
rect 316132 254584 316184 254590
rect 316132 254526 316184 254532
rect 321572 252006 321600 305186
rect 321664 261526 321692 305322
rect 321848 294778 321876 310406
rect 321836 294772 321888 294778
rect 321836 294714 321888 294720
rect 321940 292574 321968 310420
rect 322124 307086 322152 310420
rect 322112 307080 322164 307086
rect 322112 307022 322164 307028
rect 322308 305386 322336 310420
rect 322400 310406 322598 310434
rect 322296 305380 322348 305386
rect 322296 305322 322348 305328
rect 322400 305250 322428 310406
rect 322388 305244 322440 305250
rect 322388 305186 322440 305192
rect 322768 298926 322796 310420
rect 322940 306672 322992 306678
rect 322940 306614 322992 306620
rect 322756 298920 322808 298926
rect 322756 298862 322808 298868
rect 321756 292546 321968 292574
rect 321756 274038 321784 292546
rect 321744 274032 321796 274038
rect 321744 273974 321796 273980
rect 321652 261520 321704 261526
rect 321652 261462 321704 261468
rect 321560 252000 321612 252006
rect 321560 251942 321612 251948
rect 313280 249144 313332 249150
rect 313280 249086 313332 249092
rect 322952 247790 322980 306614
rect 323044 306592 323072 310420
rect 323228 306610 323256 310420
rect 323216 306604 323268 306610
rect 323044 306564 323164 306592
rect 323136 306490 323164 306564
rect 323216 306546 323268 306552
rect 323136 306462 323256 306490
rect 323124 306400 323176 306406
rect 323124 306342 323176 306348
rect 323136 306218 323164 306342
rect 323044 306190 323164 306218
rect 323044 251938 323072 306190
rect 323124 305380 323176 305386
rect 323124 305322 323176 305328
rect 323136 271250 323164 305322
rect 323228 278050 323256 306462
rect 323308 306400 323360 306406
rect 323308 306342 323360 306348
rect 323320 296138 323348 306342
rect 323412 297498 323440 310420
rect 323504 310406 323702 310434
rect 323504 306678 323532 310406
rect 323492 306672 323544 306678
rect 323492 306614 323544 306620
rect 323872 305386 323900 310420
rect 324056 306406 324084 310420
rect 324332 306406 324360 310420
rect 324516 309134 324544 310420
rect 324424 309106 324544 309134
rect 324044 306400 324096 306406
rect 324044 306342 324096 306348
rect 324320 306400 324372 306406
rect 324320 306342 324372 306348
rect 323860 305380 323912 305386
rect 323860 305322 323912 305328
rect 324320 305312 324372 305318
rect 324320 305254 324372 305260
rect 323400 297492 323452 297498
rect 323400 297434 323452 297440
rect 323308 296132 323360 296138
rect 323308 296074 323360 296080
rect 323216 278044 323268 278050
rect 323216 277986 323268 277992
rect 323124 271244 323176 271250
rect 323124 271186 323176 271192
rect 323032 251932 323084 251938
rect 323032 251874 323084 251880
rect 322940 247784 322992 247790
rect 322940 247726 322992 247732
rect 311900 246492 311952 246498
rect 311900 246434 311952 246440
rect 309322 245032 309378 245041
rect 309322 244967 309378 244976
rect 324332 244934 324360 305254
rect 324424 250510 324452 309106
rect 324596 306400 324648 306406
rect 324596 306342 324648 306348
rect 324504 305380 324556 305386
rect 324504 305322 324556 305328
rect 324516 272542 324544 305322
rect 324608 276690 324636 306342
rect 324700 304366 324728 310420
rect 324792 310406 324990 310434
rect 324688 304360 324740 304366
rect 324688 304302 324740 304308
rect 324792 292574 324820 310406
rect 325160 305386 325188 310420
rect 325344 305969 325372 310420
rect 325436 310406 325634 310434
rect 325818 310406 326016 310434
rect 325330 305960 325386 305969
rect 325330 305895 325386 305904
rect 325148 305380 325200 305386
rect 325148 305322 325200 305328
rect 325436 305318 325464 310406
rect 325792 306536 325844 306542
rect 325792 306478 325844 306484
rect 325700 306468 325752 306474
rect 325700 306410 325752 306416
rect 325424 305312 325476 305318
rect 325424 305254 325476 305260
rect 324700 292546 324820 292574
rect 324700 285054 324728 292546
rect 324688 285048 324740 285054
rect 324688 284990 324740 284996
rect 324596 276684 324648 276690
rect 324596 276626 324648 276632
rect 324504 272536 324556 272542
rect 324504 272478 324556 272484
rect 325712 269890 325740 306410
rect 325804 275330 325832 306478
rect 325884 306400 325936 306406
rect 325884 306342 325936 306348
rect 325896 293418 325924 306342
rect 325988 294710 326016 310406
rect 326080 302977 326108 310420
rect 326264 306406 326292 310420
rect 326448 306474 326476 310420
rect 326724 307290 326752 310420
rect 326712 307284 326764 307290
rect 326712 307226 326764 307232
rect 326908 306542 326936 310420
rect 327106 310406 327212 310434
rect 326896 306536 326948 306542
rect 326896 306478 326948 306484
rect 326436 306468 326488 306474
rect 326436 306410 326488 306416
rect 327080 306468 327132 306474
rect 327080 306410 327132 306416
rect 326252 306400 326304 306406
rect 326252 306342 326304 306348
rect 326066 302968 326122 302977
rect 326066 302903 326122 302912
rect 325976 294704 326028 294710
rect 325976 294646 326028 294652
rect 325884 293412 325936 293418
rect 325884 293354 325936 293360
rect 325792 275324 325844 275330
rect 325792 275266 325844 275272
rect 325700 269884 325752 269890
rect 325700 269826 325752 269832
rect 324412 250504 324464 250510
rect 324412 250446 324464 250452
rect 327092 246430 327120 306410
rect 327184 247722 327212 310406
rect 327368 306542 327396 310420
rect 327356 306536 327408 306542
rect 327356 306478 327408 306484
rect 327552 306456 327580 310420
rect 327460 306428 327580 306456
rect 327264 306400 327316 306406
rect 327460 306354 327488 306428
rect 327736 306406 327764 310420
rect 327828 310406 328026 310434
rect 327264 306342 327316 306348
rect 327276 268462 327304 306342
rect 327368 306326 327488 306354
rect 327724 306400 327776 306406
rect 327724 306342 327776 306348
rect 327368 273970 327396 306326
rect 327828 306082 327856 310406
rect 327908 306536 327960 306542
rect 327908 306478 327960 306484
rect 327460 306054 327856 306082
rect 327460 293350 327488 306054
rect 327920 305946 327948 306478
rect 328196 306474 328224 310420
rect 328368 306536 328420 306542
rect 328368 306478 328420 306484
rect 328184 306468 328236 306474
rect 328184 306410 328236 306416
rect 328380 306218 328408 306478
rect 328472 306354 328500 310420
rect 328656 307766 328684 310420
rect 328644 307760 328696 307766
rect 328644 307702 328696 307708
rect 328472 306326 328776 306354
rect 328380 306190 328500 306218
rect 327552 305918 327948 305946
rect 327552 294642 327580 305918
rect 327540 294636 327592 294642
rect 327540 294578 327592 294584
rect 327448 293344 327500 293350
rect 327448 293286 327500 293292
rect 327356 273964 327408 273970
rect 327356 273906 327408 273912
rect 327264 268456 327316 268462
rect 327264 268398 327316 268404
rect 327172 247716 327224 247722
rect 327172 247658 327224 247664
rect 327080 246424 327132 246430
rect 327080 246366 327132 246372
rect 324320 244928 324372 244934
rect 328472 244905 328500 306190
rect 328644 305380 328696 305386
rect 328644 305322 328696 305328
rect 328552 305312 328604 305318
rect 328552 305254 328604 305260
rect 328564 267170 328592 305254
rect 328656 271182 328684 305322
rect 328748 284986 328776 306326
rect 328840 291922 328868 310420
rect 328932 310406 329130 310434
rect 328932 306542 328960 310406
rect 328920 306536 328972 306542
rect 328920 306478 328972 306484
rect 329300 299474 329328 310420
rect 329380 307760 329432 307766
rect 329380 307702 329432 307708
rect 329392 301510 329420 307702
rect 329484 305386 329512 310420
rect 329576 310406 329774 310434
rect 329472 305380 329524 305386
rect 329472 305322 329524 305328
rect 329576 305318 329604 310406
rect 329840 306740 329892 306746
rect 329840 306682 329892 306688
rect 329564 305312 329616 305318
rect 329564 305254 329616 305260
rect 329380 301504 329432 301510
rect 329380 301446 329432 301452
rect 328932 299446 329328 299474
rect 328828 291916 328880 291922
rect 328828 291858 328880 291864
rect 328932 291854 328960 299446
rect 328920 291848 328972 291854
rect 328920 291790 328972 291796
rect 328736 284980 328788 284986
rect 328736 284922 328788 284928
rect 328644 271176 328696 271182
rect 328644 271118 328696 271124
rect 328552 267164 328604 267170
rect 328552 267106 328604 267112
rect 329852 265742 329880 306682
rect 329944 306592 329972 310420
rect 329944 306564 330064 306592
rect 330036 306354 330064 306564
rect 330128 306456 330156 310420
rect 330220 310406 330418 310434
rect 330220 306746 330248 310406
rect 330208 306740 330260 306746
rect 330208 306682 330260 306688
rect 330128 306428 330340 306456
rect 330036 306326 330248 306354
rect 330024 305380 330076 305386
rect 330024 305322 330076 305328
rect 329932 305244 329984 305250
rect 329932 305186 329984 305192
rect 329944 269822 329972 305186
rect 330036 290562 330064 305322
rect 330116 305312 330168 305318
rect 330116 305254 330168 305260
rect 330128 296070 330156 305254
rect 330220 300121 330248 306326
rect 330312 302841 330340 306428
rect 330588 305386 330616 310420
rect 330576 305380 330628 305386
rect 330576 305322 330628 305328
rect 330772 305250 330800 310420
rect 330864 310406 331062 310434
rect 330864 305318 330892 310406
rect 331128 306264 331180 306270
rect 331128 306206 331180 306212
rect 331140 305833 331168 306206
rect 331126 305824 331182 305833
rect 331126 305759 331182 305768
rect 331232 305386 331260 310420
rect 331312 306468 331364 306474
rect 331312 306410 331364 306416
rect 331220 305380 331272 305386
rect 331220 305322 331272 305328
rect 330852 305312 330904 305318
rect 330852 305254 330904 305260
rect 330760 305244 330812 305250
rect 330760 305186 330812 305192
rect 331220 305040 331272 305046
rect 331220 304982 331272 304988
rect 330298 302832 330354 302841
rect 330298 302767 330354 302776
rect 330206 300112 330262 300121
rect 330206 300047 330262 300056
rect 330116 296064 330168 296070
rect 330116 296006 330168 296012
rect 330024 290556 330076 290562
rect 330024 290498 330076 290504
rect 329932 269816 329984 269822
rect 329932 269758 329984 269764
rect 329840 265736 329892 265742
rect 329840 265678 329892 265684
rect 331232 246362 331260 304982
rect 331324 249082 331352 306410
rect 331404 306264 331456 306270
rect 331404 306206 331456 306212
rect 331416 267102 331444 306206
rect 331508 268394 331536 310420
rect 331692 306474 331720 310420
rect 331680 306468 331732 306474
rect 331680 306410 331732 306416
rect 331588 306400 331640 306406
rect 331876 306354 331904 310420
rect 331588 306342 331640 306348
rect 331600 287706 331628 306342
rect 331692 306326 331904 306354
rect 331968 310406 332166 310434
rect 331692 289202 331720 306326
rect 331968 306270 331996 310406
rect 331956 306264 332008 306270
rect 331956 306206 332008 306212
rect 332230 305824 332286 305833
rect 332230 305759 332286 305768
rect 331864 305516 331916 305522
rect 331864 305458 331916 305464
rect 331772 305380 331824 305386
rect 331772 305322 331824 305328
rect 331784 298858 331812 305322
rect 331876 305114 331904 305458
rect 332244 305386 332272 305759
rect 332232 305380 332284 305386
rect 332232 305322 332284 305328
rect 331864 305108 331916 305114
rect 331864 305050 331916 305056
rect 332336 305046 332364 310420
rect 332520 306406 332548 310420
rect 332508 306400 332560 306406
rect 332508 306342 332560 306348
rect 332600 306264 332652 306270
rect 332600 306206 332652 306212
rect 332324 305040 332376 305046
rect 332324 304982 332376 304988
rect 331772 298852 331824 298858
rect 331772 298794 331824 298800
rect 331680 289196 331732 289202
rect 331680 289138 331732 289144
rect 331588 287700 331640 287706
rect 331588 287642 331640 287648
rect 331496 268388 331548 268394
rect 331496 268330 331548 268336
rect 331404 267096 331456 267102
rect 331404 267038 331456 267044
rect 332612 251870 332640 306206
rect 332796 305674 332824 310420
rect 332980 306270 333008 310420
rect 332968 306264 333020 306270
rect 332968 306206 333020 306212
rect 332796 305646 332916 305674
rect 332784 305516 332836 305522
rect 332784 305458 332836 305464
rect 332692 305448 332744 305454
rect 332692 305390 332744 305396
rect 332704 260166 332732 305390
rect 332796 265674 332824 305458
rect 332888 283626 332916 305646
rect 332968 305584 333020 305590
rect 332968 305526 333020 305532
rect 332980 286346 333008 305526
rect 333164 297430 333192 310420
rect 333256 310406 333454 310434
rect 333256 305522 333284 310406
rect 333244 305516 333296 305522
rect 333244 305458 333296 305464
rect 333624 305454 333652 310420
rect 333716 310406 333914 310434
rect 333716 305590 333744 310406
rect 334084 306474 334112 310420
rect 334268 309134 334296 310420
rect 334176 309106 334296 309134
rect 334072 306468 334124 306474
rect 334072 306410 334124 306416
rect 333980 306400 334032 306406
rect 334176 306354 334204 309106
rect 334348 306468 334400 306474
rect 334348 306410 334400 306416
rect 333980 306342 334032 306348
rect 333704 305584 333756 305590
rect 333704 305526 333756 305532
rect 333612 305448 333664 305454
rect 333612 305390 333664 305396
rect 333152 297424 333204 297430
rect 333152 297366 333204 297372
rect 332968 286340 333020 286346
rect 332968 286282 333020 286288
rect 332876 283620 332928 283626
rect 332876 283562 332928 283568
rect 332784 265668 332836 265674
rect 332784 265610 332836 265616
rect 332692 260160 332744 260166
rect 332692 260102 332744 260108
rect 333992 253298 334020 306342
rect 334084 306326 334204 306354
rect 334084 280838 334112 306326
rect 334164 306264 334216 306270
rect 334164 306206 334216 306212
rect 334176 290494 334204 306206
rect 334256 305584 334308 305590
rect 334256 305526 334308 305532
rect 334268 296002 334296 305526
rect 334360 298790 334388 306410
rect 334544 304298 334572 310420
rect 334728 306270 334756 310420
rect 334912 306406 334940 310420
rect 335004 310406 335202 310434
rect 334900 306400 334952 306406
rect 334900 306342 334952 306348
rect 334716 306264 334768 306270
rect 334716 306206 334768 306212
rect 335004 305590 335032 310406
rect 335372 306270 335400 310420
rect 335556 306320 335584 310420
rect 335832 306746 335860 310420
rect 335820 306740 335872 306746
rect 335820 306682 335872 306688
rect 336016 306626 336044 310420
rect 336096 306740 336148 306746
rect 336096 306682 336148 306688
rect 335464 306292 335584 306320
rect 335648 306598 336044 306626
rect 335360 306264 335412 306270
rect 335360 306206 335412 306212
rect 334992 305584 335044 305590
rect 334992 305526 335044 305532
rect 335360 305516 335412 305522
rect 335360 305458 335412 305464
rect 334532 304292 334584 304298
rect 334532 304234 334584 304240
rect 334348 298784 334400 298790
rect 334348 298726 334400 298732
rect 334256 295996 334308 296002
rect 334256 295938 334308 295944
rect 334164 290488 334216 290494
rect 334164 290430 334216 290436
rect 334072 280832 334124 280838
rect 334072 280774 334124 280780
rect 333980 253292 334032 253298
rect 333980 253234 334032 253240
rect 332600 251864 332652 251870
rect 332600 251806 332652 251812
rect 331312 249076 331364 249082
rect 331312 249018 331364 249024
rect 331220 246356 331272 246362
rect 331220 246298 331272 246304
rect 324320 244870 324372 244876
rect 328458 244896 328514 244905
rect 328458 244831 328514 244840
rect 335372 244798 335400 305458
rect 335464 253230 335492 306292
rect 335544 305584 335596 305590
rect 335544 305526 335596 305532
rect 335556 267034 335584 305526
rect 335648 282198 335676 306598
rect 335728 306264 335780 306270
rect 335728 306206 335780 306212
rect 335740 289134 335768 306206
rect 336108 305833 336136 306682
rect 336094 305824 336150 305833
rect 336094 305759 336150 305768
rect 336200 302234 336228 310420
rect 336292 310406 336490 310434
rect 336292 305522 336320 310406
rect 336660 305590 336688 310420
rect 336648 305584 336700 305590
rect 336648 305526 336700 305532
rect 336280 305516 336332 305522
rect 336280 305458 336332 305464
rect 335832 302206 336228 302234
rect 335832 293282 335860 302206
rect 335820 293276 335872 293282
rect 335820 293218 335872 293224
rect 335728 289128 335780 289134
rect 335728 289070 335780 289076
rect 335636 282192 335688 282198
rect 335636 282134 335688 282140
rect 335544 267028 335596 267034
rect 335544 266970 335596 266976
rect 336936 254794 336964 310420
rect 337120 300014 337148 310420
rect 337304 308310 337332 310420
rect 337292 308304 337344 308310
rect 337292 308246 337344 308252
rect 337580 308242 337608 310420
rect 337764 308417 337792 310420
rect 337750 308408 337806 308417
rect 337750 308343 337806 308352
rect 337568 308236 337620 308242
rect 337568 308178 337620 308184
rect 337948 305318 337976 310420
rect 337936 305312 337988 305318
rect 337936 305254 337988 305260
rect 338224 300558 338252 310420
rect 338408 308378 338436 310420
rect 338396 308372 338448 308378
rect 338396 308314 338448 308320
rect 338304 306400 338356 306406
rect 338304 306342 338356 306348
rect 338316 300694 338344 306342
rect 338592 305386 338620 310420
rect 338868 306377 338896 310420
rect 338854 306368 338910 306377
rect 338854 306303 338910 306312
rect 338580 305380 338632 305386
rect 338580 305322 338632 305328
rect 339052 302234 339080 310420
rect 339144 310406 339342 310434
rect 339144 306406 339172 310406
rect 339132 306400 339184 306406
rect 339132 306342 339184 306348
rect 339512 306354 339540 310420
rect 339710 310406 339908 310434
rect 339880 306490 339908 310406
rect 339972 306626 340000 310420
rect 339972 306598 340092 306626
rect 339880 306462 340000 306490
rect 339512 306326 339908 306354
rect 339684 306264 339736 306270
rect 339684 306206 339736 306212
rect 339592 305584 339644 305590
rect 339592 305526 339644 305532
rect 338408 302206 339080 302234
rect 338304 300688 338356 300694
rect 338304 300630 338356 300636
rect 338212 300552 338264 300558
rect 338212 300494 338264 300500
rect 337108 300008 337160 300014
rect 337108 299950 337160 299956
rect 338408 297906 338436 302206
rect 338396 297900 338448 297906
rect 338396 297842 338448 297848
rect 336924 254788 336976 254794
rect 336924 254730 336976 254736
rect 339604 253502 339632 305526
rect 339696 300082 339724 306206
rect 339684 300076 339736 300082
rect 339684 300018 339736 300024
rect 339592 253496 339644 253502
rect 339592 253438 339644 253444
rect 335452 253224 335504 253230
rect 335452 253166 335504 253172
rect 339880 244866 339908 306326
rect 339972 305182 340000 306462
rect 339960 305176 340012 305182
rect 339960 305118 340012 305124
rect 340064 303521 340092 306598
rect 340050 303512 340106 303521
rect 340050 303447 340106 303456
rect 340156 299946 340184 310420
rect 340340 306270 340368 310420
rect 340432 310406 340630 310434
rect 340328 306264 340380 306270
rect 340328 306206 340380 306212
rect 340432 305590 340460 310406
rect 340420 305584 340472 305590
rect 340420 305526 340472 305532
rect 340800 305114 340828 310420
rect 340788 305108 340840 305114
rect 340788 305050 340840 305056
rect 340984 302734 341012 310420
rect 341064 308644 341116 308650
rect 341064 308586 341116 308592
rect 341076 308174 341104 308586
rect 341064 308168 341116 308174
rect 341064 308110 341116 308116
rect 341156 306400 341208 306406
rect 341156 306342 341208 306348
rect 341064 306332 341116 306338
rect 341064 306274 341116 306280
rect 340972 302728 341024 302734
rect 340972 302670 341024 302676
rect 341076 300762 341104 306274
rect 341064 300756 341116 300762
rect 341064 300698 341116 300704
rect 340144 299940 340196 299946
rect 340144 299882 340196 299888
rect 341168 252074 341196 306342
rect 341260 302234 341288 310420
rect 341444 306338 341472 310420
rect 341628 306406 341656 310420
rect 341616 306400 341668 306406
rect 341616 306342 341668 306348
rect 341432 306332 341484 306338
rect 341432 306274 341484 306280
rect 341904 306202 341932 310420
rect 341892 306196 341944 306202
rect 341892 306138 341944 306144
rect 342088 302802 342116 310420
rect 342076 302796 342128 302802
rect 342076 302738 342128 302744
rect 342364 302234 342392 310420
rect 342548 306354 342576 310420
rect 342548 306326 342668 306354
rect 342732 306338 342760 310420
rect 342536 306264 342588 306270
rect 342536 306206 342588 306212
rect 341260 302206 341564 302234
rect 342364 302206 342484 302234
rect 341536 297838 341564 302206
rect 342456 300830 342484 302206
rect 342444 300824 342496 300830
rect 342444 300766 342496 300772
rect 341524 297832 341576 297838
rect 341524 297774 341576 297780
rect 341156 252068 341208 252074
rect 341156 252010 341208 252016
rect 339868 244860 339920 244866
rect 339868 244802 339920 244808
rect 335360 244792 335412 244798
rect 335360 244734 335412 244740
rect 306840 244724 306892 244730
rect 306840 244666 306892 244672
rect 342548 244662 342576 306206
rect 342640 254726 342668 306326
rect 342720 306332 342772 306338
rect 342720 306274 342772 306280
rect 343008 302870 343036 310420
rect 342996 302864 343048 302870
rect 342996 302806 343048 302812
rect 343192 300490 343220 310420
rect 343376 306270 343404 310420
rect 343652 306610 343680 310420
rect 343640 306604 343692 306610
rect 343640 306546 343692 306552
rect 343364 306264 343416 306270
rect 343364 306206 343416 306212
rect 343836 303482 343864 310420
rect 344034 310406 344232 310434
rect 344008 306604 344060 306610
rect 344008 306546 344060 306552
rect 343824 303476 343876 303482
rect 343824 303418 343876 303424
rect 343824 302252 343876 302258
rect 343824 302194 343876 302200
rect 343180 300484 343232 300490
rect 343180 300426 343232 300432
rect 342628 254720 342680 254726
rect 342628 254662 342680 254668
rect 343836 253434 343864 302194
rect 343824 253428 343876 253434
rect 343824 253370 343876 253376
rect 342536 244656 342588 244662
rect 342536 244598 342588 244604
rect 303620 244384 303672 244390
rect 300950 244352 301006 244361
rect 303620 244326 303672 244332
rect 300950 244287 301006 244296
rect 300768 243976 300820 243982
rect 300768 243918 300820 243924
rect 344020 243914 344048 306546
rect 344100 306332 344152 306338
rect 344100 306274 344152 306280
rect 344112 248266 344140 306274
rect 344204 300626 344232 310406
rect 344296 302258 344324 310420
rect 344480 306134 344508 310420
rect 344468 306128 344520 306134
rect 344468 306070 344520 306076
rect 344756 303550 344784 310420
rect 344940 306338 344968 310420
rect 345138 310406 345336 310434
rect 345204 306400 345256 306406
rect 345204 306342 345256 306348
rect 344928 306332 344980 306338
rect 344928 306274 344980 306280
rect 345020 306264 345072 306270
rect 345020 306206 345072 306212
rect 344744 303544 344796 303550
rect 344744 303486 344796 303492
rect 344284 302252 344336 302258
rect 344284 302194 344336 302200
rect 344192 300620 344244 300626
rect 344192 300562 344244 300568
rect 345032 300354 345060 306206
rect 345020 300348 345072 300354
rect 345020 300290 345072 300296
rect 344100 248260 344152 248266
rect 344100 248202 344152 248208
rect 345216 248198 345244 306342
rect 345308 306338 345336 310406
rect 345296 306332 345348 306338
rect 345296 306274 345348 306280
rect 345296 306196 345348 306202
rect 345296 306138 345348 306144
rect 345308 300529 345336 306138
rect 345294 300520 345350 300529
rect 345294 300455 345350 300464
rect 345204 248192 345256 248198
rect 345204 248134 345256 248140
rect 344008 243908 344060 243914
rect 344008 243850 344060 243856
rect 345400 243846 345428 310420
rect 345480 306332 345532 306338
rect 345480 306274 345532 306280
rect 345492 248334 345520 306274
rect 345584 303278 345612 310420
rect 345768 306406 345796 310420
rect 345860 310406 346058 310434
rect 345756 306400 345808 306406
rect 345756 306342 345808 306348
rect 345860 306270 345888 310406
rect 345848 306264 345900 306270
rect 345848 306206 345900 306212
rect 346228 306202 346256 310420
rect 346426 310406 346532 310434
rect 346216 306196 346268 306202
rect 346216 306138 346268 306144
rect 345572 303272 345624 303278
rect 345572 303214 345624 303220
rect 345480 248328 345532 248334
rect 345480 248270 345532 248276
rect 346504 246702 346532 310406
rect 346596 310406 346702 310434
rect 346596 300422 346624 310406
rect 346872 308553 346900 310420
rect 346858 308544 346914 308553
rect 346858 308479 346914 308488
rect 346584 300416 346636 300422
rect 346584 300358 346636 300364
rect 347056 296714 347084 310420
rect 347332 308990 347360 310420
rect 347320 308984 347372 308990
rect 347320 308926 347372 308932
rect 347516 308825 347544 310420
rect 347502 308816 347558 308825
rect 347502 308751 347558 308760
rect 347792 306354 347820 310420
rect 347976 308922 348004 310420
rect 347964 308916 348016 308922
rect 347964 308858 348016 308864
rect 348160 308582 348188 310420
rect 348252 310406 348450 310434
rect 348148 308576 348200 308582
rect 348148 308518 348200 308524
rect 347792 306326 348096 306354
rect 347964 306264 348016 306270
rect 347964 306206 348016 306212
rect 346872 296686 347084 296714
rect 346492 246696 346544 246702
rect 346492 246638 346544 246644
rect 345388 243840 345440 243846
rect 345388 243782 345440 243788
rect 346872 243642 346900 296686
rect 347976 248062 348004 306206
rect 347964 248056 348016 248062
rect 347964 247998 348016 248004
rect 348068 243778 348096 306326
rect 348252 306270 348280 310406
rect 348620 308854 348648 310420
rect 348608 308848 348660 308854
rect 348608 308790 348660 308796
rect 348804 308718 348832 310420
rect 348896 310406 349094 310434
rect 348792 308712 348844 308718
rect 348792 308654 348844 308660
rect 348240 306264 348292 306270
rect 348240 306206 348292 306212
rect 348896 296714 348924 310406
rect 349264 306354 349292 310420
rect 349448 309126 349476 310420
rect 349632 310406 349738 310434
rect 349436 309120 349488 309126
rect 349436 309062 349488 309068
rect 349264 306326 349568 306354
rect 349344 306264 349396 306270
rect 349344 306206 349396 306212
rect 349252 306196 349304 306202
rect 349252 306138 349304 306144
rect 348344 296686 348924 296714
rect 348344 247994 348372 296686
rect 348332 247988 348384 247994
rect 348332 247930 348384 247936
rect 349264 246566 349292 306138
rect 349356 300150 349384 306206
rect 349436 306128 349488 306134
rect 349436 306070 349488 306076
rect 349344 300144 349396 300150
rect 349344 300086 349396 300092
rect 349448 246634 349476 306070
rect 349540 300218 349568 306326
rect 349632 306202 349660 310406
rect 349908 306270 349936 310420
rect 350184 308514 350212 310420
rect 350172 308508 350224 308514
rect 350172 308450 350224 308456
rect 349896 306264 349948 306270
rect 349896 306206 349948 306212
rect 349620 306196 349672 306202
rect 349620 306138 349672 306144
rect 350368 306134 350396 310420
rect 350566 310406 350672 310434
rect 350356 306128 350408 306134
rect 350356 306070 350408 306076
rect 350644 305998 350672 310406
rect 350828 309058 350856 310420
rect 350816 309052 350868 309058
rect 350816 308994 350868 309000
rect 351012 308394 351040 310420
rect 350724 308372 350776 308378
rect 350724 308314 350776 308320
rect 350920 308366 351040 308394
rect 350632 305992 350684 305998
rect 350632 305934 350684 305940
rect 350736 300801 350764 308314
rect 350722 300792 350778 300801
rect 350722 300727 350778 300736
rect 349528 300212 349580 300218
rect 349528 300154 349580 300160
rect 350920 248130 350948 308366
rect 351000 308304 351052 308310
rect 351000 308246 351052 308252
rect 351012 265878 351040 308246
rect 351196 306066 351224 310420
rect 351288 310406 351486 310434
rect 351288 308310 351316 310406
rect 351656 308514 351684 310420
rect 351644 308508 351696 308514
rect 351644 308450 351696 308456
rect 351840 308378 351868 310420
rect 352116 308689 352144 310420
rect 352102 308680 352158 308689
rect 352102 308615 352158 308624
rect 352300 308582 352328 310420
rect 352288 308576 352340 308582
rect 352288 308518 352340 308524
rect 351828 308372 351880 308378
rect 351828 308314 351880 308320
rect 352012 308372 352064 308378
rect 352012 308314 352064 308320
rect 351276 308304 351328 308310
rect 351276 308246 351328 308252
rect 351184 306060 351236 306066
rect 351184 306002 351236 306008
rect 352024 305930 352052 308314
rect 352012 305924 352064 305930
rect 352012 305866 352064 305872
rect 352484 300286 352512 310420
rect 352576 310406 352774 310434
rect 352576 308378 352604 310406
rect 352944 308718 352972 310420
rect 353220 308786 353248 310420
rect 353208 308780 353260 308786
rect 353208 308722 353260 308728
rect 352932 308712 352984 308718
rect 352932 308654 352984 308660
rect 353404 308394 353432 310420
rect 353588 308650 353616 310420
rect 353576 308644 353628 308650
rect 353576 308586 353628 308592
rect 352564 308372 352616 308378
rect 353404 308366 353800 308394
rect 352564 308314 352616 308320
rect 353668 308304 353720 308310
rect 353668 308246 353720 308252
rect 353392 308236 353444 308242
rect 353392 308178 353444 308184
rect 353404 305794 353432 308178
rect 353392 305788 353444 305794
rect 353392 305730 353444 305736
rect 353680 305726 353708 308246
rect 353772 305862 353800 308366
rect 353864 308174 353892 310420
rect 354048 308242 354076 310420
rect 354232 308854 354260 310420
rect 354324 310406 354522 310434
rect 354220 308848 354272 308854
rect 354220 308790 354272 308796
rect 354324 308310 354352 310406
rect 354692 308786 354720 310420
rect 354876 309126 354904 310420
rect 354968 310406 355166 310434
rect 354864 309120 354916 309126
rect 354864 309062 354916 309068
rect 354680 308780 354732 308786
rect 354680 308722 354732 308728
rect 354968 308666 354996 310406
rect 354692 308638 354996 308666
rect 354312 308304 354364 308310
rect 354312 308246 354364 308252
rect 354036 308236 354088 308242
rect 354036 308178 354088 308184
rect 353852 308168 353904 308174
rect 353852 308110 353904 308116
rect 353760 305856 353812 305862
rect 353760 305798 353812 305804
rect 353668 305720 353720 305726
rect 353668 305662 353720 305668
rect 354692 303618 354720 308638
rect 355336 308394 355364 310420
rect 355612 308854 355640 310420
rect 355600 308848 355652 308854
rect 355600 308790 355652 308796
rect 355416 308780 355468 308786
rect 355416 308722 355468 308728
rect 354876 308366 355364 308394
rect 354772 308032 354824 308038
rect 354772 307974 354824 307980
rect 354680 303612 354732 303618
rect 354680 303554 354732 303560
rect 354784 300665 354812 307974
rect 354876 303385 354904 308366
rect 355140 308304 355192 308310
rect 355140 308246 355192 308252
rect 354862 303376 354918 303385
rect 354862 303311 354918 303320
rect 354770 300656 354826 300665
rect 354770 300591 354826 300600
rect 352472 300280 352524 300286
rect 352472 300222 352524 300228
rect 351000 265872 351052 265878
rect 351000 265814 351052 265820
rect 355152 250646 355180 308246
rect 355428 306241 355456 308722
rect 355796 308038 355824 310420
rect 355980 308310 356008 310420
rect 356256 308786 356284 310420
rect 356244 308780 356296 308786
rect 356244 308722 356296 308728
rect 356440 308530 356468 310420
rect 356520 308780 356572 308786
rect 356520 308722 356572 308728
rect 356256 308502 356468 308530
rect 356060 308372 356112 308378
rect 356060 308314 356112 308320
rect 355968 308304 356020 308310
rect 355968 308246 356020 308252
rect 355784 308032 355836 308038
rect 355784 307974 355836 307980
rect 355414 306232 355470 306241
rect 355414 306167 355470 306176
rect 356072 303414 356100 308314
rect 356152 308304 356204 308310
rect 356152 308246 356204 308252
rect 356060 303408 356112 303414
rect 356060 303350 356112 303356
rect 356164 303346 356192 308246
rect 356152 303340 356204 303346
rect 356152 303282 356204 303288
rect 356256 297974 356284 308502
rect 356532 308292 356560 308722
rect 356624 308378 356652 310420
rect 356716 310406 356914 310434
rect 356612 308372 356664 308378
rect 356612 308314 356664 308320
rect 356440 308264 356560 308292
rect 356336 308168 356388 308174
rect 356336 308110 356388 308116
rect 356348 298042 356376 308110
rect 356336 298036 356388 298042
rect 356336 297978 356388 297984
rect 356244 297968 356296 297974
rect 356244 297910 356296 297916
rect 355140 250640 355192 250646
rect 355140 250582 355192 250588
rect 356440 248130 356468 308264
rect 356716 296714 356744 310406
rect 357084 308174 357112 310420
rect 357268 308310 357296 310420
rect 357440 308780 357492 308786
rect 357440 308722 357492 308728
rect 357256 308304 357308 308310
rect 357256 308246 357308 308252
rect 357072 308168 357124 308174
rect 357072 308110 357124 308116
rect 357452 303142 357480 308722
rect 357544 308292 357572 310420
rect 357728 308394 357756 310420
rect 357912 308786 357940 310420
rect 358004 310406 358202 310434
rect 357900 308780 357952 308786
rect 357900 308722 357952 308728
rect 357728 308366 357940 308394
rect 357808 308304 357860 308310
rect 357544 308264 357756 308292
rect 357624 308168 357676 308174
rect 357624 308110 357676 308116
rect 357532 308100 357584 308106
rect 357532 308042 357584 308048
rect 357544 303210 357572 308042
rect 357532 303204 357584 303210
rect 357532 303146 357584 303152
rect 357440 303136 357492 303142
rect 357440 303078 357492 303084
rect 356532 296686 356744 296714
rect 350908 248124 350960 248130
rect 350908 248066 350960 248072
rect 356428 248124 356480 248130
rect 356428 248066 356480 248072
rect 349436 246628 349488 246634
rect 349436 246570 349488 246576
rect 349252 246560 349304 246566
rect 349252 246502 349304 246508
rect 356532 244798 356560 296686
rect 357636 245614 357664 308110
rect 357728 248062 357756 308264
rect 357808 308246 357860 308252
rect 357716 248056 357768 248062
rect 357716 247998 357768 248004
rect 357624 245608 357676 245614
rect 357624 245550 357676 245556
rect 356520 244792 356572 244798
rect 356520 244734 356572 244740
rect 348056 243772 348108 243778
rect 348056 243714 348108 243720
rect 346860 243636 346912 243642
rect 346860 243578 346912 243584
rect 357820 243574 357848 308246
rect 357912 243710 357940 308366
rect 358004 308174 358032 310406
rect 358372 308310 358400 310420
rect 358464 310406 358662 310434
rect 358360 308304 358412 308310
rect 358360 308246 358412 308252
rect 357992 308168 358044 308174
rect 357992 308110 358044 308116
rect 358464 308106 358492 310406
rect 358832 308174 358860 310420
rect 359030 310406 359136 310434
rect 358912 308372 358964 308378
rect 358912 308314 358964 308320
rect 358820 308168 358872 308174
rect 358820 308110 358872 308116
rect 358452 308100 358504 308106
rect 358452 308042 358504 308048
rect 358820 307964 358872 307970
rect 358820 307906 358872 307912
rect 358832 305658 358860 307906
rect 358820 305652 358872 305658
rect 358820 305594 358872 305600
rect 358924 303006 358952 308314
rect 359004 308304 359056 308310
rect 359004 308246 359056 308252
rect 358912 303000 358964 303006
rect 358912 302942 358964 302948
rect 359016 248198 359044 308246
rect 359108 297702 359136 310406
rect 359292 308258 359320 310420
rect 359292 308230 359412 308258
rect 359280 308168 359332 308174
rect 359280 308110 359332 308116
rect 359188 308100 359240 308106
rect 359188 308042 359240 308048
rect 359096 297696 359148 297702
rect 359096 297638 359148 297644
rect 359004 248192 359056 248198
rect 359004 248134 359056 248140
rect 359200 244866 359228 308042
rect 359292 247994 359320 308110
rect 359384 303074 359412 308230
rect 359476 308106 359504 310420
rect 359464 308100 359516 308106
rect 359464 308042 359516 308048
rect 359660 307970 359688 310420
rect 359752 310406 359950 310434
rect 359752 308378 359780 310406
rect 359740 308372 359792 308378
rect 359740 308314 359792 308320
rect 360120 308310 360148 310420
rect 360108 308304 360160 308310
rect 360108 308246 360160 308252
rect 359648 307964 359700 307970
rect 359648 307906 359700 307912
rect 359372 303068 359424 303074
rect 359372 303010 359424 303016
rect 360304 297770 360332 310420
rect 360580 302938 360608 310420
rect 360568 302932 360620 302938
rect 360568 302874 360620 302880
rect 360292 297764 360344 297770
rect 360292 297706 360344 297712
rect 360764 296714 360792 310420
rect 360948 305697 360976 442734
rect 361040 442270 361068 446150
rect 361028 442264 361080 442270
rect 361028 442206 361080 442212
rect 362236 325650 362264 446354
rect 364984 446344 365036 446350
rect 364984 446286 365036 446292
rect 363604 446276 363656 446282
rect 363604 446218 363656 446224
rect 362316 443624 362368 443630
rect 362316 443566 362368 443572
rect 362328 431934 362356 443566
rect 362316 431928 362368 431934
rect 362316 431870 362368 431876
rect 362224 325644 362276 325650
rect 362224 325586 362276 325592
rect 360934 305688 360990 305697
rect 360934 305623 360990 305632
rect 360396 296686 360792 296714
rect 359280 247988 359332 247994
rect 359280 247930 359332 247936
rect 359188 244860 359240 244866
rect 359188 244802 359240 244808
rect 360396 244730 360424 296686
rect 363616 258738 363644 446218
rect 364996 260234 365024 446286
rect 373264 446140 373316 446146
rect 373264 446082 373316 446088
rect 369124 444440 369176 444446
rect 369124 444382 369176 444388
rect 367744 443556 367796 443562
rect 367744 443498 367796 443504
rect 367756 273222 367784 443498
rect 369136 379506 369164 444382
rect 369124 379500 369176 379506
rect 369124 379442 369176 379448
rect 367744 273216 367796 273222
rect 367744 273158 367796 273164
rect 364984 260228 365036 260234
rect 364984 260170 365036 260176
rect 363604 258732 363656 258738
rect 363604 258674 363656 258680
rect 373276 257378 373304 446082
rect 458824 445800 458876 445806
rect 458824 445742 458876 445748
rect 442264 444848 442316 444854
rect 442264 444790 442316 444796
rect 438124 308916 438176 308922
rect 438124 308858 438176 308864
rect 436836 308848 436888 308854
rect 436836 308790 436888 308796
rect 373264 257372 373316 257378
rect 373264 257314 373316 257320
rect 436744 253360 436796 253366
rect 436744 253302 436796 253308
rect 360384 244724 360436 244730
rect 360384 244666 360436 244672
rect 357900 243704 357952 243710
rect 357900 243646 357952 243652
rect 357808 243568 357860 243574
rect 357808 243510 357860 243516
rect 299386 168056 299442 168065
rect 299386 167991 299442 168000
rect 299386 167104 299442 167113
rect 299386 167039 299442 167048
rect 299296 159656 299348 159662
rect 299296 159598 299348 159604
rect 299296 158568 299348 158574
rect 299296 158510 299348 158516
rect 299308 157962 299336 158510
rect 299296 157956 299348 157962
rect 299296 157898 299348 157904
rect 299204 157616 299256 157622
rect 299204 157558 299256 157564
rect 299112 157548 299164 157554
rect 299112 157490 299164 157496
rect 298928 155916 298980 155922
rect 298928 155858 298980 155864
rect 299296 154488 299348 154494
rect 299296 154430 299348 154436
rect 299308 153746 299336 154430
rect 299296 153740 299348 153746
rect 299296 153682 299348 153688
rect 299400 4826 299428 167039
rect 345938 159896 345994 159905
rect 345938 159831 345994 159840
rect 348238 159896 348294 159905
rect 348238 159831 348294 159840
rect 353574 159896 353630 159905
rect 353574 159831 353630 159840
rect 365902 159896 365958 159905
rect 365902 159831 365958 159840
rect 299480 159588 299532 159594
rect 299480 159530 299532 159536
rect 299388 4820 299440 4826
rect 299388 4762 299440 4768
rect 298744 3936 298796 3942
rect 298744 3878 298796 3884
rect 299492 2774 299520 159530
rect 313280 159520 313332 159526
rect 313280 159462 313332 159468
rect 299570 158672 299626 158681
rect 299570 158607 299626 158616
rect 299584 158574 299612 158607
rect 299572 158568 299624 158574
rect 299572 158510 299624 158516
rect 302240 156732 302292 156738
rect 302240 156674 302292 156680
rect 299572 152652 299624 152658
rect 299572 152594 299624 152600
rect 299584 7614 299612 152594
rect 300858 151056 300914 151065
rect 300858 150991 300914 151000
rect 300872 16574 300900 150991
rect 302252 16574 302280 156674
rect 306380 155168 306432 155174
rect 306380 155110 306432 155116
rect 303620 147076 303672 147082
rect 303620 147018 303672 147024
rect 303632 16574 303660 147018
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 299572 7608 299624 7614
rect 299572 7550 299624 7556
rect 300768 7608 300820 7614
rect 300768 7550 300820 7556
rect 299492 2746 299704 2774
rect 299676 480 299704 2746
rect 300780 480 300808 7550
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305552 14476 305604 14482
rect 305552 14418 305604 14424
rect 305564 480 305592 14418
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 155110
rect 309138 153776 309194 153785
rect 309138 153711 309194 153720
rect 309152 16574 309180 153711
rect 310520 145648 310572 145654
rect 310520 145590 310572 145596
rect 310532 16574 310560 145590
rect 313292 16574 313320 159462
rect 320180 159452 320232 159458
rect 320180 159394 320232 159400
rect 316038 158672 316094 158681
rect 316038 158607 316094 158616
rect 316682 158672 316738 158681
rect 316682 158607 316738 158616
rect 319442 158672 319498 158681
rect 319442 158607 319498 158616
rect 316052 156806 316080 158607
rect 316040 156800 316092 156806
rect 316040 156742 316092 156748
rect 316040 156596 316092 156602
rect 316040 156538 316092 156544
rect 314660 144288 314712 144294
rect 314660 144230 314712 144236
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 313292 16546 313872 16574
rect 307944 5160 307996 5166
rect 307944 5102 307996 5108
rect 307956 480 307984 5102
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 312176 13116 312228 13122
rect 312176 13058 312228 13064
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 13058
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 144230
rect 316052 3398 316080 156538
rect 316696 156534 316724 158607
rect 319456 158166 319484 158607
rect 319444 158160 319496 158166
rect 319444 158102 319496 158108
rect 320088 157820 320140 157826
rect 320088 157762 320140 157768
rect 317694 157448 317750 157457
rect 317694 157383 317750 157392
rect 316684 156528 316736 156534
rect 316684 156470 316736 156476
rect 317708 154154 317736 157383
rect 320100 155922 320128 157762
rect 320088 155916 320140 155922
rect 320088 155858 320140 155864
rect 317696 154148 317748 154154
rect 317696 154090 317748 154096
rect 317420 149864 317472 149870
rect 317420 149806 317472 149812
rect 317432 16574 317460 149806
rect 318800 130416 318852 130422
rect 318800 130358 318852 130364
rect 318812 16574 318840 130358
rect 320192 16574 320220 159394
rect 345952 159390 345980 159831
rect 345940 159384 345992 159390
rect 345940 159326 345992 159332
rect 348252 159254 348280 159831
rect 350998 159760 351054 159769
rect 350998 159695 351054 159704
rect 351012 159322 351040 159695
rect 351000 159316 351052 159322
rect 351000 159258 351052 159264
rect 348240 159248 348292 159254
rect 348240 159190 348292 159196
rect 353588 158982 353616 159831
rect 356058 159624 356114 159633
rect 356058 159559 356114 159568
rect 358450 159624 358506 159633
rect 358450 159559 358506 159568
rect 356072 159186 356100 159559
rect 356060 159180 356112 159186
rect 356060 159122 356112 159128
rect 358464 159118 358492 159559
rect 358452 159112 358504 159118
rect 358452 159054 358504 159060
rect 365916 159050 365944 159831
rect 373998 159352 374054 159361
rect 373998 159287 374054 159296
rect 365904 159044 365956 159050
rect 365904 158986 365956 158992
rect 353576 158976 353628 158982
rect 353576 158918 353628 158924
rect 368204 158908 368256 158914
rect 368204 158850 368256 158856
rect 360844 158840 360896 158846
rect 360844 158782 360896 158788
rect 338396 158704 338448 158710
rect 320546 158672 320602 158681
rect 320546 158607 320602 158616
rect 323122 158672 323178 158681
rect 323122 158607 323178 158616
rect 324226 158672 324282 158681
rect 324226 158607 324282 158616
rect 326434 158672 326490 158681
rect 326434 158607 326490 158616
rect 328274 158672 328330 158681
rect 328274 158607 328276 158616
rect 320560 158506 320588 158607
rect 320548 158500 320600 158506
rect 320548 158442 320600 158448
rect 323136 157214 323164 158607
rect 324240 157282 324268 158607
rect 325146 157992 325202 158001
rect 325146 157927 325202 157936
rect 325160 157826 325188 157927
rect 326448 157894 326476 158607
rect 328328 158607 328330 158616
rect 328642 158672 328698 158681
rect 328642 158607 328698 158616
rect 329930 158672 329986 158681
rect 329930 158607 329986 158616
rect 330482 158672 330538 158681
rect 330482 158607 330538 158616
rect 332230 158672 332286 158681
rect 332230 158607 332286 158616
rect 333610 158672 333666 158681
rect 333610 158607 333666 158616
rect 334530 158672 334586 158681
rect 334530 158607 334586 158616
rect 335634 158672 335690 158681
rect 335634 158607 335690 158616
rect 336002 158672 336058 158681
rect 336002 158607 336058 158616
rect 336830 158672 336886 158681
rect 336830 158607 336886 158616
rect 338394 158672 338396 158681
rect 360856 158681 360884 158782
rect 363420 158772 363472 158778
rect 363420 158714 363472 158720
rect 363432 158681 363460 158714
rect 368216 158681 368244 158850
rect 371056 158704 371108 158710
rect 338448 158672 338450 158681
rect 338394 158607 338450 158616
rect 338762 158672 338818 158681
rect 338762 158607 338818 158616
rect 340970 158672 341026 158681
rect 340970 158607 341026 158616
rect 343546 158672 343602 158681
rect 343546 158607 343602 158616
rect 349802 158672 349858 158681
rect 349802 158607 349858 158616
rect 355230 158672 355286 158681
rect 355230 158607 355286 158616
rect 356978 158672 357034 158681
rect 356978 158607 357034 158616
rect 360842 158672 360898 158681
rect 360842 158607 360898 158616
rect 363418 158672 363474 158681
rect 363418 158607 363474 158616
rect 368202 158672 368258 158681
rect 368202 158607 368258 158616
rect 371054 158672 371056 158681
rect 371108 158672 371110 158681
rect 371054 158607 371110 158616
rect 373446 158672 373502 158681
rect 373446 158607 373448 158616
rect 328276 158578 328328 158584
rect 328656 158234 328684 158607
rect 328644 158228 328696 158234
rect 328644 158170 328696 158176
rect 329944 157962 329972 158607
rect 330496 158030 330524 158607
rect 332244 158574 332272 158607
rect 332232 158568 332284 158574
rect 332232 158510 332284 158516
rect 333624 158302 333652 158607
rect 333612 158296 333664 158302
rect 333612 158238 333664 158244
rect 330484 158024 330536 158030
rect 330484 157966 330536 157972
rect 329932 157956 329984 157962
rect 329932 157898 329984 157904
rect 326436 157888 326488 157894
rect 326436 157830 326488 157836
rect 325148 157820 325200 157826
rect 325148 157762 325200 157768
rect 329196 157480 329248 157486
rect 329196 157422 329248 157428
rect 327356 157412 327408 157418
rect 327356 157354 327408 157360
rect 324228 157276 324280 157282
rect 324228 157218 324280 157224
rect 323124 157208 323176 157214
rect 323124 157150 323176 157156
rect 327080 156664 327132 156670
rect 327080 156606 327132 156612
rect 324320 155372 324372 155378
rect 324320 155314 324372 155320
rect 321560 142860 321612 142866
rect 321560 142802 321612 142808
rect 321572 16574 321600 142802
rect 322940 17264 322992 17270
rect 322940 17206 322992 17212
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 11756 316276 11762
rect 316224 11698 316276 11704
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 11698
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 17206
rect 324332 3210 324360 155314
rect 324412 141432 324464 141438
rect 324412 141374 324464 141380
rect 324424 3398 324452 141374
rect 325700 129056 325752 129062
rect 325700 128998 325752 129004
rect 325712 16574 325740 128998
rect 327092 16574 327120 156606
rect 327368 154222 327396 157354
rect 329208 154290 329236 157422
rect 334544 157078 334572 158607
rect 334532 157072 334584 157078
rect 334532 157014 334584 157020
rect 335648 157010 335676 158607
rect 336016 158098 336044 158607
rect 336004 158092 336056 158098
rect 336004 158034 336056 158040
rect 335636 157004 335688 157010
rect 335636 156946 335688 156952
rect 336844 156942 336872 158607
rect 338118 158400 338174 158409
rect 338118 158335 338174 158344
rect 336832 156936 336884 156942
rect 336832 156878 336884 156884
rect 338132 156874 338160 158335
rect 338776 157146 338804 158607
rect 340984 158370 341012 158607
rect 343560 158438 343588 158607
rect 343548 158432 343600 158438
rect 343548 158374 343600 158380
rect 340972 158364 341024 158370
rect 340972 158306 341024 158312
rect 343914 158264 343970 158273
rect 343914 158199 343970 158208
rect 348698 158264 348754 158273
rect 348698 158199 348754 158208
rect 339498 157856 339554 157865
rect 339498 157791 339554 157800
rect 341154 157856 341210 157865
rect 341154 157791 341210 157800
rect 342810 157856 342866 157865
rect 342810 157791 342866 157800
rect 338764 157140 338816 157146
rect 338764 157082 338816 157088
rect 338120 156868 338172 156874
rect 338120 156810 338172 156816
rect 339512 155106 339540 157791
rect 341168 155514 341196 157791
rect 341156 155508 341208 155514
rect 341156 155450 341208 155456
rect 342824 155446 342852 157791
rect 343928 155718 343956 158199
rect 346398 157992 346454 158001
rect 346398 157927 346454 157936
rect 345110 157856 345166 157865
rect 345110 157791 345166 157800
rect 343916 155712 343968 155718
rect 343916 155654 343968 155660
rect 345124 155650 345152 157791
rect 346412 155854 346440 157927
rect 346858 157856 346914 157865
rect 346858 157791 346914 157800
rect 346400 155848 346452 155854
rect 346400 155790 346452 155796
rect 345112 155644 345164 155650
rect 345112 155586 345164 155592
rect 346872 155582 346900 157791
rect 348712 155786 348740 158199
rect 349816 157350 349844 158607
rect 353298 158264 353354 158273
rect 353298 158199 353354 158208
rect 351090 157448 351146 157457
rect 351090 157383 351146 157392
rect 352194 157448 352250 157457
rect 352194 157383 352250 157392
rect 349804 157344 349856 157350
rect 349804 157286 349856 157292
rect 348700 155780 348752 155786
rect 348700 155722 348752 155728
rect 346860 155576 346912 155582
rect 346860 155518 346912 155524
rect 342812 155440 342864 155446
rect 342812 155382 342864 155388
rect 340880 155304 340932 155310
rect 340880 155246 340932 155252
rect 339500 155100 339552 155106
rect 339500 155042 339552 155048
rect 329196 154284 329248 154290
rect 329196 154226 329248 154232
rect 327356 154216 327408 154222
rect 327356 154158 327408 154164
rect 331220 153876 331272 153882
rect 331220 153818 331272 153824
rect 328460 147008 328512 147014
rect 328460 146950 328512 146956
rect 328472 16574 328500 146950
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 15904 330444 15910
rect 330392 15846 330444 15852
rect 330404 480 330432 15846
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 153818
rect 333980 152584 334032 152590
rect 333980 152526 334032 152532
rect 332600 145580 332652 145586
rect 332600 145522 332652 145528
rect 332612 3210 332640 145522
rect 332692 127628 332744 127634
rect 332692 127570 332744 127576
rect 332704 3398 332732 127570
rect 333992 16574 334020 152526
rect 338120 151088 338172 151094
rect 338120 151030 338172 151036
rect 336740 149796 336792 149802
rect 336740 149738 336792 149744
rect 335360 140072 335412 140078
rect 335360 140014 335412 140020
rect 335372 16574 335400 140014
rect 336752 16574 336780 149738
rect 338132 16574 338160 151030
rect 339500 138712 339552 138718
rect 339500 138654 339552 138660
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 332692 3392 332744 3398
rect 332692 3334 332744 3340
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 332612 3182 332732 3210
rect 332704 480 332732 3182
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 138654
rect 340892 3398 340920 155246
rect 350540 155236 350592 155242
rect 350540 155178 350592 155184
rect 343640 152516 343692 152522
rect 343640 152458 343692 152464
rect 342260 144220 342312 144226
rect 342260 144162 342312 144168
rect 340972 126268 341024 126274
rect 340972 126210 341024 126216
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 340984 480 341012 126210
rect 342272 16574 342300 144162
rect 343652 16574 343680 152458
rect 345020 149728 345072 149734
rect 345020 149670 345072 149676
rect 345032 16574 345060 149670
rect 346400 137284 346452 137290
rect 346400 137226 346452 137232
rect 346412 16574 346440 137226
rect 347780 24132 347832 24138
rect 347780 24074 347832 24080
rect 347792 16574 347820 24074
rect 350552 16574 350580 155178
rect 351104 154562 351132 157383
rect 351092 154556 351144 154562
rect 351092 154498 351144 154504
rect 352208 154426 352236 157383
rect 353312 154494 353340 158199
rect 355244 157486 355272 158607
rect 355232 157480 355284 157486
rect 354402 157448 354458 157457
rect 355232 157422 355284 157428
rect 356992 157418 357020 158607
rect 373500 158607 373502 158616
rect 373448 158578 373500 158584
rect 354402 157383 354458 157392
rect 356980 157412 357032 157418
rect 353300 154488 353352 154494
rect 353300 154430 353352 154436
rect 352196 154420 352248 154426
rect 352196 154362 352248 154368
rect 354416 154358 354444 157383
rect 356980 157354 357032 157360
rect 354404 154352 354456 154358
rect 354404 154294 354456 154300
rect 357440 148368 357492 148374
rect 357440 148310 357492 148316
rect 354680 124908 354732 124914
rect 354680 124850 354732 124856
rect 354692 16574 354720 124850
rect 357452 16574 357480 148310
rect 360200 146940 360252 146946
rect 360200 146882 360252 146888
rect 360212 16574 360240 146882
rect 361580 18624 361632 18630
rect 361580 18566 361632 18572
rect 361592 16574 361620 18566
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 354692 16546 355272 16574
rect 357452 16546 357572 16574
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 350448 5092 350500 5098
rect 350448 5034 350500 5040
rect 349252 4140 349304 4146
rect 349252 4082 349304 4088
rect 349264 480 349292 4082
rect 350460 480 350488 5034
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 354036 5024 354088 5030
rect 354036 4966 354088 4972
rect 352840 4072 352892 4078
rect 352840 4014 352892 4020
rect 352852 480 352880 4014
rect 354048 480 354076 4966
rect 355244 480 355272 16546
rect 356336 4004 356388 4010
rect 356336 3946 356388 3952
rect 356348 480 356376 3946
rect 357544 480 357572 16546
rect 358728 6792 358780 6798
rect 358728 6734 358780 6740
rect 358740 480 358768 6734
rect 359924 3868 359976 3874
rect 359924 3810 359976 3816
rect 359936 480 359964 3810
rect 361132 480 361160 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 372894 6896 372950 6905
rect 372894 6831 372950 6840
rect 369398 6080 369454 6089
rect 369398 6015 369454 6024
rect 368202 4992 368258 5001
rect 364616 4956 364668 4962
rect 368202 4927 368258 4936
rect 364616 4898 364668 4904
rect 363510 3224 363566 3233
rect 363510 3159 363566 3168
rect 363524 480 363552 3159
rect 364628 480 364656 4898
rect 365812 3936 365864 3942
rect 365812 3878 365864 3884
rect 365824 480 365852 3878
rect 367008 3800 367060 3806
rect 367008 3742 367060 3748
rect 367020 480 367048 3742
rect 368216 480 368244 4927
rect 369412 480 369440 6015
rect 371700 4888 371752 4894
rect 370594 4856 370650 4865
rect 371700 4830 371752 4836
rect 370594 4791 370650 4800
rect 370608 480 370636 4791
rect 371712 480 371740 4830
rect 372908 480 372936 6831
rect 374012 3398 374040 159287
rect 393504 158772 393556 158778
rect 393504 158714 393556 158720
rect 393516 158681 393544 158714
rect 376022 158672 376078 158681
rect 376022 158607 376078 158616
rect 378598 158672 378654 158681
rect 378598 158607 378654 158616
rect 380990 158672 381046 158681
rect 380990 158607 381046 158616
rect 383566 158672 383622 158681
rect 383566 158607 383622 158616
rect 385958 158672 386014 158681
rect 385958 158607 386014 158616
rect 388534 158672 388590 158681
rect 388534 158607 388590 158616
rect 391478 158672 391534 158681
rect 391478 158607 391534 158616
rect 393502 158672 393558 158681
rect 393502 158607 393558 158616
rect 395894 158672 395950 158681
rect 395894 158607 395950 158616
rect 398470 158672 398526 158681
rect 398470 158607 398526 158616
rect 401414 158672 401470 158681
rect 401414 158607 401470 158616
rect 403806 158672 403862 158681
rect 403806 158607 403862 158616
rect 406750 158672 406806 158681
rect 406750 158607 406806 158616
rect 376036 158574 376064 158607
rect 376024 158568 376076 158574
rect 376024 158510 376076 158516
rect 378612 158506 378640 158607
rect 378600 158500 378652 158506
rect 378600 158442 378652 158448
rect 381004 158438 381032 158607
rect 380992 158432 381044 158438
rect 380992 158374 381044 158380
rect 383580 158370 383608 158607
rect 383568 158364 383620 158370
rect 383568 158306 383620 158312
rect 385972 158302 386000 158607
rect 385960 158296 386012 158302
rect 385960 158238 386012 158244
rect 388548 158234 388576 158607
rect 388536 158228 388588 158234
rect 388536 158170 388588 158176
rect 391492 158166 391520 158607
rect 391480 158160 391532 158166
rect 391480 158102 391532 158108
rect 395908 158098 395936 158607
rect 395896 158092 395948 158098
rect 395896 158034 395948 158040
rect 398484 158030 398512 158607
rect 398472 158024 398524 158030
rect 398472 157966 398524 157972
rect 401428 157962 401456 158607
rect 401416 157956 401468 157962
rect 401416 157898 401468 157904
rect 403820 157894 403848 158607
rect 403808 157888 403860 157894
rect 403808 157830 403860 157836
rect 406764 157826 406792 158607
rect 406752 157820 406804 157826
rect 406752 157762 406804 157768
rect 375378 75168 375434 75177
rect 375378 75103 375434 75112
rect 375392 16574 375420 75103
rect 375392 16546 376064 16574
rect 374090 9616 374146 9625
rect 374090 9551 374146 9560
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 9551
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 387154 9480 387210 9489
rect 387154 9415 387210 9424
rect 379978 8800 380034 8809
rect 379978 8735 380034 8744
rect 378876 6724 378928 6730
rect 378876 6666 378928 6672
rect 377680 4820 377732 4826
rect 377680 4762 377732 4768
rect 377692 480 377720 4762
rect 378888 480 378916 6666
rect 379992 480 380020 8735
rect 382370 6760 382426 6769
rect 382370 6695 382426 6704
rect 381174 4040 381230 4049
rect 381174 3975 381230 3984
rect 381188 480 381216 3975
rect 382384 480 382412 6695
rect 385960 6656 386012 6662
rect 385960 6598 386012 6604
rect 383566 3904 383622 3913
rect 383566 3839 383622 3848
rect 383580 480 383608 3839
rect 384764 3732 384816 3738
rect 384764 3674 384816 3680
rect 384776 480 384804 3674
rect 385972 480 386000 6598
rect 387168 480 387196 9415
rect 394238 9344 394294 9353
rect 394238 9279 394294 9288
rect 389454 6624 389510 6633
rect 389454 6559 389510 6568
rect 388258 3768 388314 3777
rect 388258 3703 388314 3712
rect 388272 480 388300 3703
rect 389468 480 389496 6559
rect 393042 6488 393098 6497
rect 393042 6423 393098 6432
rect 390650 6352 390706 6361
rect 390650 6287 390706 6296
rect 390664 480 390692 6287
rect 391846 3632 391902 3641
rect 391846 3567 391902 3576
rect 391860 480 391888 3567
rect 393056 480 393084 6423
rect 394252 480 394280 9279
rect 408406 9208 408462 9217
rect 408406 9143 408462 9152
rect 397734 9072 397790 9081
rect 397734 9007 397790 9016
rect 396538 6216 396594 6225
rect 396538 6151 396594 6160
rect 395342 3496 395398 3505
rect 395342 3431 395398 3440
rect 395356 480 395384 3431
rect 396552 480 396580 6151
rect 397748 480 397776 9007
rect 404818 8936 404874 8945
rect 404818 8871 404874 8880
rect 400128 6588 400180 6594
rect 400128 6530 400180 6536
rect 398930 3360 398986 3369
rect 398930 3295 398986 3304
rect 398944 480 398972 3295
rect 400140 480 400168 6530
rect 403624 6520 403676 6526
rect 403624 6462 403676 6468
rect 402520 3664 402572 3670
rect 402520 3606 402572 3612
rect 401324 3460 401376 3466
rect 401324 3402 401376 3408
rect 401336 480 401364 3402
rect 402532 480 402560 3606
rect 403636 480 403664 6462
rect 404832 480 404860 8871
rect 407212 6384 407264 6390
rect 407212 6326 407264 6332
rect 406016 3596 406068 3602
rect 406016 3538 406068 3544
rect 406028 480 406056 3538
rect 407224 480 407252 6326
rect 408420 480 408448 9143
rect 410800 9104 410852 9110
rect 410800 9046 410852 9052
rect 409604 3528 409656 3534
rect 409604 3470 409656 3476
rect 409616 480 409644 3470
rect 410812 480 410840 9046
rect 411904 9036 411956 9042
rect 411904 8978 411956 8984
rect 411916 480 411944 8978
rect 414296 8968 414348 8974
rect 414296 8910 414348 8916
rect 413100 6452 413152 6458
rect 413100 6394 413152 6400
rect 413112 480 413140 6394
rect 414308 480 414336 8910
rect 416688 6316 416740 6322
rect 416688 6258 416740 6264
rect 415492 6180 415544 6186
rect 415492 6122 415544 6128
rect 415504 480 415532 6122
rect 416700 480 416728 6258
rect 420184 6248 420236 6254
rect 420184 6190 420236 6196
rect 418988 3528 419040 3534
rect 418988 3470 419040 3476
rect 417884 3460 417936 3466
rect 417884 3402 417936 3408
rect 417896 480 417924 3402
rect 419000 480 419028 3470
rect 420196 480 420224 6190
rect 430856 4140 430908 4146
rect 430856 4082 430908 4088
rect 429660 4072 429712 4078
rect 429660 4014 429712 4020
rect 428464 4004 428516 4010
rect 428464 3946 428516 3952
rect 426164 3936 426216 3942
rect 426164 3878 426216 3884
rect 424968 3800 425020 3806
rect 424968 3742 425020 3748
rect 423772 3732 423824 3738
rect 423772 3674 423824 3680
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 421380 3596 421432 3602
rect 421380 3538 421432 3544
rect 421392 480 421420 3538
rect 422588 480 422616 3606
rect 423784 480 423812 3674
rect 424980 480 425008 3742
rect 426176 480 426204 3878
rect 427268 3868 427320 3874
rect 427268 3810 427320 3816
rect 427280 480 427308 3810
rect 428476 480 428504 3946
rect 429672 480 429700 4014
rect 430868 480 430896 4082
rect 435546 3768 435602 3777
rect 435546 3703 435602 3712
rect 433246 3632 433302 3641
rect 433246 3567 433302 3576
rect 434352 3596 434404 3602
rect 432050 3360 432106 3369
rect 432050 3295 432106 3304
rect 432064 480 432092 3295
rect 433260 480 433288 3567
rect 434352 3538 434404 3544
rect 434444 3596 434496 3602
rect 434444 3538 434496 3544
rect 434364 3398 434392 3538
rect 434352 3392 434404 3398
rect 434352 3334 434404 3340
rect 434456 480 434484 3538
rect 435560 480 435588 3703
rect 436756 480 436784 253302
rect 436848 158438 436876 308790
rect 438032 308712 438084 308718
rect 438032 308654 438084 308660
rect 437480 308440 437532 308446
rect 437480 308382 437532 308388
rect 436928 248124 436980 248130
rect 436928 248066 436980 248072
rect 436836 158432 436888 158438
rect 436836 158374 436888 158380
rect 436940 158234 436968 248066
rect 436928 158228 436980 158234
rect 436928 158170 436980 158176
rect 437492 3806 437520 308382
rect 437572 247920 437624 247926
rect 437572 247862 437624 247868
rect 437584 3942 437612 247862
rect 437664 245540 437716 245546
rect 437664 245482 437716 245488
rect 437676 4146 437704 245482
rect 437848 245404 437900 245410
rect 437848 245346 437900 245352
rect 437756 245200 437808 245206
rect 437756 245142 437808 245148
rect 437664 4140 437716 4146
rect 437664 4082 437716 4088
rect 437572 3936 437624 3942
rect 437572 3878 437624 3884
rect 437480 3800 437532 3806
rect 437480 3742 437532 3748
rect 437768 3466 437796 245142
rect 437860 3738 437888 245346
rect 437940 245268 437992 245274
rect 437940 245210 437992 245216
rect 437952 16574 437980 245210
rect 438044 158574 438072 308654
rect 438032 158568 438084 158574
rect 438032 158510 438084 158516
rect 438136 158370 438164 308858
rect 439504 308780 439556 308786
rect 439504 308722 439556 308728
rect 439412 308644 439464 308650
rect 439412 308586 439464 308592
rect 438216 248192 438268 248198
rect 438216 248134 438268 248140
rect 438124 158364 438176 158370
rect 438124 158306 438176 158312
rect 438228 157894 438256 248134
rect 438860 247852 438912 247858
rect 438860 247794 438912 247800
rect 438308 244792 438360 244798
rect 438308 244734 438360 244740
rect 438320 158166 438348 244734
rect 438308 158160 438360 158166
rect 438308 158102 438360 158108
rect 438216 157888 438268 157894
rect 438216 157830 438268 157836
rect 437952 16546 438072 16574
rect 437848 3732 437900 3738
rect 437848 3674 437900 3680
rect 438044 3534 438072 16546
rect 438872 4078 438900 247794
rect 439044 245472 439096 245478
rect 439044 245414 439096 245420
rect 438952 245064 439004 245070
rect 438952 245006 439004 245012
rect 438860 4072 438912 4078
rect 438860 4014 438912 4020
rect 438964 3670 438992 245006
rect 439056 11778 439084 245414
rect 439136 245336 439188 245342
rect 439136 245278 439188 245284
rect 439148 11898 439176 245278
rect 439320 245132 439372 245138
rect 439320 245074 439372 245080
rect 439228 244996 439280 245002
rect 439228 244938 439280 244944
rect 439136 11892 439188 11898
rect 439136 11834 439188 11840
rect 439056 11750 439176 11778
rect 439044 11688 439096 11694
rect 439044 11630 439096 11636
rect 439056 4010 439084 11630
rect 439044 4004 439096 4010
rect 439044 3946 439096 3952
rect 438952 3664 439004 3670
rect 438952 3606 439004 3612
rect 439148 3602 439176 11750
rect 439136 3596 439188 3602
rect 439136 3538 439188 3544
rect 438032 3528 438084 3534
rect 437938 3496 437994 3505
rect 437756 3460 437808 3466
rect 438032 3470 438084 3476
rect 439134 3496 439190 3505
rect 437938 3431 437994 3440
rect 439134 3431 439190 3440
rect 437756 3402 437808 3408
rect 437952 480 437980 3431
rect 439148 480 439176 3431
rect 439240 3398 439268 244938
rect 439332 3874 439360 245074
rect 439424 158506 439452 308586
rect 439412 158500 439464 158506
rect 439412 158442 439464 158448
rect 439516 158302 439544 308722
rect 440424 308576 440476 308582
rect 440424 308518 440476 308524
rect 439596 308508 439648 308514
rect 439596 308450 439648 308456
rect 439608 158710 439636 308450
rect 440240 289264 440292 289270
rect 440240 289206 440292 289212
rect 439688 244724 439740 244730
rect 439688 244666 439740 244672
rect 439596 158704 439648 158710
rect 439596 158646 439648 158652
rect 439504 158296 439556 158302
rect 439504 158238 439556 158244
rect 439700 157826 439728 244666
rect 439688 157820 439740 157826
rect 439688 157762 439740 157768
rect 439320 3868 439372 3874
rect 439320 3810 439372 3816
rect 439228 3392 439280 3398
rect 439228 3334 439280 3340
rect 440252 3346 440280 289206
rect 440332 285116 440384 285122
rect 440332 285058 440384 285064
rect 440344 3534 440372 285058
rect 440436 158642 440464 308518
rect 441620 250572 441672 250578
rect 441620 250514 441672 250520
rect 440516 248056 440568 248062
rect 440516 247998 440568 248004
rect 440528 158778 440556 247998
rect 440608 245608 440660 245614
rect 440608 245550 440660 245556
rect 440516 158772 440568 158778
rect 440516 158714 440568 158720
rect 440424 158636 440476 158642
rect 440424 158578 440476 158584
rect 440620 158098 440648 245550
rect 440608 158092 440660 158098
rect 440608 158034 440660 158040
rect 441632 16574 441660 250514
rect 441712 247988 441764 247994
rect 441712 247930 441764 247936
rect 441724 158030 441752 247930
rect 441804 244860 441856 244866
rect 441804 244802 441856 244808
rect 441712 158024 441764 158030
rect 441712 157966 441764 157972
rect 441816 157962 441844 244802
rect 441804 157956 441856 157962
rect 441804 157898 441856 157904
rect 442276 113150 442304 444790
rect 458836 439550 458864 445742
rect 580264 445052 580316 445058
rect 580264 444994 580316 445000
rect 526444 444780 526496 444786
rect 526444 444722 526496 444728
rect 458824 439544 458876 439550
rect 458824 439486 458876 439492
rect 445024 307284 445076 307290
rect 445024 307226 445076 307232
rect 442354 303240 442410 303249
rect 442354 303175 442410 303184
rect 442264 113144 442316 113150
rect 442264 113086 442316 113092
rect 441632 16546 442304 16574
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442276 3482 442304 16546
rect 442368 3602 442396 303175
rect 443000 283756 443052 283762
rect 443000 283698 443052 283704
rect 443012 16574 443040 283698
rect 444380 274100 444432 274106
rect 444380 274042 444432 274048
rect 443012 16546 443408 16574
rect 442356 3596 442408 3602
rect 442356 3538 442408 3544
rect 440252 3318 440372 3346
rect 440344 480 440372 3318
rect 441540 480 441568 3470
rect 442276 3454 442672 3482
rect 442644 480 442672 3454
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 444392 6914 444420 274042
rect 445036 16574 445064 307226
rect 467104 307216 467156 307222
rect 467104 307158 467156 307164
rect 458824 304496 458876 304502
rect 458824 304438 458876 304444
rect 449900 287768 449952 287774
rect 449900 287710 449952 287716
rect 448520 286544 448572 286550
rect 448520 286486 448572 286492
rect 446404 271312 446456 271318
rect 446404 271254 446456 271260
rect 445760 260296 445812 260302
rect 445760 260238 445812 260244
rect 445036 16546 445156 16574
rect 444392 6886 445064 6914
rect 445036 480 445064 6886
rect 445128 3466 445156 16546
rect 445116 3460 445168 3466
rect 445116 3402 445168 3408
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 260238
rect 446416 3398 446444 271254
rect 447416 3596 447468 3602
rect 447416 3538 447468 3544
rect 446404 3392 446456 3398
rect 446404 3334 446456 3340
rect 447428 480 447456 3538
rect 448532 3346 448560 286486
rect 448612 246492 448664 246498
rect 448612 246434 448664 246440
rect 448624 3534 448652 246434
rect 449912 16574 449940 287710
rect 456892 286476 456944 286482
rect 456892 286418 456944 286424
rect 456800 286408 456852 286414
rect 456800 286350 456852 286356
rect 454684 283688 454736 283694
rect 454684 283630 454736 283636
rect 450544 282328 450596 282334
rect 450544 282270 450596 282276
rect 449912 16546 450492 16574
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 450464 3482 450492 16546
rect 450556 3602 450584 282270
rect 452660 280968 452712 280974
rect 452660 280910 452712 280916
rect 452672 16574 452700 280910
rect 453304 269952 453356 269958
rect 453304 269894 453356 269900
rect 452672 16546 453252 16574
rect 450544 3596 450596 3602
rect 450544 3538 450596 3544
rect 453224 3482 453252 16546
rect 453316 3602 453344 269894
rect 453304 3596 453356 3602
rect 453304 3538 453356 3544
rect 454500 3528 454552 3534
rect 448532 3318 448652 3346
rect 448624 480 448652 3318
rect 449820 480 449848 3470
rect 450464 3454 450952 3482
rect 453224 3454 453344 3482
rect 454500 3470 454552 3476
rect 450924 480 450952 3454
rect 452108 3392 452160 3398
rect 452108 3334 452160 3340
rect 452120 480 452148 3334
rect 453316 480 453344 3454
rect 454512 480 454540 3470
rect 454696 3330 454724 283630
rect 455696 3596 455748 3602
rect 455696 3538 455748 3544
rect 454684 3324 454736 3330
rect 454684 3266 454736 3272
rect 455708 480 455736 3538
rect 456812 3346 456840 286350
rect 456904 3534 456932 286418
rect 458836 3602 458864 304438
rect 462964 297628 463016 297634
rect 462964 297570 463016 297576
rect 460940 279608 460992 279614
rect 460940 279550 460992 279556
rect 460204 268524 460256 268530
rect 460204 268466 460256 268472
rect 459560 249144 459612 249150
rect 459560 249086 459612 249092
rect 459572 16574 459600 249086
rect 459572 16546 459968 16574
rect 458824 3596 458876 3602
rect 458824 3538 458876 3544
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456812 3318 456932 3346
rect 456904 480 456932 3318
rect 458100 480 458128 3470
rect 459192 3324 459244 3330
rect 459192 3266 459244 3272
rect 459204 480 459232 3266
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 460216 4146 460244 268466
rect 460952 16574 460980 279550
rect 460952 16546 461624 16574
rect 460204 4140 460256 4146
rect 460204 4082 460256 4088
rect 461596 480 461624 16546
rect 462780 4140 462832 4146
rect 462780 4082 462832 4088
rect 462792 480 462820 4082
rect 462976 3534 463004 297570
rect 463700 279540 463752 279546
rect 463700 279482 463752 279488
rect 463712 16574 463740 279482
rect 464344 267232 464396 267238
rect 464344 267174 464396 267180
rect 463712 16546 464016 16574
rect 462964 3528 463016 3534
rect 462964 3470 463016 3476
rect 463988 480 464016 16546
rect 464356 3058 464384 267174
rect 466460 258868 466512 258874
rect 466460 258810 466512 258816
rect 466472 16574 466500 258810
rect 466472 16546 467052 16574
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 3538
rect 467024 3482 467052 16546
rect 467116 3602 467144 307158
rect 476764 307148 476816 307154
rect 476764 307090 476816 307096
rect 468484 301640 468536 301646
rect 468484 301582 468536 301588
rect 467840 254652 467892 254658
rect 467840 254594 467892 254600
rect 467852 16574 467880 254594
rect 467852 16546 468248 16574
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 467024 3454 467512 3482
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 3454
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 4146 468524 301582
rect 471242 300384 471298 300393
rect 471242 300319 471298 300328
rect 468484 4140 468536 4146
rect 468484 4082 468536 4088
rect 471060 4140 471112 4146
rect 471060 4082 471112 4088
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 471072 480 471100 4082
rect 471256 3534 471284 300319
rect 473452 297560 473504 297566
rect 473452 297502 473504 297508
rect 471980 258800 472032 258806
rect 471980 258742 472032 258748
rect 471992 16574 472020 258742
rect 473464 16574 473492 297502
rect 475384 282260 475436 282266
rect 475384 282202 475436 282208
rect 474740 254584 474792 254590
rect 474740 254526 474792 254532
rect 474752 16574 474780 254526
rect 471992 16546 472296 16574
rect 473464 16546 474136 16574
rect 474752 16546 475332 16574
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 472268 480 472296 16546
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475304 3482 475332 16546
rect 475396 3602 475424 282202
rect 476776 3942 476804 307090
rect 500224 307080 500276 307086
rect 500224 307022 500276 307028
rect 489918 306096 489974 306105
rect 489918 306031 489974 306040
rect 478144 304428 478196 304434
rect 478144 304370 478196 304376
rect 477500 276752 477552 276758
rect 477500 276694 477552 276700
rect 477512 6914 477540 276694
rect 478156 16574 478184 304370
rect 485042 303104 485098 303113
rect 485042 303039 485098 303048
rect 481640 265804 481692 265810
rect 481640 265746 481692 265752
rect 478156 16546 478276 16574
rect 477512 6886 478184 6914
rect 476764 3936 476816 3942
rect 476764 3878 476816 3884
rect 475384 3596 475436 3602
rect 475384 3538 475436 3544
rect 476948 3596 477000 3602
rect 476948 3538 477000 3544
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 476960 480 476988 3538
rect 478156 480 478184 6886
rect 478248 3602 478276 16546
rect 481652 6914 481680 265746
rect 481732 264308 481784 264314
rect 481732 264250 481784 264256
rect 481744 16574 481772 264250
rect 484400 264240 484452 264246
rect 484400 264182 484452 264188
rect 484412 16574 484440 264182
rect 481744 16546 482416 16574
rect 484412 16546 484808 16574
rect 481652 6886 481772 6914
rect 480536 3936 480588 3942
rect 480536 3878 480588 3884
rect 478236 3596 478288 3602
rect 478236 3538 478288 3544
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 3878
rect 481744 480 481772 6886
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484032 3596 484084 3602
rect 484032 3538 484084 3544
rect 484044 480 484072 3538
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485056 3194 485084 303039
rect 488540 280900 488592 280906
rect 488540 280842 488592 280848
rect 485780 278112 485832 278118
rect 485780 278054 485832 278060
rect 485792 16574 485820 278054
rect 488552 16574 488580 280842
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 485044 3188 485096 3194
rect 485044 3130 485096 3136
rect 486436 480 486464 16546
rect 487620 3188 487672 3194
rect 487620 3130 487672 3136
rect 487632 480 487660 3130
rect 488828 480 488856 16546
rect 489932 3534 489960 306031
rect 494060 301572 494112 301578
rect 494060 301514 494112 301520
rect 493324 294772 493376 294778
rect 493324 294714 493376 294720
rect 491300 279472 491352 279478
rect 491300 279414 491352 279420
rect 490012 262948 490064 262954
rect 490012 262890 490064 262896
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 262890
rect 491312 16574 491340 279414
rect 492680 275392 492732 275398
rect 492680 275334 492732 275340
rect 492692 16574 492720 275334
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 493336 3398 493364 294714
rect 494072 16574 494100 301514
rect 498290 300248 498346 300257
rect 498290 300183 498346 300192
rect 495440 262880 495492 262886
rect 495440 262822 495492 262828
rect 494072 16546 494744 16574
rect 493324 3392 493376 3398
rect 493324 3334 493376 3340
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 262822
rect 496084 261588 496136 261594
rect 496084 261530 496136 261536
rect 496096 3534 496124 261530
rect 498304 6914 498332 300183
rect 499580 274032 499632 274038
rect 499580 273974 499632 273980
rect 499592 16574 499620 273974
rect 499592 16546 500172 16574
rect 498212 6886 498332 6914
rect 496084 3528 496136 3534
rect 496084 3470 496136 3476
rect 497096 3528 497148 3534
rect 497096 3470 497148 3476
rect 497108 480 497136 3470
rect 498212 480 498240 6886
rect 500144 3482 500172 16546
rect 500236 3602 500264 307022
rect 516782 305960 516838 305969
rect 516782 305895 516838 305904
rect 514024 304360 514076 304366
rect 514024 304302 514076 304308
rect 502984 298920 503036 298926
rect 502984 298862 503036 298868
rect 502340 261520 502392 261526
rect 502340 261462 502392 261468
rect 502352 6914 502380 261462
rect 502996 16574 503024 298862
rect 507860 297492 507912 297498
rect 507860 297434 507912 297440
rect 506480 278044 506532 278050
rect 506480 277986 506532 277992
rect 503720 252000 503772 252006
rect 503720 251942 503772 251948
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 500144 3454 500632 3482
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500604 480 500632 3454
rect 501800 480 501828 3538
rect 502996 480 503024 6886
rect 503088 3058 503116 16546
rect 503076 3052 503128 3058
rect 503076 2994 503128 3000
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 251942
rect 505376 3052 505428 3058
rect 505376 2994 505428 3000
rect 505388 480 505416 2994
rect 506492 480 506520 277986
rect 506572 251932 506624 251938
rect 506572 251874 506624 251880
rect 506584 16574 506612 251874
rect 507872 16574 507900 297434
rect 512000 296132 512052 296138
rect 512000 296074 512052 296080
rect 509884 276684 509936 276690
rect 509884 276626 509936 276632
rect 509240 247784 509292 247790
rect 509240 247726 509292 247732
rect 509252 16574 509280 247726
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 509896 3330 509924 276626
rect 510620 271244 510672 271250
rect 510620 271186 510672 271192
rect 510632 16574 510660 271186
rect 510632 16546 511304 16574
rect 509884 3324 509936 3330
rect 509884 3266 509936 3272
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 296074
rect 514036 3534 514064 304302
rect 516140 285048 516192 285054
rect 516140 284990 516192 284996
rect 514116 250504 514168 250510
rect 514116 250446 514168 250452
rect 514024 3528 514076 3534
rect 514024 3470 514076 3476
rect 514128 3466 514156 250446
rect 516152 16574 516180 284990
rect 516152 16546 516732 16574
rect 515956 3528 516008 3534
rect 515956 3470 516008 3476
rect 516704 3482 516732 16546
rect 516796 3874 516824 305895
rect 520922 302968 520978 302977
rect 520922 302903 520978 302912
rect 517520 272536 517572 272542
rect 517520 272478 517572 272484
rect 517532 16574 517560 272478
rect 520280 244928 520332 244934
rect 520280 244870 520332 244876
rect 517532 16546 517928 16574
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 514116 3460 514168 3466
rect 514116 3402 514168 3408
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 513564 3324 513616 3330
rect 513564 3266 513616 3272
rect 513576 480 513604 3266
rect 514772 480 514800 3402
rect 515968 480 515996 3470
rect 516704 3454 517192 3482
rect 517164 480 517192 3454
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3868 519596 3874
rect 519544 3810 519596 3816
rect 519556 480 519584 3810
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 244870
rect 520936 3466 520964 302903
rect 521660 294704 521712 294710
rect 521660 294646 521712 294652
rect 520924 3460 520976 3466
rect 520924 3402 520976 3408
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 294646
rect 522304 293412 522356 293418
rect 522304 293354 522356 293360
rect 522316 3534 522344 293354
rect 524420 269884 524472 269890
rect 524420 269826 524472 269832
rect 524432 16574 524460 269826
rect 526456 33114 526484 444722
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 575478 305824 575534 305833
rect 575478 305759 575534 305768
rect 566464 304292 566516 304298
rect 566464 304234 566516 304240
rect 545118 302832 545174 302841
rect 545118 302767 545174 302776
rect 534724 301504 534776 301510
rect 534724 301446 534776 301452
rect 529940 294636 529992 294642
rect 529940 294578 529992 294584
rect 527824 293344 527876 293350
rect 527824 293286 527876 293292
rect 526536 275324 526588 275330
rect 526536 275266 526588 275272
rect 526444 33108 526496 33114
rect 526444 33050 526496 33056
rect 524432 16546 525472 16574
rect 522304 3528 522356 3534
rect 522304 3470 522356 3476
rect 524236 3528 524288 3534
rect 524236 3470 524288 3476
rect 523040 3460 523092 3466
rect 523040 3402 523092 3408
rect 523052 480 523080 3402
rect 524248 480 524276 3470
rect 525444 480 525472 16546
rect 526548 2990 526576 275266
rect 527836 16574 527864 293286
rect 528560 247716 528612 247722
rect 528560 247658 528612 247664
rect 527836 16546 527956 16574
rect 527928 3466 527956 16546
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 526628 3392 526680 3398
rect 526628 3334 526680 3340
rect 526536 2984 526588 2990
rect 526536 2926 526588 2932
rect 526640 480 526668 3334
rect 527824 2984 527876 2990
rect 527824 2926 527876 2932
rect 527836 480 527864 2926
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 247658
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 294578
rect 531320 273964 531372 273970
rect 531320 273906 531372 273912
rect 531332 480 531360 273906
rect 531412 268456 531464 268462
rect 531412 268398 531464 268404
rect 531424 16574 531452 268398
rect 534080 246424 534132 246430
rect 534080 246366 534132 246372
rect 534092 16574 534120 246366
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3460 533764 3466
rect 533712 3402 533764 3408
rect 533724 480 533752 3402
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3194 534764 301446
rect 543738 300112 543794 300121
rect 543738 300047 543794 300056
rect 536104 291916 536156 291922
rect 536104 291858 536156 291864
rect 535460 284980 535512 284986
rect 535460 284922 535512 284928
rect 535472 6914 535500 284922
rect 536116 16574 536144 291858
rect 538864 291848 538916 291854
rect 538864 291790 538916 291796
rect 536116 16546 536236 16574
rect 535472 6886 536144 6914
rect 534724 3188 534776 3194
rect 534724 3130 534776 3136
rect 536116 480 536144 6886
rect 536208 4146 536236 16546
rect 536196 4140 536248 4146
rect 536196 4082 536248 4088
rect 538404 4140 538456 4146
rect 538404 4082 538456 4088
rect 537208 3188 537260 3194
rect 537208 3130 537260 3136
rect 537220 480 537248 3130
rect 538416 480 538444 4082
rect 538876 3534 538904 291790
rect 540244 271176 540296 271182
rect 540244 271118 540296 271124
rect 539690 244896 539746 244905
rect 539690 244831 539746 244840
rect 539704 6914 539732 244831
rect 539612 6886 539732 6914
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539612 480 539640 6886
rect 540256 2990 540284 271118
rect 543004 269816 543056 269822
rect 543004 269758 543056 269764
rect 542360 267164 542412 267170
rect 542360 267106 542412 267112
rect 542372 16574 542400 267106
rect 542372 16546 542768 16574
rect 540796 3528 540848 3534
rect 540796 3470 540848 3476
rect 540244 2984 540296 2990
rect 540244 2926 540296 2932
rect 540808 480 540836 3470
rect 541992 2984 542044 2990
rect 541992 2926 542044 2932
rect 542004 480 542032 2926
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3466 543044 269758
rect 543752 16574 543780 300047
rect 545132 16574 545160 302767
rect 549904 298852 549956 298858
rect 549904 298794 549956 298800
rect 548524 296064 548576 296070
rect 548524 296006 548576 296012
rect 547972 290556 548024 290562
rect 547972 290498 548024 290504
rect 546500 265736 546552 265742
rect 546500 265678 546552 265684
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 543004 3460 543056 3466
rect 543004 3402 543056 3408
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 265678
rect 547984 6914 548012 290498
rect 547892 6886 548012 6914
rect 547892 480 547920 6886
rect 548536 3602 548564 296006
rect 548524 3596 548576 3602
rect 548524 3538 548576 3544
rect 549916 3534 549944 298794
rect 563704 298784 563756 298790
rect 563704 298726 563756 298732
rect 561680 297424 561732 297430
rect 561680 297366 561732 297372
rect 552664 289196 552716 289202
rect 552664 289138 552716 289144
rect 552020 268388 552072 268394
rect 552020 268330 552072 268336
rect 552032 6914 552060 268330
rect 552676 16574 552704 289138
rect 557540 287700 557592 287706
rect 557540 287642 557592 287648
rect 554044 283620 554096 283626
rect 554044 283562 554096 283568
rect 553400 249076 553452 249082
rect 553400 249018 553452 249024
rect 553412 16574 553440 249018
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 550272 3596 550324 3602
rect 550272 3538 550324 3544
rect 549904 3528 549956 3534
rect 549904 3470 549956 3476
rect 549076 3460 549128 3466
rect 549076 3402 549128 3408
rect 549088 480 549116 3402
rect 550284 480 550312 3538
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 551480 480 551508 3470
rect 552676 480 552704 6886
rect 552768 3058 552796 16546
rect 552756 3052 552808 3058
rect 552756 2994 552808 3000
rect 553780 480 553808 16546
rect 554056 3398 554084 283562
rect 556160 267096 556212 267102
rect 556160 267038 556212 267044
rect 554044 3392 554096 3398
rect 554044 3334 554096 3340
rect 554964 3052 555016 3058
rect 554964 2994 555016 3000
rect 554976 480 555004 2994
rect 556172 480 556200 267038
rect 556252 246356 556304 246362
rect 556252 246298 556304 246304
rect 556264 16574 556292 246298
rect 557552 16574 557580 287642
rect 560944 265668 560996 265674
rect 560944 265610 560996 265616
rect 560300 251864 560352 251870
rect 560300 251806 560352 251812
rect 560312 16574 560340 251806
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 559748 3392 559800 3398
rect 559748 3334 559800 3340
rect 559760 480 559788 3334
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 560956 3194 560984 265610
rect 561692 16574 561720 297366
rect 561692 16546 562088 16574
rect 560944 3188 560996 3194
rect 560944 3130 560996 3136
rect 562060 480 562088 16546
rect 563716 3534 563744 298726
rect 563796 286340 563848 286346
rect 563796 286282 563848 286288
rect 563704 3528 563756 3534
rect 563704 3470 563756 3476
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 563808 3058 563836 286282
rect 564532 260160 564584 260166
rect 564532 260102 564584 260108
rect 564544 6914 564572 260102
rect 564452 6886 564572 6914
rect 563796 3052 563848 3058
rect 563796 2994 563848 3000
rect 564452 480 564480 6886
rect 566476 4146 566504 304234
rect 570604 295996 570656 296002
rect 570604 295938 570656 295944
rect 567844 290488 567896 290494
rect 567844 290430 567896 290436
rect 567200 280832 567252 280838
rect 567200 280774 567252 280780
rect 567212 16574 567240 280774
rect 567212 16546 567608 16574
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 566832 3528 566884 3534
rect 566832 3470 566884 3476
rect 565636 3052 565688 3058
rect 565636 2994 565688 3000
rect 565648 480 565676 2994
rect 566844 480 566872 3470
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3194 567884 290430
rect 569132 4140 569184 4146
rect 569132 4082 569184 4088
rect 567844 3188 567896 3194
rect 567844 3130 567896 3136
rect 569144 480 569172 4082
rect 570328 3188 570380 3194
rect 570328 3130 570380 3136
rect 570340 480 570368 3130
rect 570616 3126 570644 295938
rect 571984 289128 572036 289134
rect 571984 289070 572036 289076
rect 571340 253292 571392 253298
rect 571340 253234 571392 253240
rect 570604 3120 570656 3126
rect 570604 3062 570656 3068
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 253234
rect 571996 3330 572024 289070
rect 574744 282192 574796 282198
rect 574744 282134 574796 282140
rect 574100 253224 574152 253230
rect 574100 253166 574152 253172
rect 574112 16574 574140 253166
rect 574112 16546 574692 16574
rect 574664 3482 574692 16546
rect 574756 3874 574784 282134
rect 575492 16574 575520 305759
rect 578240 293276 578292 293282
rect 578240 293218 578292 293224
rect 578252 16574 578280 293218
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580276 152697 580304 444994
rect 581000 442264 581052 442270
rect 581000 442206 581052 442212
rect 580448 260228 580500 260234
rect 580448 260170 580500 260176
rect 580356 258732 580408 258738
rect 580356 258674 580408 258680
rect 580368 192545 580396 258674
rect 580460 232393 580488 260170
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 574744 3868 574796 3874
rect 574744 3810 574796 3816
rect 574664 3454 575152 3482
rect 571984 3324 572036 3330
rect 571984 3266 572036 3272
rect 573916 3324 573968 3330
rect 573916 3266 573968 3272
rect 572720 3120 572772 3126
rect 572720 3062 572772 3068
rect 572732 480 572760 3062
rect 573928 480 573956 3266
rect 575124 480 575152 3454
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 577424 480 577452 3810
rect 578620 480 578648 16546
rect 581012 3534 581040 442206
rect 582380 439544 582432 439550
rect 582380 439486 582432 439492
rect 581092 257372 581144 257378
rect 581092 257314 581144 257320
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581104 3346 581132 257314
rect 582392 16574 582420 439486
rect 582392 16546 583432 16574
rect 581828 3528 581880 3534
rect 581828 3470 581880 3476
rect 581012 3318 581132 3346
rect 581012 480 581040 3318
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581840 354 581868 3470
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581840 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 619112 3478 619168
rect 3330 579944 3386 580000
rect 2962 527856 3018 527912
rect 3330 501744 3386 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 2870 449520 2926 449576
rect 3514 606076 3570 606112
rect 3514 606056 3516 606076
rect 3516 606056 3568 606076
rect 3568 606056 3570 606076
rect 3514 566888 3570 566944
rect 3606 553832 3662 553888
rect 3606 514800 3662 514856
rect 217874 516840 217930 516896
rect 217782 515888 217838 515944
rect 217598 513712 217654 513768
rect 217322 488280 217378 488336
rect 217506 488008 217562 488064
rect 217690 489912 217746 489968
rect 219162 512760 219218 512816
rect 219070 508136 219126 508192
rect 219346 510992 219402 511048
rect 219254 509904 219310 509960
rect 247038 477400 247094 477456
rect 242898 476992 242954 477048
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 397432 3386 397488
rect 3054 371320 3110 371376
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3146 214920 3202 214976
rect 3146 188808 3202 188864
rect 3606 358400 3662 358456
rect 3514 201864 3570 201920
rect 3514 162832 3570 162888
rect 3422 149776 3478 149832
rect 3146 136720 3202 136776
rect 3146 110608 3202 110664
rect 3422 84632 3478 84688
rect 3698 97552 3754 97608
rect 3606 45464 3662 45520
rect 3422 6432 3478 6488
rect 40682 305632 40738 305688
rect 97814 196832 97870 196888
rect 97906 195880 97962 195936
rect 97906 193704 97962 193760
rect 97814 192752 97870 192808
rect 97722 190984 97778 191040
rect 97630 189896 97686 189952
rect 97538 188128 97594 188184
rect 97446 169904 97502 169960
rect 97354 168272 97410 168328
rect 235998 476332 236054 476368
rect 235998 476312 236000 476332
rect 236000 476312 236052 476332
rect 236052 476312 236054 476332
rect 235998 476176 236054 476232
rect 237378 476196 237434 476232
rect 237378 476176 237380 476196
rect 237380 476176 237432 476196
rect 237432 476176 237434 476196
rect 248418 476992 248474 477048
rect 244646 476856 244702 476912
rect 239126 476468 239182 476504
rect 239126 476448 239128 476468
rect 239128 476448 239180 476468
rect 239180 476448 239182 476468
rect 244278 476468 244334 476504
rect 244278 476448 244280 476468
rect 244280 476448 244332 476468
rect 244332 476448 244334 476468
rect 240230 476176 240286 476232
rect 242806 476176 242862 476232
rect 245658 476196 245714 476232
rect 245658 476176 245660 476196
rect 245660 476176 245712 476196
rect 245712 476176 245714 476196
rect 247038 476584 247094 476640
rect 249890 477400 249946 477456
rect 252466 477400 252522 477456
rect 253846 477400 253902 477456
rect 249798 476448 249854 476504
rect 252374 476196 252430 476232
rect 252374 476176 252376 476196
rect 252376 476176 252428 476196
rect 252428 476176 252430 476196
rect 252558 476604 252614 476640
rect 252558 476584 252560 476604
rect 252560 476584 252612 476604
rect 252612 476584 252614 476604
rect 268014 477264 268070 477320
rect 255410 476992 255466 477048
rect 258078 477012 258134 477048
rect 258078 476992 258080 477012
rect 258080 476992 258132 477012
rect 258132 476992 258134 477012
rect 258078 476740 258134 476776
rect 258078 476720 258080 476740
rect 258080 476720 258132 476740
rect 258132 476720 258134 476740
rect 258262 476720 258318 476776
rect 255962 476312 256018 476368
rect 256606 476176 256662 476232
rect 260838 476584 260894 476640
rect 260746 476176 260802 476232
rect 261482 476312 261538 476368
rect 263598 476584 263654 476640
rect 264978 476604 265034 476640
rect 264978 476584 264980 476604
rect 264980 476584 265032 476604
rect 265032 476584 265034 476604
rect 264242 476448 264298 476504
rect 270498 476992 270554 477048
rect 304998 476992 305054 477048
rect 307758 476992 307814 477048
rect 262862 476176 262918 476232
rect 265622 476312 265678 476368
rect 267554 476312 267610 476368
rect 302238 476856 302294 476912
rect 277950 476584 278006 476640
rect 273258 476448 273314 476504
rect 266266 476176 266322 476232
rect 274454 476312 274510 476368
rect 276018 476312 276074 476368
rect 267646 476176 267702 476232
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476176 271842 476232
rect 273166 476176 273222 476232
rect 274546 476176 274602 476232
rect 275926 476176 275982 476232
rect 277306 476176 277362 476232
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 280250 476176 280306 476232
rect 283102 476176 283158 476232
rect 285770 476176 285826 476232
rect 287058 476176 287114 476232
rect 289910 476176 289966 476232
rect 292578 476176 292634 476232
rect 295430 476176 295486 476232
rect 298190 476176 298246 476232
rect 300858 476176 300914 476232
rect 310518 476856 310574 476912
rect 313278 476468 313334 476504
rect 313278 476448 313280 476468
rect 313280 476448 313332 476468
rect 313332 476448 313334 476468
rect 314658 476448 314714 476504
rect 322938 476856 322994 476912
rect 325790 476856 325846 476912
rect 317418 476332 317474 476368
rect 317418 476312 317420 476332
rect 317420 476312 317472 476332
rect 317472 476312 317474 476332
rect 320178 476312 320234 476368
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 484608 580226 484664
rect 298006 442992 298062 443048
rect 359462 442720 359518 442776
rect 99286 168000 99342 168056
rect 160926 159840 160982 159896
rect 163502 159840 163558 159896
rect 165986 159840 166042 159896
rect 203430 159840 203486 159896
rect 200118 159296 200174 159352
rect 116858 158616 116914 158672
rect 119710 158652 119712 158672
rect 119712 158652 119764 158672
rect 119764 158652 119766 158672
rect 119710 158616 119766 158652
rect 121182 158616 121238 158672
rect 122102 158616 122158 158672
rect 123206 158616 123262 158672
rect 125322 158616 125378 158672
rect 126518 158616 126574 158672
rect 127622 158616 127678 158672
rect 128726 158616 128782 158672
rect 130198 158616 130254 158672
rect 131302 158636 131358 158672
rect 131302 158616 131304 158636
rect 131304 158616 131356 158636
rect 131356 158616 131358 158636
rect 117226 158208 117282 158264
rect 118238 157392 118294 157448
rect 125414 157936 125470 157992
rect 132406 158616 132462 158672
rect 133510 158616 133566 158672
rect 134890 158616 134946 158672
rect 158166 158616 158222 158672
rect 158534 158616 158590 158672
rect 159822 158616 159878 158672
rect 168286 158616 168342 158672
rect 191102 158616 191158 158672
rect 135902 158480 135958 158536
rect 137006 158480 137062 158536
rect 139214 158480 139270 158536
rect 140686 158480 140742 158536
rect 136086 157392 136142 157448
rect 125598 156576 125654 156632
rect 138938 157392 138994 157448
rect 140594 157936 140650 157992
rect 150254 158344 150310 158400
rect 141422 158208 141478 158264
rect 141790 158208 141846 158264
rect 146022 158208 146078 158264
rect 146390 158208 146446 158264
rect 144274 157800 144330 157856
rect 145286 157800 145342 157856
rect 143078 157528 143134 157584
rect 144366 157392 144422 157448
rect 148782 157800 148838 157856
rect 147770 157528 147826 157584
rect 148414 157392 148470 157448
rect 150990 158208 151046 158264
rect 178958 158344 179014 158400
rect 181718 158344 181774 158400
rect 151358 157392 151414 157448
rect 152646 157392 152702 157448
rect 153934 157392 153990 157448
rect 154486 157392 154542 157448
rect 155774 157392 155830 157448
rect 157062 157392 157118 157448
rect 178038 156712 178094 156768
rect 160098 155216 160154 155272
rect 185950 158072 186006 158128
rect 195886 158344 195942 158400
rect 198462 158344 198518 158400
rect 193954 157800 194010 157856
rect 185950 155896 186006 155952
rect 182178 155352 182234 155408
rect 213918 159432 213974 159488
rect 201038 157528 201094 157584
rect 206282 157528 206338 157584
rect 202878 156848 202934 156904
rect 220818 155488 220874 155544
rect 238022 308352 238078 308408
rect 238022 159024 238078 159080
rect 238206 158208 238262 158264
rect 238390 158072 238446 158128
rect 247774 308488 247830 308544
rect 247774 159160 247830 159216
rect 252834 156576 252890 156632
rect 255962 156712 256018 156768
rect 256974 306584 257030 306640
rect 257158 306312 257214 306368
rect 259918 155216 259974 155272
rect 260194 160656 260250 160712
rect 262494 155352 262550 155408
rect 265622 159296 265678 159352
rect 266818 156848 266874 156904
rect 268658 300464 268714 300520
rect 269670 159432 269726 159488
rect 269762 150320 269818 150376
rect 270958 155488 271014 155544
rect 273994 303456 274050 303512
rect 274638 158208 274694 158264
rect 273994 157256 274050 157312
rect 276018 158344 276074 158400
rect 275926 158208 275982 158264
rect 277582 307944 277638 308000
rect 277398 307808 277454 307864
rect 277306 158344 277362 158400
rect 278594 300600 278650 300656
rect 278686 157528 278742 157584
rect 280066 300736 280122 300792
rect 282366 158480 282422 158536
rect 284758 247016 284814 247072
rect 284666 158480 284722 158536
rect 284850 158480 284906 158536
rect 284574 158108 284576 158128
rect 284576 158108 284628 158128
rect 284628 158108 284630 158128
rect 284574 158072 284630 158108
rect 285402 307808 285458 307864
rect 285402 158752 285458 158808
rect 285310 158072 285366 158128
rect 285586 247152 285642 247208
rect 285586 169768 285642 169824
rect 286966 307808 287022 307864
rect 286690 247016 286746 247072
rect 286966 247016 287022 247072
rect 286966 158752 287022 158808
rect 287978 247152 288034 247208
rect 287886 247016 287942 247072
rect 288070 159024 288126 159080
rect 287978 158888 288034 158944
rect 287886 158752 287942 158808
rect 289358 247152 289414 247208
rect 289174 247016 289230 247072
rect 289358 158752 289414 158808
rect 289726 158888 289782 158944
rect 289634 157936 289690 157992
rect 290186 309032 290242 309088
rect 290462 308896 290518 308952
rect 290646 244296 290702 244352
rect 290646 158752 290702 158808
rect 291750 244296 291806 244352
rect 292118 244296 292174 244352
rect 292486 158752 292542 158808
rect 293498 309032 293554 309088
rect 293406 308896 293462 308952
rect 293406 244296 293462 244352
rect 293866 307808 293922 307864
rect 293774 244296 293830 244352
rect 293866 196016 293922 196072
rect 294878 168408 294934 168464
rect 295062 244296 295118 244352
rect 295982 307808 296038 307864
rect 297178 307808 297234 307864
rect 297546 308080 297602 308136
rect 298006 307944 298062 308000
rect 297822 307808 297878 307864
rect 298466 307808 298522 307864
rect 296810 244976 296866 245032
rect 297086 244976 297142 245032
rect 297086 244568 297142 244624
rect 297362 195880 297418 195936
rect 297362 193160 297418 193216
rect 297362 192752 297418 192808
rect 297546 193160 297602 193216
rect 297454 190984 297510 191040
rect 297546 189896 297602 189952
rect 297638 188128 297694 188184
rect 297822 244332 297824 244352
rect 297824 244332 297876 244352
rect 297876 244332 297878 244352
rect 297822 244296 297878 244332
rect 297730 168272 297786 168328
rect 298190 244840 298246 244896
rect 298926 307944 298982 308000
rect 298282 244432 298338 244488
rect 298374 244296 298430 244352
rect 298006 169904 298062 169960
rect 298006 167048 298062 167104
rect 299110 245520 299166 245576
rect 298742 244568 298798 244624
rect 298650 196832 298706 196888
rect 298834 193704 298890 193760
rect 298926 188128 298982 188184
rect 299110 158616 299166 158672
rect 299662 244976 299718 245032
rect 299938 248104 299994 248160
rect 299846 247424 299902 247480
rect 299478 244704 299534 244760
rect 301318 308216 301374 308272
rect 301962 308896 302018 308952
rect 301134 248240 301190 248296
rect 301226 247968 301282 248024
rect 302238 245248 302294 245304
rect 302514 247832 302570 247888
rect 302606 247696 302662 247752
rect 302698 247560 302754 247616
rect 301042 245112 301098 245168
rect 304998 308896 305054 308952
rect 309138 245112 309194 245168
rect 309598 275168 309654 275224
rect 310886 287680 310942 287736
rect 309414 247560 309470 247616
rect 312818 308216 312874 308272
rect 312358 303184 312414 303240
rect 313922 308216 313978 308272
rect 314106 307944 314162 308000
rect 316682 308216 316738 308272
rect 316314 300328 316370 300384
rect 318062 307944 318118 308000
rect 319442 308216 319498 308272
rect 319166 303048 319222 303104
rect 320730 306040 320786 306096
rect 320546 300192 320602 300248
rect 309322 244976 309378 245032
rect 325330 305904 325386 305960
rect 326066 302912 326122 302968
rect 331126 305768 331182 305824
rect 330298 302776 330354 302832
rect 330206 300056 330262 300112
rect 332230 305768 332286 305824
rect 328458 244840 328514 244896
rect 336094 305768 336150 305824
rect 337750 308352 337806 308408
rect 338854 306312 338910 306368
rect 340050 303456 340106 303512
rect 300950 244296 301006 244352
rect 345294 300464 345350 300520
rect 346858 308488 346914 308544
rect 347502 308760 347558 308816
rect 350722 300736 350778 300792
rect 352102 308624 352158 308680
rect 354862 303320 354918 303376
rect 354770 300600 354826 300656
rect 355414 306176 355470 306232
rect 360934 305632 360990 305688
rect 299386 168000 299442 168056
rect 299386 167048 299442 167104
rect 345938 159840 345994 159896
rect 348238 159840 348294 159896
rect 353574 159840 353630 159896
rect 365902 159840 365958 159896
rect 299570 158616 299626 158672
rect 300858 151000 300914 151056
rect 309138 153720 309194 153776
rect 316038 158616 316094 158672
rect 316682 158616 316738 158672
rect 319442 158616 319498 158672
rect 317694 157392 317750 157448
rect 350998 159704 351054 159760
rect 356058 159568 356114 159624
rect 358450 159568 358506 159624
rect 373998 159296 374054 159352
rect 320546 158616 320602 158672
rect 323122 158616 323178 158672
rect 324226 158616 324282 158672
rect 326434 158616 326490 158672
rect 328274 158636 328330 158672
rect 328274 158616 328276 158636
rect 328276 158616 328328 158636
rect 328328 158616 328330 158636
rect 325146 157936 325202 157992
rect 328642 158616 328698 158672
rect 329930 158616 329986 158672
rect 330482 158616 330538 158672
rect 332230 158616 332286 158672
rect 333610 158616 333666 158672
rect 334530 158616 334586 158672
rect 335634 158616 335690 158672
rect 336002 158616 336058 158672
rect 336830 158616 336886 158672
rect 338394 158652 338396 158672
rect 338396 158652 338448 158672
rect 338448 158652 338450 158672
rect 338394 158616 338450 158652
rect 338762 158616 338818 158672
rect 340970 158616 341026 158672
rect 343546 158616 343602 158672
rect 349802 158616 349858 158672
rect 355230 158616 355286 158672
rect 356978 158616 357034 158672
rect 360842 158616 360898 158672
rect 363418 158616 363474 158672
rect 368202 158616 368258 158672
rect 371054 158652 371056 158672
rect 371056 158652 371108 158672
rect 371108 158652 371110 158672
rect 371054 158616 371110 158652
rect 373446 158636 373502 158672
rect 373446 158616 373448 158636
rect 373448 158616 373500 158636
rect 373500 158616 373502 158636
rect 338118 158344 338174 158400
rect 343914 158208 343970 158264
rect 348698 158208 348754 158264
rect 339498 157800 339554 157856
rect 341154 157800 341210 157856
rect 342810 157800 342866 157856
rect 346398 157936 346454 157992
rect 345110 157800 345166 157856
rect 346858 157800 346914 157856
rect 353298 158208 353354 158264
rect 351090 157392 351146 157448
rect 352194 157392 352250 157448
rect 354402 157392 354458 157448
rect 372894 6840 372950 6896
rect 369398 6024 369454 6080
rect 368202 4936 368258 4992
rect 363510 3168 363566 3224
rect 370594 4800 370650 4856
rect 376022 158616 376078 158672
rect 378598 158616 378654 158672
rect 380990 158616 381046 158672
rect 383566 158616 383622 158672
rect 385958 158616 386014 158672
rect 388534 158616 388590 158672
rect 391478 158616 391534 158672
rect 393502 158616 393558 158672
rect 395894 158616 395950 158672
rect 398470 158616 398526 158672
rect 401414 158616 401470 158672
rect 403806 158616 403862 158672
rect 406750 158616 406806 158672
rect 375378 75112 375434 75168
rect 374090 9560 374146 9616
rect 387154 9424 387210 9480
rect 379978 8744 380034 8800
rect 382370 6704 382426 6760
rect 381174 3984 381230 4040
rect 383566 3848 383622 3904
rect 394238 9288 394294 9344
rect 389454 6568 389510 6624
rect 388258 3712 388314 3768
rect 393042 6432 393098 6488
rect 390650 6296 390706 6352
rect 391846 3576 391902 3632
rect 408406 9152 408462 9208
rect 397734 9016 397790 9072
rect 396538 6160 396594 6216
rect 395342 3440 395398 3496
rect 404818 8880 404874 8936
rect 398930 3304 398986 3360
rect 435546 3712 435602 3768
rect 433246 3576 433302 3632
rect 432050 3304 432106 3360
rect 437938 3440 437994 3496
rect 439134 3440 439190 3496
rect 442354 303184 442410 303240
rect 471242 300328 471298 300384
rect 489918 306040 489974 306096
rect 485042 303048 485098 303104
rect 498290 300192 498346 300248
rect 516782 305904 516838 305960
rect 520922 302912 520978 302968
rect 580170 431568 580226 431624
rect 580170 378392 580226 378448
rect 579894 325216 579950 325272
rect 575478 305768 575534 305824
rect 545118 302776 545174 302832
rect 543738 300056 543794 300112
rect 539690 244840 539746 244896
rect 579894 272176 579950 272232
rect 580446 232328 580502 232384
rect 580354 192480 580410 192536
rect 580262 152632 580318 152688
rect 579802 112784 579858 112840
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3601 553890 3667 553893
rect -960 553888 3667 553890
rect -960 553832 3606 553888
rect 3662 553832 3667 553888
rect -960 553830 3667 553832
rect -960 553740 480 553830
rect 3601 553827 3667 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 583520 524364 584960 524604
rect 217869 516898 217935 516901
rect 219390 516898 220064 516924
rect 217869 516896 220064 516898
rect 217869 516840 217874 516896
rect 217930 516864 220064 516896
rect 217930 516840 219450 516864
rect 217869 516838 219450 516840
rect 217869 516835 217935 516838
rect 217777 515946 217843 515949
rect 219390 515946 220064 515972
rect 217777 515944 220064 515946
rect 217777 515888 217782 515944
rect 217838 515912 220064 515944
rect 217838 515888 219450 515912
rect 217777 515886 219450 515888
rect 217777 515883 217843 515886
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 217593 513770 217659 513773
rect 219390 513770 220064 513796
rect 217593 513768 220064 513770
rect 217593 513712 217598 513768
rect 217654 513736 220064 513768
rect 217654 513712 219450 513736
rect 217593 513710 219450 513712
rect 217593 513707 217659 513710
rect 219157 512818 219223 512821
rect 219390 512818 220064 512844
rect 219157 512816 220064 512818
rect 219157 512760 219162 512816
rect 219218 512784 220064 512816
rect 219218 512760 219450 512784
rect 219157 512758 219450 512760
rect 219157 512755 219223 512758
rect 583520 511172 584960 511412
rect 219390 511053 220064 511076
rect 219341 511048 220064 511053
rect 219341 510992 219346 511048
rect 219402 511016 220064 511048
rect 219402 510992 219450 511016
rect 219341 510990 219450 510992
rect 219341 510987 219407 510990
rect 219249 509962 219315 509965
rect 219390 509962 220064 509988
rect 219249 509960 220064 509962
rect 219249 509904 219254 509960
rect 219310 509928 220064 509960
rect 219310 509904 219450 509928
rect 219249 509902 219450 509904
rect 219249 509899 219315 509902
rect 219065 508194 219131 508197
rect 219390 508194 220064 508220
rect 219065 508192 220064 508194
rect 219065 508136 219070 508192
rect 219126 508160 220064 508192
rect 219126 508136 219450 508160
rect 219065 508134 219450 508136
rect 219065 508131 219131 508134
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect 217685 489970 217751 489973
rect 219390 489970 220064 489996
rect 217685 489968 220064 489970
rect 217685 489912 217690 489968
rect 217746 489936 220064 489968
rect 217746 489912 219450 489936
rect 217685 489910 219450 489912
rect 217685 489907 217751 489910
rect -960 488596 480 488836
rect 217317 488338 217383 488341
rect 219390 488338 220064 488364
rect 217317 488336 220064 488338
rect 217317 488280 217322 488336
rect 217378 488304 220064 488336
rect 217378 488280 219450 488304
rect 217317 488278 219450 488280
rect 217317 488275 217383 488278
rect 217501 488066 217567 488069
rect 219390 488066 220064 488092
rect 217501 488064 220064 488066
rect 217501 488008 217506 488064
rect 217562 488032 220064 488064
rect 217562 488008 219450 488032
rect 217501 488006 219450 488008
rect 217501 488003 217567 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 247033 477458 247099 477461
rect 247534 477458 247540 477460
rect 247033 477456 247540 477458
rect 247033 477400 247038 477456
rect 247094 477400 247540 477456
rect 247033 477398 247540 477400
rect 247033 477395 247099 477398
rect 247534 477396 247540 477398
rect 247604 477396 247610 477460
rect 249885 477458 249951 477461
rect 250110 477458 250116 477460
rect 249885 477456 250116 477458
rect 249885 477400 249890 477456
rect 249946 477400 250116 477456
rect 249885 477398 250116 477400
rect 249885 477395 249951 477398
rect 250110 477396 250116 477398
rect 250180 477396 250186 477460
rect 251398 477396 251404 477460
rect 251468 477458 251474 477460
rect 252461 477458 252527 477461
rect 251468 477456 252527 477458
rect 251468 477400 252466 477456
rect 252522 477400 252527 477456
rect 251468 477398 252527 477400
rect 251468 477396 251474 477398
rect 252461 477395 252527 477398
rect 253422 477396 253428 477460
rect 253492 477458 253498 477460
rect 253841 477458 253907 477461
rect 253492 477456 253907 477458
rect 253492 477400 253846 477456
rect 253902 477400 253907 477456
rect 253492 477398 253907 477400
rect 253492 477396 253498 477398
rect 253841 477395 253907 477398
rect 268009 477322 268075 477325
rect 268326 477322 268332 477324
rect 268009 477320 268332 477322
rect 268009 477264 268014 477320
rect 268070 477264 268332 477320
rect 268009 477262 268332 477264
rect 268009 477259 268075 477262
rect 268326 477260 268332 477262
rect 268396 477260 268402 477324
rect 242893 477050 242959 477053
rect 243118 477050 243124 477052
rect 242893 477048 243124 477050
rect 242893 476992 242898 477048
rect 242954 476992 243124 477048
rect 242893 476990 243124 476992
rect 242893 476987 242959 476990
rect 243118 476988 243124 476990
rect 243188 476988 243194 477052
rect 248413 477050 248479 477053
rect 248638 477050 248644 477052
rect 248413 477048 248644 477050
rect 248413 476992 248418 477048
rect 248474 476992 248644 477048
rect 248413 476990 248644 476992
rect 248413 476987 248479 476990
rect 248638 476988 248644 476990
rect 248708 476988 248714 477052
rect 255405 477050 255471 477053
rect 258073 477052 258139 477053
rect 256182 477050 256188 477052
rect 255405 477048 256188 477050
rect 255405 476992 255410 477048
rect 255466 476992 256188 477048
rect 255405 476990 256188 476992
rect 255405 476987 255471 476990
rect 256182 476988 256188 476990
rect 256252 476988 256258 477052
rect 258022 476988 258028 477052
rect 258092 477050 258139 477052
rect 270493 477050 270559 477053
rect 270902 477050 270908 477052
rect 258092 477048 258184 477050
rect 258134 476992 258184 477048
rect 258092 476990 258184 476992
rect 270493 477048 270908 477050
rect 270493 476992 270498 477048
rect 270554 476992 270908 477048
rect 270493 476990 270908 476992
rect 258092 476988 258139 476990
rect 258073 476987 258139 476988
rect 270493 476987 270559 476990
rect 270902 476988 270908 476990
rect 270972 476988 270978 477052
rect 304993 477050 305059 477053
rect 305862 477050 305868 477052
rect 304993 477048 305868 477050
rect 304993 476992 304998 477048
rect 305054 476992 305868 477048
rect 304993 476990 305868 476992
rect 304993 476987 305059 476990
rect 305862 476988 305868 476990
rect 305932 476988 305938 477052
rect 307753 477050 307819 477053
rect 308438 477050 308444 477052
rect 307753 477048 308444 477050
rect 307753 476992 307758 477048
rect 307814 476992 308444 477048
rect 307753 476990 308444 476992
rect 307753 476987 307819 476990
rect 308438 476988 308444 476990
rect 308508 476988 308514 477052
rect 244641 476914 244707 476917
rect 245326 476914 245332 476916
rect 244641 476912 245332 476914
rect 244641 476856 244646 476912
rect 244702 476856 245332 476912
rect 244641 476854 245332 476856
rect 244641 476851 244707 476854
rect 245326 476852 245332 476854
rect 245396 476852 245402 476916
rect 302233 476914 302299 476917
rect 303470 476914 303476 476916
rect 302233 476912 303476 476914
rect 302233 476856 302238 476912
rect 302294 476856 303476 476912
rect 302233 476854 303476 476856
rect 302233 476851 302299 476854
rect 303470 476852 303476 476854
rect 303540 476852 303546 476916
rect 310513 476914 310579 476917
rect 311014 476914 311020 476916
rect 310513 476912 311020 476914
rect 310513 476856 310518 476912
rect 310574 476856 311020 476912
rect 310513 476854 311020 476856
rect 310513 476851 310579 476854
rect 311014 476852 311020 476854
rect 311084 476852 311090 476916
rect 322933 476914 322999 476917
rect 323342 476914 323348 476916
rect 322933 476912 323348 476914
rect 322933 476856 322938 476912
rect 322994 476856 323348 476912
rect 322933 476854 323348 476856
rect 322933 476851 322999 476854
rect 323342 476852 323348 476854
rect 323412 476852 323418 476916
rect 325785 476914 325851 476917
rect 325918 476914 325924 476916
rect 325785 476912 325924 476914
rect 325785 476856 325790 476912
rect 325846 476856 325924 476912
rect 325785 476854 325924 476856
rect 325785 476851 325851 476854
rect 325918 476852 325924 476854
rect 325988 476852 325994 476916
rect 257102 476716 257108 476780
rect 257172 476778 257178 476780
rect 258073 476778 258139 476781
rect 257172 476776 258139 476778
rect 257172 476720 258078 476776
rect 258134 476720 258139 476776
rect 257172 476718 258139 476720
rect 257172 476716 257178 476718
rect 258073 476715 258139 476718
rect 258257 476778 258323 476781
rect 258390 476778 258396 476780
rect 258257 476776 258396 476778
rect 258257 476720 258262 476776
rect 258318 476720 258396 476776
rect 258257 476718 258396 476720
rect 258257 476715 258323 476718
rect 258390 476716 258396 476718
rect 258460 476716 258466 476780
rect 247033 476642 247099 476645
rect 248270 476642 248276 476644
rect 247033 476640 248276 476642
rect 247033 476584 247038 476640
rect 247094 476584 248276 476640
rect 247033 476582 248276 476584
rect 247033 476579 247099 476582
rect 248270 476580 248276 476582
rect 248340 476580 248346 476644
rect 252553 476642 252619 476645
rect 253606 476642 253612 476644
rect 252553 476640 253612 476642
rect 252553 476584 252558 476640
rect 252614 476584 253612 476640
rect 252553 476582 253612 476584
rect 252553 476579 252619 476582
rect 253606 476580 253612 476582
rect 253676 476580 253682 476644
rect 260833 476642 260899 476645
rect 263593 476644 263659 476645
rect 260966 476642 260972 476644
rect 260833 476640 260972 476642
rect 260833 476584 260838 476640
rect 260894 476584 260972 476640
rect 260833 476582 260972 476584
rect 260833 476579 260899 476582
rect 260966 476580 260972 476582
rect 261036 476580 261042 476644
rect 263542 476580 263548 476644
rect 263612 476642 263659 476644
rect 264973 476642 265039 476645
rect 265934 476642 265940 476644
rect 263612 476640 263704 476642
rect 263654 476584 263704 476640
rect 263612 476582 263704 476584
rect 264973 476640 265940 476642
rect 264973 476584 264978 476640
rect 265034 476584 265940 476640
rect 264973 476582 265940 476584
rect 263612 476580 263659 476582
rect 263593 476579 263659 476580
rect 264973 476579 265039 476582
rect 265934 476580 265940 476582
rect 266004 476580 266010 476644
rect 277945 476642 278011 476645
rect 278446 476642 278452 476644
rect 277945 476640 278452 476642
rect 277945 476584 277950 476640
rect 278006 476584 278452 476640
rect 277945 476582 278452 476584
rect 277945 476579 278011 476582
rect 278446 476580 278452 476582
rect 278516 476580 278522 476644
rect 239121 476506 239187 476509
rect 239622 476506 239628 476508
rect 239121 476504 239628 476506
rect 239121 476448 239126 476504
rect 239182 476448 239628 476504
rect 239121 476446 239628 476448
rect 239121 476443 239187 476446
rect 239622 476444 239628 476446
rect 239692 476444 239698 476508
rect 244273 476506 244339 476509
rect 244406 476506 244412 476508
rect 244273 476504 244412 476506
rect 244273 476448 244278 476504
rect 244334 476448 244412 476504
rect 244273 476446 244412 476448
rect 244273 476443 244339 476446
rect 244406 476444 244412 476446
rect 244476 476444 244482 476508
rect 249793 476506 249859 476509
rect 250662 476506 250668 476508
rect 249793 476504 250668 476506
rect 249793 476448 249798 476504
rect 249854 476448 250668 476504
rect 249793 476446 250668 476448
rect 249793 476443 249859 476446
rect 250662 476444 250668 476446
rect 250732 476444 250738 476508
rect 262806 476444 262812 476508
rect 262876 476506 262882 476508
rect 264237 476506 264303 476509
rect 262876 476504 264303 476506
rect 262876 476448 264242 476504
rect 264298 476448 264303 476504
rect 262876 476446 264303 476448
rect 262876 476444 262882 476446
rect 264237 476443 264303 476446
rect 273253 476506 273319 476509
rect 273478 476506 273484 476508
rect 273253 476504 273484 476506
rect 273253 476448 273258 476504
rect 273314 476448 273484 476504
rect 273253 476446 273484 476448
rect 273253 476443 273319 476446
rect 273478 476444 273484 476446
rect 273548 476444 273554 476508
rect 313273 476506 313339 476509
rect 313406 476506 313412 476508
rect 313273 476504 313412 476506
rect 313273 476448 313278 476504
rect 313334 476448 313412 476504
rect 313273 476446 313412 476448
rect 313273 476443 313339 476446
rect 313406 476444 313412 476446
rect 313476 476444 313482 476508
rect 314653 476506 314719 476509
rect 315798 476506 315804 476508
rect 314653 476504 315804 476506
rect 314653 476448 314658 476504
rect 314714 476448 315804 476504
rect 314653 476446 315804 476448
rect 314653 476443 314719 476446
rect 315798 476444 315804 476446
rect 315868 476444 315874 476508
rect 235993 476372 236059 476373
rect 235942 476308 235948 476372
rect 236012 476370 236059 476372
rect 236012 476368 236104 476370
rect 236054 476312 236104 476368
rect 236012 476310 236104 476312
rect 236012 476308 236059 476310
rect 254526 476308 254532 476372
rect 254596 476370 254602 476372
rect 255957 476370 256023 476373
rect 254596 476368 256023 476370
rect 254596 476312 255962 476368
rect 256018 476312 256023 476368
rect 254596 476310 256023 476312
rect 254596 476308 254602 476310
rect 235993 476307 236059 476308
rect 255957 476307 256023 476310
rect 260782 476308 260788 476372
rect 260852 476370 260858 476372
rect 261477 476370 261543 476373
rect 260852 476368 261543 476370
rect 260852 476312 261482 476368
rect 261538 476312 261543 476368
rect 260852 476310 261543 476312
rect 260852 476308 260858 476310
rect 261477 476307 261543 476310
rect 263910 476308 263916 476372
rect 263980 476370 263986 476372
rect 265617 476370 265683 476373
rect 267549 476372 267615 476373
rect 267549 476370 267596 476372
rect 263980 476368 265683 476370
rect 263980 476312 265622 476368
rect 265678 476312 265683 476368
rect 263980 476310 265683 476312
rect 267504 476368 267596 476370
rect 267504 476312 267554 476368
rect 267504 476310 267596 476312
rect 263980 476308 263986 476310
rect 265617 476307 265683 476310
rect 267549 476308 267596 476310
rect 267660 476308 267666 476372
rect 273294 476308 273300 476372
rect 273364 476370 273370 476372
rect 274449 476370 274515 476373
rect 276013 476372 276079 476373
rect 276013 476370 276060 476372
rect 273364 476368 274515 476370
rect 273364 476312 274454 476368
rect 274510 476312 274515 476368
rect 273364 476310 274515 476312
rect 275968 476368 276060 476370
rect 275968 476312 276018 476368
rect 275968 476310 276060 476312
rect 273364 476308 273370 476310
rect 267549 476307 267615 476308
rect 274449 476307 274515 476310
rect 276013 476308 276060 476310
rect 276124 476308 276130 476372
rect 317413 476370 317479 476373
rect 318374 476370 318380 476372
rect 317413 476368 318380 476370
rect 317413 476312 317418 476368
rect 317474 476312 318380 476368
rect 317413 476310 318380 476312
rect 276013 476307 276079 476308
rect 317413 476307 317479 476310
rect 318374 476308 318380 476310
rect 318444 476308 318450 476372
rect 320173 476370 320239 476373
rect 320950 476370 320956 476372
rect 320173 476368 320956 476370
rect 320173 476312 320178 476368
rect 320234 476312 320956 476368
rect 320173 476310 320956 476312
rect 320173 476307 320239 476310
rect 320950 476308 320956 476310
rect 321020 476308 321026 476372
rect 235993 476234 236059 476237
rect 237046 476234 237052 476236
rect 235993 476232 237052 476234
rect 235993 476176 235998 476232
rect 236054 476176 237052 476232
rect 235993 476174 237052 476176
rect 235993 476171 236059 476174
rect 237046 476172 237052 476174
rect 237116 476172 237122 476236
rect 237373 476234 237439 476237
rect 238150 476234 238156 476236
rect 237373 476232 238156 476234
rect 237373 476176 237378 476232
rect 237434 476176 238156 476232
rect 237373 476174 238156 476176
rect 237373 476171 237439 476174
rect 238150 476172 238156 476174
rect 238220 476172 238226 476236
rect 240225 476234 240291 476237
rect 240542 476234 240548 476236
rect 240225 476232 240548 476234
rect 240225 476176 240230 476232
rect 240286 476176 240548 476232
rect 240225 476174 240548 476176
rect 240225 476171 240291 476174
rect 240542 476172 240548 476174
rect 240612 476172 240618 476236
rect 241830 476172 241836 476236
rect 241900 476234 241906 476236
rect 242801 476234 242867 476237
rect 241900 476232 242867 476234
rect 241900 476176 242806 476232
rect 242862 476176 242867 476232
rect 241900 476174 242867 476176
rect 241900 476172 241906 476174
rect 242801 476171 242867 476174
rect 245653 476234 245719 476237
rect 252369 476236 252435 476237
rect 246430 476234 246436 476236
rect 245653 476232 246436 476234
rect 245653 476176 245658 476232
rect 245714 476176 246436 476232
rect 245653 476174 246436 476176
rect 245653 476171 245719 476174
rect 246430 476172 246436 476174
rect 246500 476172 246506 476236
rect 252318 476172 252324 476236
rect 252388 476234 252435 476236
rect 252388 476232 252480 476234
rect 252430 476176 252480 476232
rect 252388 476174 252480 476176
rect 252388 476172 252435 476174
rect 255814 476172 255820 476236
rect 255884 476234 255890 476236
rect 256601 476234 256667 476237
rect 255884 476232 256667 476234
rect 255884 476176 256606 476232
rect 256662 476176 256667 476232
rect 255884 476174 256667 476176
rect 255884 476172 255890 476174
rect 252369 476171 252435 476172
rect 256601 476171 256667 476174
rect 259494 476172 259500 476236
rect 259564 476234 259570 476236
rect 260741 476234 260807 476237
rect 259564 476232 260807 476234
rect 259564 476176 260746 476232
rect 260802 476176 260807 476232
rect 259564 476174 260807 476176
rect 259564 476172 259570 476174
rect 260741 476171 260807 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262857 476234 262923 476237
rect 261772 476232 262923 476234
rect 261772 476176 262862 476232
rect 262918 476176 262923 476232
rect 261772 476174 262923 476176
rect 261772 476172 261778 476174
rect 262857 476171 262923 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266261 476234 266327 476237
rect 265452 476232 266327 476234
rect 265452 476176 266266 476232
rect 266322 476176 266327 476232
rect 265452 476174 266327 476176
rect 265452 476172 265458 476174
rect 266261 476171 266327 476174
rect 266486 476172 266492 476236
rect 266556 476234 266562 476236
rect 267641 476234 267707 476237
rect 266556 476232 267707 476234
rect 266556 476176 267646 476232
rect 267702 476176 267707 476232
rect 266556 476174 267707 476176
rect 266556 476172 266562 476174
rect 267641 476171 267707 476174
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271781 476234 271847 476237
rect 271340 476232 271847 476234
rect 271340 476176 271786 476232
rect 271842 476176 271847 476232
rect 271340 476174 271847 476176
rect 271340 476172 271346 476174
rect 271781 476171 271847 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 274398 476172 274404 476236
rect 274468 476234 274474 476236
rect 274541 476234 274607 476237
rect 275921 476236 275987 476237
rect 274468 476232 274607 476234
rect 274468 476176 274546 476232
rect 274602 476176 274607 476232
rect 274468 476174 274607 476176
rect 274468 476172 274474 476174
rect 274541 476171 274607 476174
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277301 476234 277367 476237
rect 277044 476232 277367 476234
rect 277044 476176 277306 476232
rect 277362 476176 277367 476232
rect 277044 476174 277367 476176
rect 277044 476172 277050 476174
rect 275921 476171 275987 476172
rect 277301 476171 277367 476174
rect 278078 476172 278084 476236
rect 278148 476234 278154 476236
rect 278681 476234 278747 476237
rect 278148 476232 278747 476234
rect 278148 476176 278686 476232
rect 278742 476176 278747 476232
rect 278148 476174 278747 476176
rect 278148 476172 278154 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 280245 476234 280311 476237
rect 280838 476234 280844 476236
rect 280245 476232 280844 476234
rect 280245 476176 280250 476232
rect 280306 476176 280844 476232
rect 280245 476174 280844 476176
rect 280245 476171 280311 476174
rect 280838 476172 280844 476174
rect 280908 476172 280914 476236
rect 283097 476234 283163 476237
rect 283414 476234 283420 476236
rect 283097 476232 283420 476234
rect 283097 476176 283102 476232
rect 283158 476176 283420 476232
rect 283097 476174 283420 476176
rect 283097 476171 283163 476174
rect 283414 476172 283420 476174
rect 283484 476172 283490 476236
rect 285765 476234 285831 476237
rect 285990 476234 285996 476236
rect 285765 476232 285996 476234
rect 285765 476176 285770 476232
rect 285826 476176 285996 476232
rect 285765 476174 285996 476176
rect 285765 476171 285831 476174
rect 285990 476172 285996 476174
rect 286060 476172 286066 476236
rect 287053 476234 287119 476237
rect 288198 476234 288204 476236
rect 287053 476232 288204 476234
rect 287053 476176 287058 476232
rect 287114 476176 288204 476232
rect 287053 476174 288204 476176
rect 287053 476171 287119 476174
rect 288198 476172 288204 476174
rect 288268 476172 288274 476236
rect 289905 476234 289971 476237
rect 290958 476234 290964 476236
rect 289905 476232 290964 476234
rect 289905 476176 289910 476232
rect 289966 476176 290964 476232
rect 289905 476174 290964 476176
rect 289905 476171 289971 476174
rect 290958 476172 290964 476174
rect 291028 476172 291034 476236
rect 292573 476234 292639 476237
rect 293350 476234 293356 476236
rect 292573 476232 293356 476234
rect 292573 476176 292578 476232
rect 292634 476176 293356 476232
rect 292573 476174 293356 476176
rect 292573 476171 292639 476174
rect 293350 476172 293356 476174
rect 293420 476172 293426 476236
rect 295425 476234 295491 476237
rect 295926 476234 295932 476236
rect 295425 476232 295932 476234
rect 295425 476176 295430 476232
rect 295486 476176 295932 476232
rect 295425 476174 295932 476176
rect 295425 476171 295491 476174
rect 295926 476172 295932 476174
rect 295996 476172 296002 476236
rect 298185 476234 298251 476237
rect 300853 476236 300919 476237
rect 298502 476234 298508 476236
rect 298185 476232 298508 476234
rect 298185 476176 298190 476232
rect 298246 476176 298508 476232
rect 298185 476174 298508 476176
rect 298185 476171 298251 476174
rect 298502 476172 298508 476174
rect 298572 476172 298578 476236
rect 300853 476234 300900 476236
rect 300808 476232 300900 476234
rect 300808 476176 300858 476232
rect 300808 476174 300900 476176
rect 300853 476172 300900 476174
rect 300964 476172 300970 476236
rect 300853 476171 300919 476172
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 583520 471324 584960 471564
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 2865 449578 2931 449581
rect -960 449576 2931 449578
rect -960 449520 2870 449576
rect 2926 449520 2931 449576
rect -960 449518 2931 449520
rect -960 449428 480 449518
rect 2865 449515 2931 449518
rect 583520 444668 584960 444908
rect 298001 443050 298067 443053
rect 439446 443050 439452 443052
rect 298001 443048 439452 443050
rect 298001 442992 298006 443048
rect 298062 442992 439452 443048
rect 298001 442990 439452 442992
rect 298001 442987 298067 442990
rect 439446 442988 439452 442990
rect 439516 442988 439522 443052
rect 358854 442716 358860 442780
rect 358924 442778 358930 442780
rect 359457 442778 359523 442781
rect 358924 442776 359523 442778
rect 358924 442720 359462 442776
rect 359518 442720 359523 442776
rect 358924 442718 359523 442720
rect 358924 442716 358930 442718
rect 359457 442715 359523 442718
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 583520 311932 584960 312172
rect 290181 309090 290247 309093
rect 293493 309090 293559 309093
rect 290181 309088 293559 309090
rect 290181 309032 290186 309088
rect 290242 309032 293498 309088
rect 293554 309032 293559 309088
rect 290181 309030 293559 309032
rect 290181 309027 290247 309030
rect 293493 309027 293559 309030
rect 295190 309028 295196 309092
rect 295260 309090 295266 309092
rect 295260 309030 302250 309090
rect 295260 309028 295266 309030
rect 290457 308954 290523 308957
rect 293401 308954 293467 308957
rect 290457 308952 293467 308954
rect 290457 308896 290462 308952
rect 290518 308896 293406 308952
rect 293462 308896 293467 308952
rect 290457 308894 293467 308896
rect 290457 308891 290523 308894
rect 293401 308891 293467 308894
rect 296294 308892 296300 308956
rect 296364 308954 296370 308956
rect 301957 308954 302023 308957
rect 296364 308952 302023 308954
rect 296364 308896 301962 308952
rect 302018 308896 302023 308952
rect 296364 308894 302023 308896
rect 302190 308954 302250 309030
rect 304993 308954 305059 308957
rect 302190 308952 305059 308954
rect 302190 308896 304998 308952
rect 305054 308896 305059 308952
rect 302190 308894 305059 308896
rect 296364 308892 296370 308894
rect 301957 308891 302023 308894
rect 304993 308891 305059 308894
rect 282126 308756 282132 308820
rect 282196 308818 282202 308820
rect 347497 308818 347563 308821
rect 282196 308816 347563 308818
rect 282196 308760 347502 308816
rect 347558 308760 347563 308816
rect 282196 308758 347563 308760
rect 282196 308756 282202 308758
rect 347497 308755 347563 308758
rect 286174 308620 286180 308684
rect 286244 308682 286250 308684
rect 352097 308682 352163 308685
rect 286244 308680 352163 308682
rect 286244 308624 352102 308680
rect 352158 308624 352163 308680
rect 286244 308622 352163 308624
rect 286244 308620 286250 308622
rect 352097 308619 352163 308622
rect 247769 308546 247835 308549
rect 346853 308546 346919 308549
rect 247769 308544 346919 308546
rect 247769 308488 247774 308544
rect 247830 308488 346858 308544
rect 346914 308488 346919 308544
rect 247769 308486 346919 308488
rect 247769 308483 247835 308486
rect 346853 308483 346919 308486
rect 238017 308410 238083 308413
rect 337745 308410 337811 308413
rect 238017 308408 337811 308410
rect 238017 308352 238022 308408
rect 238078 308352 337750 308408
rect 337806 308352 337811 308408
rect 238017 308350 337811 308352
rect 238017 308347 238083 308350
rect 337745 308347 337811 308350
rect 296478 308212 296484 308276
rect 296548 308274 296554 308276
rect 301313 308274 301379 308277
rect 296548 308272 301379 308274
rect 296548 308216 301318 308272
rect 301374 308216 301379 308272
rect 296548 308214 301379 308216
rect 296548 308212 296554 308214
rect 301313 308211 301379 308214
rect 312813 308274 312879 308277
rect 313917 308274 313983 308277
rect 312813 308272 313983 308274
rect 312813 308216 312818 308272
rect 312874 308216 313922 308272
rect 313978 308216 313983 308272
rect 312813 308214 313983 308216
rect 312813 308211 312879 308214
rect 313917 308211 313983 308214
rect 316677 308274 316743 308277
rect 319437 308274 319503 308277
rect 316677 308272 319503 308274
rect 316677 308216 316682 308272
rect 316738 308216 319442 308272
rect 319498 308216 319503 308272
rect 316677 308214 319503 308216
rect 316677 308211 316743 308214
rect 319437 308211 319503 308214
rect 297541 308138 297607 308141
rect 297950 308138 297956 308140
rect 297541 308136 297956 308138
rect 297541 308080 297546 308136
rect 297602 308080 297956 308136
rect 297541 308078 297956 308080
rect 297541 308075 297607 308078
rect 297950 308076 297956 308078
rect 298020 308076 298026 308140
rect 277342 307940 277348 308004
rect 277412 308002 277418 308004
rect 277577 308002 277643 308005
rect 277412 308000 277643 308002
rect 277412 307944 277582 308000
rect 277638 307944 277643 308000
rect 277412 307942 277643 307944
rect 277412 307940 277418 307942
rect 277577 307939 277643 307942
rect 297766 307940 297772 308004
rect 297836 308002 297842 308004
rect 298001 308002 298067 308005
rect 297836 308000 298067 308002
rect 297836 307944 298006 308000
rect 298062 307944 298067 308000
rect 297836 307942 298067 307944
rect 297836 307940 297842 307942
rect 298001 307939 298067 307942
rect 298134 307940 298140 308004
rect 298204 308002 298210 308004
rect 298921 308002 298987 308005
rect 298204 308000 298987 308002
rect 298204 307944 298926 308000
rect 298982 307944 298987 308000
rect 298204 307942 298987 307944
rect 298204 307940 298210 307942
rect 298921 307939 298987 307942
rect 314101 308002 314167 308005
rect 318057 308002 318123 308005
rect 314101 308000 318123 308002
rect 314101 307944 314106 308000
rect 314162 307944 318062 308000
rect 318118 307944 318123 308000
rect 314101 307942 318123 307944
rect 314101 307939 314167 307942
rect 318057 307939 318123 307942
rect 277393 307866 277459 307869
rect 277526 307866 277532 307868
rect 277393 307864 277532 307866
rect 277393 307808 277398 307864
rect 277454 307808 277532 307864
rect 277393 307806 277532 307808
rect 277393 307803 277459 307806
rect 277526 307804 277532 307806
rect 277596 307804 277602 307868
rect 284886 307804 284892 307868
rect 284956 307866 284962 307868
rect 285397 307866 285463 307869
rect 284956 307864 285463 307866
rect 284956 307808 285402 307864
rect 285458 307808 285463 307864
rect 284956 307806 285463 307808
rect 284956 307804 284962 307806
rect 285397 307803 285463 307806
rect 286726 307804 286732 307868
rect 286796 307866 286802 307868
rect 286961 307866 287027 307869
rect 286796 307864 287027 307866
rect 286796 307808 286966 307864
rect 287022 307808 287027 307864
rect 286796 307806 287027 307808
rect 286796 307804 286802 307806
rect 286961 307803 287027 307806
rect 293861 307866 293927 307869
rect 295977 307866 296043 307869
rect 293861 307864 296043 307866
rect 293861 307808 293866 307864
rect 293922 307808 295982 307864
rect 296038 307808 296043 307864
rect 293861 307806 296043 307808
rect 293861 307803 293927 307806
rect 295977 307803 296043 307806
rect 297173 307866 297239 307869
rect 297398 307866 297404 307868
rect 297173 307864 297404 307866
rect 297173 307808 297178 307864
rect 297234 307808 297404 307864
rect 297173 307806 297404 307808
rect 297173 307803 297239 307806
rect 297398 307804 297404 307806
rect 297468 307804 297474 307868
rect 297582 307804 297588 307868
rect 297652 307866 297658 307868
rect 297817 307866 297883 307869
rect 297652 307864 297883 307866
rect 297652 307808 297822 307864
rect 297878 307808 297883 307864
rect 297652 307806 297883 307808
rect 297652 307804 297658 307806
rect 297817 307803 297883 307806
rect 298461 307868 298527 307869
rect 298461 307864 298508 307868
rect 298572 307866 298578 307868
rect 298461 307808 298466 307864
rect 298461 307804 298508 307808
rect 298572 307806 298618 307866
rect 298572 307804 298578 307806
rect 298461 307803 298527 307804
rect 256969 306642 257035 306645
rect 256969 306640 257170 306642
rect 256969 306584 256974 306640
rect 257030 306584 257170 306640
rect 256969 306582 257170 306584
rect 256969 306579 257035 306582
rect 257110 306373 257170 306582
rect 257110 306368 257219 306373
rect -960 306234 480 306324
rect 257110 306312 257158 306368
rect 257214 306312 257219 306368
rect 257110 306310 257219 306312
rect 257153 306307 257219 306310
rect 282494 306308 282500 306372
rect 282564 306370 282570 306372
rect 338849 306370 338915 306373
rect 282564 306368 338915 306370
rect 282564 306312 338854 306368
rect 338910 306312 338915 306368
rect 282564 306310 338915 306312
rect 282564 306308 282570 306310
rect 338849 306307 338915 306310
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 279366 306172 279372 306236
rect 279436 306234 279442 306236
rect 355409 306234 355475 306237
rect 279436 306232 355475 306234
rect 279436 306176 355414 306232
rect 355470 306176 355475 306232
rect 279436 306174 355475 306176
rect 279436 306172 279442 306174
rect 355409 306171 355475 306174
rect 320725 306098 320791 306101
rect 489913 306098 489979 306101
rect 320725 306096 489979 306098
rect 320725 306040 320730 306096
rect 320786 306040 489918 306096
rect 489974 306040 489979 306096
rect 320725 306038 489979 306040
rect 320725 306035 320791 306038
rect 489913 306035 489979 306038
rect 325325 305962 325391 305965
rect 516777 305962 516843 305965
rect 325325 305960 516843 305962
rect 325325 305904 325330 305960
rect 325386 305904 516782 305960
rect 516838 305904 516843 305960
rect 325325 305902 516843 305904
rect 325325 305899 325391 305902
rect 516777 305899 516843 305902
rect 331121 305826 331187 305829
rect 332225 305826 332291 305829
rect 331121 305824 332291 305826
rect 331121 305768 331126 305824
rect 331182 305768 332230 305824
rect 332286 305768 332291 305824
rect 331121 305766 332291 305768
rect 331121 305763 331187 305766
rect 332225 305763 332291 305766
rect 336089 305826 336155 305829
rect 575473 305826 575539 305829
rect 336089 305824 575539 305826
rect 336089 305768 336094 305824
rect 336150 305768 575478 305824
rect 575534 305768 575539 305824
rect 336089 305766 575539 305768
rect 336089 305763 336155 305766
rect 575473 305763 575539 305766
rect 40677 305690 40743 305693
rect 360929 305690 360995 305693
rect 40677 305688 360995 305690
rect 40677 305632 40682 305688
rect 40738 305632 360934 305688
rect 360990 305632 360995 305688
rect 40677 305630 360995 305632
rect 40677 305627 40743 305630
rect 360929 305627 360995 305630
rect 273989 303514 274055 303517
rect 340045 303514 340111 303517
rect 273989 303512 340111 303514
rect 273989 303456 273994 303512
rect 274050 303456 340050 303512
rect 340106 303456 340111 303512
rect 273989 303454 340111 303456
rect 273989 303451 274055 303454
rect 340045 303451 340111 303454
rect 279550 303316 279556 303380
rect 279620 303378 279626 303380
rect 354857 303378 354923 303381
rect 279620 303376 354923 303378
rect 279620 303320 354862 303376
rect 354918 303320 354923 303376
rect 279620 303318 354923 303320
rect 279620 303316 279626 303318
rect 354857 303315 354923 303318
rect 312353 303242 312419 303245
rect 442349 303242 442415 303245
rect 312353 303240 442415 303242
rect 312353 303184 312358 303240
rect 312414 303184 442354 303240
rect 442410 303184 442415 303240
rect 312353 303182 442415 303184
rect 312353 303179 312419 303182
rect 442349 303179 442415 303182
rect 319161 303106 319227 303109
rect 485037 303106 485103 303109
rect 319161 303104 485103 303106
rect 319161 303048 319166 303104
rect 319222 303048 485042 303104
rect 485098 303048 485103 303104
rect 319161 303046 485103 303048
rect 319161 303043 319227 303046
rect 485037 303043 485103 303046
rect 326061 302970 326127 302973
rect 520917 302970 520983 302973
rect 326061 302968 520983 302970
rect 326061 302912 326066 302968
rect 326122 302912 520922 302968
rect 520978 302912 520983 302968
rect 326061 302910 520983 302912
rect 326061 302907 326127 302910
rect 520917 302907 520983 302910
rect 330293 302834 330359 302837
rect 545113 302834 545179 302837
rect 330293 302832 545179 302834
rect 330293 302776 330298 302832
rect 330354 302776 545118 302832
rect 545174 302776 545179 302832
rect 330293 302774 545179 302776
rect 330293 302771 330359 302774
rect 545113 302771 545179 302774
rect 280061 300794 280127 300797
rect 350717 300794 350783 300797
rect 280061 300792 350783 300794
rect 280061 300736 280066 300792
rect 280122 300736 350722 300792
rect 350778 300736 350783 300792
rect 280061 300734 350783 300736
rect 280061 300731 280127 300734
rect 350717 300731 350783 300734
rect 278589 300658 278655 300661
rect 354765 300658 354831 300661
rect 278589 300656 354831 300658
rect 278589 300600 278594 300656
rect 278650 300600 354770 300656
rect 354826 300600 354831 300656
rect 278589 300598 354831 300600
rect 278589 300595 278655 300598
rect 354765 300595 354831 300598
rect 268653 300522 268719 300525
rect 345289 300522 345355 300525
rect 268653 300520 345355 300522
rect 268653 300464 268658 300520
rect 268714 300464 345294 300520
rect 345350 300464 345355 300520
rect 268653 300462 345355 300464
rect 268653 300459 268719 300462
rect 345289 300459 345355 300462
rect 316309 300386 316375 300389
rect 471237 300386 471303 300389
rect 316309 300384 471303 300386
rect 316309 300328 316314 300384
rect 316370 300328 471242 300384
rect 471298 300328 471303 300384
rect 316309 300326 471303 300328
rect 316309 300323 316375 300326
rect 471237 300323 471303 300326
rect 320541 300250 320607 300253
rect 498285 300250 498351 300253
rect 320541 300248 498351 300250
rect 320541 300192 320546 300248
rect 320602 300192 498290 300248
rect 498346 300192 498351 300248
rect 320541 300190 498351 300192
rect 320541 300187 320607 300190
rect 498285 300187 498351 300190
rect 330201 300114 330267 300117
rect 543733 300114 543799 300117
rect 330201 300112 543799 300114
rect 330201 300056 330206 300112
rect 330262 300056 543738 300112
rect 543794 300056 543799 300112
rect 330201 300054 543799 300056
rect 330201 300051 330267 300054
rect 543733 300051 543799 300054
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 310881 287738 310947 287741
rect 439078 287738 439084 287740
rect 310881 287736 439084 287738
rect 310881 287680 310886 287736
rect 310942 287680 439084 287736
rect 310881 287678 439084 287680
rect 310881 287675 310947 287678
rect 439078 287676 439084 287678
rect 439148 287676 439154 287740
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 309593 275226 309659 275229
rect 437422 275226 437428 275228
rect 309593 275224 437428 275226
rect 309593 275168 309598 275224
rect 309654 275168 437428 275224
rect 309593 275166 437428 275168
rect 309593 275163 309659 275166
rect 437422 275164 437428 275166
rect 437492 275164 437498 275228
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 293350 248236 293356 248300
rect 293420 248298 293426 248300
rect 301129 248298 301195 248301
rect 293420 248296 301195 248298
rect 293420 248240 301134 248296
rect 301190 248240 301195 248296
rect 293420 248238 301195 248240
rect 293420 248236 293426 248238
rect 301129 248235 301195 248238
rect 289486 248100 289492 248164
rect 289556 248162 289562 248164
rect 299933 248162 299999 248165
rect 289556 248160 299999 248162
rect 289556 248104 299938 248160
rect 299994 248104 299999 248160
rect 289556 248102 299999 248104
rect 289556 248100 289562 248102
rect 299933 248099 299999 248102
rect 288198 247964 288204 248028
rect 288268 248026 288274 248028
rect 301221 248026 301287 248029
rect 288268 248024 301287 248026
rect 288268 247968 301226 248024
rect 301282 247968 301287 248024
rect 288268 247966 301287 247968
rect 288268 247964 288274 247966
rect 301221 247963 301287 247966
rect 289302 247828 289308 247892
rect 289372 247890 289378 247892
rect 302509 247890 302575 247893
rect 289372 247888 302575 247890
rect 289372 247832 302514 247888
rect 302570 247832 302575 247888
rect 289372 247830 302575 247832
rect 289372 247828 289378 247830
rect 302509 247827 302575 247830
rect 288014 247692 288020 247756
rect 288084 247754 288090 247756
rect 302601 247754 302667 247757
rect 288084 247752 302667 247754
rect 288084 247696 302606 247752
rect 302662 247696 302667 247752
rect 288084 247694 302667 247696
rect 288084 247692 288090 247694
rect 302601 247691 302667 247694
rect 285070 247556 285076 247620
rect 285140 247618 285146 247620
rect 302693 247618 302759 247621
rect 285140 247616 302759 247618
rect 285140 247560 302698 247616
rect 302754 247560 302759 247616
rect 285140 247558 302759 247560
rect 285140 247556 285146 247558
rect 302693 247555 302759 247558
rect 309409 247618 309475 247621
rect 437606 247618 437612 247620
rect 309409 247616 437612 247618
rect 309409 247560 309414 247616
rect 309470 247560 437612 247616
rect 309409 247558 437612 247560
rect 309409 247555 309475 247558
rect 437606 247556 437612 247558
rect 437676 247556 437682 247620
rect 296110 247420 296116 247484
rect 296180 247482 296186 247484
rect 299841 247482 299907 247485
rect 296180 247480 299907 247482
rect 296180 247424 299846 247480
rect 299902 247424 299907 247480
rect 296180 247422 299907 247424
rect 296180 247420 296186 247422
rect 299841 247419 299907 247422
rect 284518 247148 284524 247212
rect 284588 247210 284594 247212
rect 285581 247210 285647 247213
rect 284588 247208 285647 247210
rect 284588 247152 285586 247208
rect 285642 247152 285647 247208
rect 284588 247150 285647 247152
rect 284588 247148 284594 247150
rect 285581 247147 285647 247150
rect 287646 247148 287652 247212
rect 287716 247210 287722 247212
rect 287973 247210 288039 247213
rect 287716 247208 288039 247210
rect 287716 247152 287978 247208
rect 288034 247152 288039 247208
rect 287716 247150 288039 247152
rect 287716 247148 287722 247150
rect 287973 247147 288039 247150
rect 288934 247148 288940 247212
rect 289004 247210 289010 247212
rect 289353 247210 289419 247213
rect 289004 247208 289419 247210
rect 289004 247152 289358 247208
rect 289414 247152 289419 247208
rect 289004 247150 289419 247152
rect 289004 247148 289010 247150
rect 289353 247147 289419 247150
rect 284753 247076 284819 247077
rect 284702 247074 284708 247076
rect 284662 247014 284708 247074
rect 284772 247072 284819 247076
rect 284814 247016 284819 247072
rect 284702 247012 284708 247014
rect 284772 247012 284819 247016
rect 286358 247012 286364 247076
rect 286428 247074 286434 247076
rect 286685 247074 286751 247077
rect 286961 247076 287027 247077
rect 287881 247076 287947 247077
rect 289169 247076 289235 247077
rect 286910 247074 286916 247076
rect 286428 247072 286751 247074
rect 286428 247016 286690 247072
rect 286746 247016 286751 247072
rect 286428 247014 286751 247016
rect 286870 247014 286916 247074
rect 286980 247072 287027 247076
rect 287830 247074 287836 247076
rect 287022 247016 287027 247072
rect 286428 247012 286434 247014
rect 284753 247011 284819 247012
rect 286685 247011 286751 247014
rect 286910 247012 286916 247014
rect 286980 247012 287027 247016
rect 287790 247014 287836 247074
rect 287900 247072 287947 247076
rect 289118 247074 289124 247076
rect 287942 247016 287947 247072
rect 287830 247012 287836 247014
rect 287900 247012 287947 247016
rect 289078 247014 289124 247074
rect 289188 247072 289235 247076
rect 289230 247016 289235 247072
rect 289118 247012 289124 247014
rect 289188 247012 289235 247016
rect 286961 247011 287027 247012
rect 287881 247011 287947 247012
rect 289169 247011 289235 247012
rect 299105 245578 299171 245581
rect 358854 245578 358860 245580
rect 299105 245576 358860 245578
rect 299105 245520 299110 245576
rect 299166 245520 358860 245576
rect 299105 245518 358860 245520
rect 299105 245515 299171 245518
rect 358854 245516 358860 245518
rect 358924 245516 358930 245580
rect 583520 245428 584960 245668
rect 293534 245244 293540 245308
rect 293604 245306 293610 245308
rect 302233 245306 302299 245309
rect 293604 245304 302299 245306
rect 293604 245248 302238 245304
rect 302294 245248 302299 245304
rect 293604 245246 302299 245248
rect 293604 245244 293610 245246
rect 302233 245243 302299 245246
rect 290958 245108 290964 245172
rect 291028 245170 291034 245172
rect 301037 245170 301103 245173
rect 291028 245168 301103 245170
rect 291028 245112 301042 245168
rect 301098 245112 301103 245168
rect 291028 245110 301103 245112
rect 291028 245108 291034 245110
rect 301037 245107 301103 245110
rect 309133 245170 309199 245173
rect 437790 245170 437796 245172
rect 309133 245168 437796 245170
rect 309133 245112 309138 245168
rect 309194 245112 437796 245168
rect 309133 245110 437796 245112
rect 309133 245107 309199 245110
rect 437790 245108 437796 245110
rect 437860 245108 437866 245172
rect 284150 244972 284156 245036
rect 284220 245034 284226 245036
rect 296805 245034 296871 245037
rect 284220 245032 296871 245034
rect 284220 244976 296810 245032
rect 296866 244976 296871 245032
rect 284220 244974 296871 244976
rect 284220 244972 284226 244974
rect 296805 244971 296871 244974
rect 297081 245034 297147 245037
rect 299657 245034 299723 245037
rect 297081 245032 299723 245034
rect 297081 244976 297086 245032
rect 297142 244976 299662 245032
rect 299718 244976 299723 245032
rect 297081 244974 299723 244976
rect 297081 244971 297147 244974
rect 299657 244971 299723 244974
rect 309317 245034 309383 245037
rect 439262 245034 439268 245036
rect 309317 245032 439268 245034
rect 309317 244976 309322 245032
rect 309378 244976 439268 245032
rect 309317 244974 439268 244976
rect 309317 244971 309383 244974
rect 439262 244972 439268 244974
rect 439332 244972 439338 245036
rect 283966 244836 283972 244900
rect 284036 244898 284042 244900
rect 298185 244898 298251 244901
rect 284036 244896 298251 244898
rect 284036 244840 298190 244896
rect 298246 244840 298251 244896
rect 284036 244838 298251 244840
rect 284036 244836 284042 244838
rect 298185 244835 298251 244838
rect 328453 244898 328519 244901
rect 539685 244898 539751 244901
rect 328453 244896 539751 244898
rect 328453 244840 328458 244896
rect 328514 244840 539690 244896
rect 539746 244840 539751 244896
rect 328453 244838 539751 244840
rect 328453 244835 328519 244838
rect 539685 244835 539751 244838
rect 292430 244700 292436 244764
rect 292500 244762 292506 244764
rect 299473 244762 299539 244765
rect 292500 244760 299539 244762
rect 292500 244704 299478 244760
rect 299534 244704 299539 244760
rect 292500 244702 299539 244704
rect 292500 244700 292506 244702
rect 299473 244699 299539 244702
rect 295926 244564 295932 244628
rect 295996 244626 296002 244628
rect 297081 244626 297147 244629
rect 295996 244624 297147 244626
rect 295996 244568 297086 244624
rect 297142 244568 297147 244624
rect 295996 244566 297147 244568
rect 295996 244564 296002 244566
rect 297081 244563 297147 244566
rect 297398 244564 297404 244628
rect 297468 244626 297474 244628
rect 298737 244626 298803 244629
rect 297468 244624 298803 244626
rect 297468 244568 298742 244624
rect 298798 244568 298803 244624
rect 297468 244566 298803 244568
rect 297468 244564 297474 244566
rect 298737 244563 298803 244566
rect 292246 244428 292252 244492
rect 292316 244490 292322 244492
rect 298277 244490 298343 244493
rect 298686 244490 298692 244492
rect 292316 244430 298202 244490
rect 292316 244428 292322 244430
rect 290641 244356 290707 244357
rect 291745 244356 291811 244357
rect 292113 244356 292179 244357
rect 290590 244354 290596 244356
rect 290550 244294 290596 244354
rect 290660 244352 290707 244356
rect 291694 244354 291700 244356
rect 290702 244296 290707 244352
rect 290590 244292 290596 244294
rect 290660 244292 290707 244296
rect 291654 244294 291700 244354
rect 291764 244352 291811 244356
rect 292062 244354 292068 244356
rect 291806 244296 291811 244352
rect 291694 244292 291700 244294
rect 291764 244292 291811 244296
rect 292022 244294 292068 244354
rect 292132 244352 292179 244356
rect 292174 244296 292179 244352
rect 292062 244292 292068 244294
rect 292132 244292 292179 244296
rect 293166 244292 293172 244356
rect 293236 244354 293242 244356
rect 293401 244354 293467 244357
rect 293769 244356 293835 244357
rect 295057 244356 295123 244357
rect 293718 244354 293724 244356
rect 293236 244352 293467 244354
rect 293236 244296 293406 244352
rect 293462 244296 293467 244352
rect 293236 244294 293467 244296
rect 293678 244294 293724 244354
rect 293788 244352 293835 244356
rect 295006 244354 295012 244356
rect 293830 244296 293835 244352
rect 293236 244292 293242 244294
rect 290641 244291 290707 244292
rect 291745 244291 291811 244292
rect 292113 244291 292179 244292
rect 293401 244291 293467 244294
rect 293718 244292 293724 244294
rect 293788 244292 293835 244296
rect 294966 244294 295012 244354
rect 295076 244352 295123 244356
rect 295118 244296 295123 244352
rect 295006 244292 295012 244294
rect 295076 244292 295123 244296
rect 297214 244292 297220 244356
rect 297284 244354 297290 244356
rect 297817 244354 297883 244357
rect 297284 244352 297883 244354
rect 297284 244296 297822 244352
rect 297878 244296 297883 244352
rect 297284 244294 297883 244296
rect 297284 244292 297290 244294
rect 293769 244291 293835 244292
rect 295057 244291 295123 244292
rect 297817 244291 297883 244294
rect 298142 244218 298202 244430
rect 298277 244488 298692 244490
rect 298277 244432 298282 244488
rect 298338 244432 298692 244488
rect 298277 244430 298692 244432
rect 298277 244427 298343 244430
rect 298686 244428 298692 244430
rect 298756 244428 298762 244492
rect 298369 244356 298435 244357
rect 298318 244354 298324 244356
rect 298278 244294 298324 244354
rect 298388 244352 298435 244356
rect 300945 244354 301011 244357
rect 298430 244296 298435 244352
rect 298318 244292 298324 244294
rect 298388 244292 298435 244296
rect 298369 244291 298435 244292
rect 298510 244352 301011 244354
rect 298510 244296 300950 244352
rect 301006 244296 301011 244352
rect 298510 244294 301011 244296
rect 298510 244218 298570 244294
rect 300945 244291 301011 244294
rect 298142 244158 298570 244218
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 97809 196890 97875 196893
rect 99422 196890 100004 196924
rect 97809 196888 100004 196890
rect 97809 196832 97814 196888
rect 97870 196864 100004 196888
rect 298645 196890 298711 196893
rect 299430 196890 300012 196924
rect 298645 196888 300012 196890
rect 97870 196832 99482 196864
rect 97809 196830 99482 196832
rect 298645 196832 298650 196888
rect 298706 196864 300012 196888
rect 298706 196832 299490 196864
rect 298645 196830 299490 196832
rect 97809 196827 97875 196830
rect 298645 196827 298711 196830
rect 293166 196012 293172 196076
rect 293236 196074 293242 196076
rect 293861 196074 293927 196077
rect 293236 196072 293927 196074
rect 293236 196016 293866 196072
rect 293922 196016 293927 196072
rect 293236 196014 293927 196016
rect 293236 196012 293242 196014
rect 293861 196011 293927 196014
rect 97901 195938 97967 195941
rect 99422 195938 100004 195972
rect 97901 195936 100004 195938
rect 97901 195880 97906 195936
rect 97962 195912 100004 195936
rect 297357 195938 297423 195941
rect 299430 195938 300012 195972
rect 297357 195936 300012 195938
rect 97962 195880 99482 195912
rect 97901 195878 99482 195880
rect 297357 195880 297362 195936
rect 297418 195912 300012 195936
rect 297418 195880 299490 195912
rect 297357 195878 299490 195880
rect 97901 195875 97967 195878
rect 297357 195875 297423 195878
rect 97901 193762 97967 193765
rect 99422 193762 100004 193796
rect 97901 193760 100004 193762
rect 97901 193704 97906 193760
rect 97962 193736 100004 193760
rect 298829 193762 298895 193765
rect 299430 193762 300012 193796
rect 298829 193760 300012 193762
rect 97962 193704 99482 193736
rect 97901 193702 99482 193704
rect 298829 193704 298834 193760
rect 298890 193736 300012 193760
rect 298890 193704 299490 193736
rect 298829 193702 299490 193704
rect 97901 193699 97967 193702
rect 298829 193699 298895 193702
rect 297357 193218 297423 193221
rect 297541 193218 297607 193221
rect 297357 193216 297607 193218
rect 297357 193160 297362 193216
rect 297418 193160 297546 193216
rect 297602 193160 297607 193216
rect 297357 193158 297607 193160
rect 297357 193155 297423 193158
rect 297541 193155 297607 193158
rect 97809 192810 97875 192813
rect 99422 192810 100004 192844
rect 97809 192808 100004 192810
rect 97809 192752 97814 192808
rect 97870 192784 100004 192808
rect 297357 192810 297423 192813
rect 299430 192810 300012 192844
rect 297357 192808 300012 192810
rect 97870 192752 99482 192784
rect 97809 192750 99482 192752
rect 297357 192752 297362 192808
rect 297418 192784 300012 192808
rect 297418 192752 299490 192784
rect 297357 192750 299490 192752
rect 97809 192747 97875 192750
rect 297357 192747 297423 192750
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 97717 191042 97783 191045
rect 99422 191042 100004 191076
rect 97717 191040 100004 191042
rect 97717 190984 97722 191040
rect 97778 191016 100004 191040
rect 297449 191042 297515 191045
rect 299430 191042 300012 191076
rect 297449 191040 300012 191042
rect 97778 190984 99482 191016
rect 97717 190982 99482 190984
rect 297449 190984 297454 191040
rect 297510 191016 300012 191040
rect 297510 190984 299490 191016
rect 297449 190982 299490 190984
rect 97717 190979 97783 190982
rect 297449 190979 297515 190982
rect 97625 189954 97691 189957
rect 99422 189954 100004 189988
rect 97625 189952 100004 189954
rect 97625 189896 97630 189952
rect 97686 189928 100004 189952
rect 297541 189954 297607 189957
rect 299430 189954 300012 189988
rect 297541 189952 300012 189954
rect 97686 189896 99482 189928
rect 97625 189894 99482 189896
rect 297541 189896 297546 189952
rect 297602 189928 300012 189952
rect 297602 189896 299490 189928
rect 297541 189894 299490 189896
rect 97625 189891 97691 189894
rect 297541 189891 297607 189894
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 97533 188186 97599 188189
rect 99422 188186 100004 188220
rect 97533 188184 100004 188186
rect 97533 188128 97538 188184
rect 97594 188160 100004 188184
rect 297633 188186 297699 188189
rect 298921 188186 298987 188189
rect 299430 188186 300012 188220
rect 297633 188184 300012 188186
rect 97594 188128 99482 188160
rect 97533 188126 99482 188128
rect 297633 188128 297638 188184
rect 297694 188128 298926 188184
rect 298982 188160 300012 188184
rect 298982 188128 299490 188160
rect 297633 188126 299490 188128
rect 97533 188123 97599 188126
rect 297633 188123 297699 188126
rect 298921 188123 298987 188126
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 97441 169962 97507 169965
rect 99422 169962 100004 169996
rect 97441 169960 100004 169962
rect 97441 169904 97446 169960
rect 97502 169936 100004 169960
rect 298001 169962 298067 169965
rect 299430 169962 300012 169996
rect 298001 169960 300012 169962
rect 97502 169904 99482 169936
rect 97441 169902 99482 169904
rect 298001 169904 298006 169960
rect 298062 169936 300012 169960
rect 298062 169904 299490 169936
rect 298001 169902 299490 169904
rect 97441 169899 97507 169902
rect 298001 169899 298067 169902
rect 284518 169764 284524 169828
rect 284588 169826 284594 169828
rect 285581 169826 285647 169829
rect 284588 169824 285647 169826
rect 284588 169768 285586 169824
rect 285642 169768 285647 169824
rect 284588 169766 285647 169768
rect 284588 169764 284594 169766
rect 285581 169763 285647 169766
rect 294873 168466 294939 168469
rect 295006 168466 295012 168468
rect 294873 168464 295012 168466
rect 294873 168408 294878 168464
rect 294934 168408 295012 168464
rect 294873 168406 295012 168408
rect 294873 168403 294939 168406
rect 295006 168404 295012 168406
rect 295076 168404 295082 168468
rect 97349 168330 97415 168333
rect 99422 168330 100004 168364
rect 97349 168328 100004 168330
rect 97349 168272 97354 168328
rect 97410 168304 100004 168328
rect 297725 168330 297791 168333
rect 299430 168330 300012 168364
rect 297725 168328 300012 168330
rect 97410 168272 99482 168304
rect 97349 168270 99482 168272
rect 297725 168272 297730 168328
rect 297786 168304 300012 168328
rect 297786 168272 299490 168304
rect 297725 168270 299490 168272
rect 97349 168267 97415 168270
rect 297725 168267 297791 168270
rect 99281 168058 99347 168061
rect 99422 168058 100004 168092
rect 299430 168061 300012 168092
rect 99281 168056 100004 168058
rect 99281 168000 99286 168056
rect 99342 168032 100004 168056
rect 299381 168056 300012 168061
rect 99342 168000 99482 168032
rect 99281 167998 99482 168000
rect 299381 168000 299386 168056
rect 299442 168032 300012 168056
rect 299442 168000 299490 168032
rect 299381 167998 299490 168000
rect 99281 167995 99347 167998
rect 299381 167995 299447 167998
rect 297214 167044 297220 167108
rect 297284 167106 297290 167108
rect 298001 167106 298067 167109
rect 297284 167104 298067 167106
rect 297284 167048 298006 167104
rect 298062 167048 298067 167104
rect 297284 167046 298067 167048
rect 297284 167044 297290 167046
rect 298001 167043 298067 167046
rect 298686 167044 298692 167108
rect 298756 167106 298762 167108
rect 299381 167106 299447 167109
rect 298756 167104 299447 167106
rect 298756 167048 299386 167104
rect 299442 167048 299447 167104
rect 298756 167046 299447 167048
rect 298756 167044 298762 167046
rect 299381 167043 299447 167046
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 260189 160714 260255 160717
rect 277526 160714 277532 160716
rect 260189 160712 277532 160714
rect 260189 160656 260194 160712
rect 260250 160656 277532 160712
rect 260189 160654 277532 160656
rect 260189 160651 260255 160654
rect 277526 160652 277532 160654
rect 277596 160652 277602 160716
rect 160921 159900 160987 159901
rect 163497 159900 163563 159901
rect 165981 159900 166047 159901
rect 203425 159900 203491 159901
rect 160921 159896 160934 159900
rect 160998 159898 161004 159900
rect 160921 159840 160926 159896
rect 160921 159836 160934 159840
rect 160998 159838 161078 159898
rect 163497 159896 163518 159900
rect 163582 159898 163588 159900
rect 165960 159898 165966 159900
rect 163497 159840 163502 159896
rect 160998 159836 161004 159838
rect 163497 159836 163518 159840
rect 163582 159838 163654 159898
rect 165890 159838 165966 159898
rect 166030 159896 166047 159900
rect 203360 159898 203366 159900
rect 166042 159840 166047 159896
rect 163582 159836 163588 159838
rect 165960 159836 165966 159838
rect 166030 159836 166047 159840
rect 203334 159838 203366 159898
rect 203360 159836 203366 159838
rect 203430 159896 203491 159900
rect 203486 159840 203491 159896
rect 203430 159836 203491 159840
rect 160921 159835 160987 159836
rect 163497 159835 163563 159836
rect 165981 159835 166047 159836
rect 203425 159835 203491 159836
rect 345933 159900 345999 159901
rect 348233 159900 348299 159901
rect 353569 159900 353635 159901
rect 365897 159900 365963 159901
rect 345933 159896 345974 159900
rect 346038 159898 346044 159900
rect 345933 159840 345938 159896
rect 345933 159836 345974 159840
rect 346038 159838 346090 159898
rect 348233 159896 348286 159900
rect 348350 159898 348356 159900
rect 348233 159840 348238 159896
rect 346038 159836 346044 159838
rect 348233 159836 348286 159840
rect 348350 159838 348390 159898
rect 353569 159896 353590 159900
rect 353654 159898 353660 159900
rect 353569 159840 353574 159896
rect 348350 159836 348356 159838
rect 353569 159836 353590 159840
rect 353654 159838 353726 159898
rect 365897 159896 365966 159900
rect 365897 159840 365902 159896
rect 365958 159840 365966 159896
rect 353654 159836 353660 159838
rect 365897 159836 365966 159840
rect 366030 159898 366036 159900
rect 366030 159838 366054 159898
rect 366030 159836 366036 159838
rect 345933 159835 345999 159836
rect 348233 159835 348299 159836
rect 353569 159835 353635 159836
rect 365897 159835 365963 159836
rect 350993 159764 351059 159765
rect 350993 159760 351006 159764
rect 351070 159762 351076 159764
rect 350993 159704 350998 159760
rect 350993 159700 351006 159704
rect 351070 159702 351150 159762
rect 351070 159700 351076 159702
rect 350993 159699 351059 159700
rect 356053 159628 356119 159629
rect 356032 159626 356038 159628
rect 355962 159566 356038 159626
rect 356102 159624 356119 159628
rect 356114 159568 356119 159624
rect 356032 159564 356038 159566
rect 356102 159564 356119 159568
rect 356053 159563 356119 159564
rect 358445 159628 358511 159629
rect 358445 159624 358486 159628
rect 358550 159626 358556 159628
rect 358445 159568 358450 159624
rect 358445 159564 358486 159568
rect 358550 159566 358602 159626
rect 358550 159564 358556 159566
rect 358445 159563 358511 159564
rect 213913 159490 213979 159493
rect 269665 159490 269731 159493
rect 213913 159488 269731 159490
rect 213913 159432 213918 159488
rect 213974 159432 269670 159488
rect 269726 159432 269731 159488
rect 213913 159430 269731 159432
rect 213913 159427 213979 159430
rect 269665 159427 269731 159430
rect 200113 159354 200179 159357
rect 265617 159354 265683 159357
rect 200113 159352 265683 159354
rect 200113 159296 200118 159352
rect 200174 159296 265622 159352
rect 265678 159296 265683 159352
rect 200113 159294 265683 159296
rect 200113 159291 200179 159294
rect 265617 159291 265683 159294
rect 298134 159292 298140 159356
rect 298204 159354 298210 159356
rect 373993 159354 374059 159357
rect 298204 159352 374059 159354
rect 298204 159296 373998 159352
rect 374054 159296 374059 159352
rect 298204 159294 374059 159296
rect 298204 159292 298210 159294
rect 373993 159291 374059 159294
rect 153694 159156 153700 159220
rect 153764 159218 153770 159220
rect 247769 159218 247835 159221
rect 153764 159216 247835 159218
rect 153764 159160 247774 159216
rect 247830 159160 247835 159216
rect 153764 159158 247835 159160
rect 153764 159156 153770 159158
rect 247769 159155 247835 159158
rect 128302 159020 128308 159084
rect 128372 159082 128378 159084
rect 238017 159082 238083 159085
rect 128372 159080 238083 159082
rect 128372 159024 238022 159080
rect 238078 159024 238083 159080
rect 128372 159022 238083 159024
rect 128372 159020 128378 159022
rect 238017 159019 238083 159022
rect 287646 159020 287652 159084
rect 287716 159082 287722 159084
rect 288065 159082 288131 159085
rect 287716 159080 288131 159082
rect 287716 159024 288070 159080
rect 288126 159024 288131 159080
rect 287716 159022 288131 159024
rect 287716 159020 287722 159022
rect 288065 159019 288131 159022
rect 173382 158884 173388 158948
rect 173452 158946 173458 158948
rect 286174 158946 286180 158948
rect 173452 158886 286180 158946
rect 173452 158884 173458 158886
rect 286174 158884 286180 158886
rect 286244 158884 286250 158948
rect 287830 158884 287836 158948
rect 287900 158946 287906 158948
rect 287973 158946 288039 158949
rect 287900 158944 288039 158946
rect 287900 158888 287978 158944
rect 288034 158888 288039 158944
rect 287900 158886 288039 158888
rect 287900 158884 287906 158886
rect 287973 158883 288039 158886
rect 288934 158884 288940 158948
rect 289004 158946 289010 158948
rect 289721 158946 289787 158949
rect 289004 158944 289787 158946
rect 289004 158888 289726 158944
rect 289782 158888 289787 158944
rect 289004 158886 289787 158888
rect 289004 158884 289010 158886
rect 289721 158883 289787 158886
rect 156086 158748 156092 158812
rect 156156 158810 156162 158812
rect 282126 158810 282132 158812
rect 156156 158750 282132 158810
rect 156156 158748 156162 158750
rect 282126 158748 282132 158750
rect 282196 158748 282202 158812
rect 284702 158748 284708 158812
rect 284772 158810 284778 158812
rect 285397 158810 285463 158813
rect 284772 158808 285463 158810
rect 284772 158752 285402 158808
rect 285458 158752 285463 158808
rect 284772 158750 285463 158752
rect 284772 158748 284778 158750
rect 285397 158747 285463 158750
rect 286358 158748 286364 158812
rect 286428 158810 286434 158812
rect 286961 158810 287027 158813
rect 286428 158808 287027 158810
rect 286428 158752 286966 158808
rect 287022 158752 287027 158808
rect 286428 158750 287027 158752
rect 286428 158748 286434 158750
rect 286961 158747 287027 158750
rect 287881 158810 287947 158813
rect 288014 158810 288020 158812
rect 287881 158808 288020 158810
rect 287881 158752 287886 158808
rect 287942 158752 288020 158808
rect 287881 158750 288020 158752
rect 287881 158747 287947 158750
rect 288014 158748 288020 158750
rect 288084 158748 288090 158812
rect 289118 158748 289124 158812
rect 289188 158810 289194 158812
rect 289353 158810 289419 158813
rect 290641 158812 290707 158813
rect 290590 158810 290596 158812
rect 289188 158808 289419 158810
rect 289188 158752 289358 158808
rect 289414 158752 289419 158808
rect 289188 158750 289419 158752
rect 290550 158750 290596 158810
rect 290660 158808 290707 158812
rect 290702 158752 290707 158808
rect 289188 158748 289194 158750
rect 289353 158747 289419 158750
rect 290590 158748 290596 158750
rect 290660 158748 290707 158752
rect 291694 158748 291700 158812
rect 291764 158810 291770 158812
rect 292481 158810 292547 158813
rect 291764 158808 292547 158810
rect 291764 158752 292486 158808
rect 292542 158752 292547 158808
rect 291764 158750 292547 158752
rect 291764 158748 291770 158750
rect 290641 158747 290707 158748
rect 292481 158747 292547 158750
rect 116158 158612 116164 158676
rect 116228 158674 116234 158676
rect 116853 158674 116919 158677
rect 119705 158676 119771 158677
rect 119654 158674 119660 158676
rect 116228 158672 116919 158674
rect 116228 158616 116858 158672
rect 116914 158616 116919 158672
rect 116228 158614 116919 158616
rect 119614 158614 119660 158674
rect 119724 158672 119771 158676
rect 119766 158616 119771 158672
rect 116228 158612 116234 158614
rect 116853 158611 116919 158614
rect 119654 158612 119660 158614
rect 119724 158612 119771 158616
rect 120574 158612 120580 158676
rect 120644 158674 120650 158676
rect 121177 158674 121243 158677
rect 120644 158672 121243 158674
rect 120644 158616 121182 158672
rect 121238 158616 121243 158672
rect 120644 158614 121243 158616
rect 120644 158612 120650 158614
rect 119705 158611 119771 158612
rect 121177 158611 121243 158614
rect 121862 158612 121868 158676
rect 121932 158674 121938 158676
rect 122097 158674 122163 158677
rect 123201 158676 123267 158677
rect 123150 158674 123156 158676
rect 121932 158672 122163 158674
rect 121932 158616 122102 158672
rect 122158 158616 122163 158672
rect 121932 158614 122163 158616
rect 123110 158614 123156 158674
rect 123220 158672 123267 158676
rect 123262 158616 123267 158672
rect 121932 158612 121938 158614
rect 122097 158611 122163 158614
rect 123150 158612 123156 158614
rect 123220 158612 123267 158616
rect 124254 158612 124260 158676
rect 124324 158674 124330 158676
rect 125317 158674 125383 158677
rect 126513 158676 126579 158677
rect 127617 158676 127683 158677
rect 128721 158676 128787 158677
rect 130193 158676 130259 158677
rect 131297 158676 131363 158677
rect 132401 158676 132467 158677
rect 133505 158676 133571 158677
rect 126462 158674 126468 158676
rect 124324 158672 125383 158674
rect 124324 158616 125322 158672
rect 125378 158616 125383 158672
rect 124324 158614 125383 158616
rect 126422 158614 126468 158674
rect 126532 158672 126579 158676
rect 127566 158674 127572 158676
rect 126574 158616 126579 158672
rect 124324 158612 124330 158614
rect 123201 158611 123267 158612
rect 125317 158611 125383 158614
rect 126462 158612 126468 158614
rect 126532 158612 126579 158616
rect 127526 158614 127572 158674
rect 127636 158672 127683 158676
rect 128670 158674 128676 158676
rect 127678 158616 127683 158672
rect 127566 158612 127572 158614
rect 127636 158612 127683 158616
rect 128630 158614 128676 158674
rect 128740 158672 128787 158676
rect 130142 158674 130148 158676
rect 128782 158616 128787 158672
rect 128670 158612 128676 158614
rect 128740 158612 128787 158616
rect 130102 158614 130148 158674
rect 130212 158672 130259 158676
rect 131246 158674 131252 158676
rect 130254 158616 130259 158672
rect 130142 158612 130148 158614
rect 130212 158612 130259 158616
rect 131206 158614 131252 158674
rect 131316 158672 131363 158676
rect 132350 158674 132356 158676
rect 131358 158616 131363 158672
rect 131246 158612 131252 158614
rect 131316 158612 131363 158616
rect 132310 158614 132356 158674
rect 132420 158672 132467 158676
rect 133454 158674 133460 158676
rect 132462 158616 132467 158672
rect 132350 158612 132356 158614
rect 132420 158612 132467 158616
rect 133414 158614 133460 158674
rect 133524 158672 133571 158676
rect 133566 158616 133571 158672
rect 133454 158612 133460 158614
rect 133524 158612 133571 158616
rect 134558 158612 134564 158676
rect 134628 158674 134634 158676
rect 134885 158674 134951 158677
rect 158161 158676 158227 158677
rect 158529 158676 158595 158677
rect 158110 158674 158116 158676
rect 134628 158672 134951 158674
rect 134628 158616 134890 158672
rect 134946 158616 134951 158672
rect 134628 158614 134951 158616
rect 158070 158614 158116 158674
rect 158180 158672 158227 158676
rect 158478 158674 158484 158676
rect 158222 158616 158227 158672
rect 134628 158612 134634 158614
rect 126513 158611 126579 158612
rect 127617 158611 127683 158612
rect 128721 158611 128787 158612
rect 130193 158611 130259 158612
rect 131297 158611 131363 158612
rect 132401 158611 132467 158612
rect 133505 158611 133571 158612
rect 134885 158611 134951 158614
rect 158110 158612 158116 158614
rect 158180 158612 158227 158616
rect 158438 158614 158484 158674
rect 158548 158672 158595 158676
rect 158590 158616 158595 158672
rect 158478 158612 158484 158614
rect 158548 158612 158595 158616
rect 159214 158612 159220 158676
rect 159284 158674 159290 158676
rect 159817 158674 159883 158677
rect 168281 158676 168347 158677
rect 191097 158676 191163 158677
rect 168230 158674 168236 158676
rect 159284 158672 159883 158674
rect 159284 158616 159822 158672
rect 159878 158616 159883 158672
rect 159284 158614 159883 158616
rect 168190 158614 168236 158674
rect 168300 158672 168347 158676
rect 191046 158674 191052 158676
rect 168342 158616 168347 158672
rect 159284 158612 159290 158614
rect 158161 158611 158227 158612
rect 158529 158611 158595 158612
rect 159817 158611 159883 158614
rect 168230 158612 168236 158614
rect 168300 158612 168347 158616
rect 191006 158614 191052 158674
rect 191116 158672 191163 158676
rect 191158 158616 191163 158672
rect 191046 158612 191052 158614
rect 191116 158612 191163 158616
rect 168281 158611 168347 158612
rect 191097 158611 191163 158612
rect 299105 158674 299171 158677
rect 299565 158674 299631 158677
rect 299105 158672 299631 158674
rect 299105 158616 299110 158672
rect 299166 158616 299570 158672
rect 299626 158616 299631 158672
rect 299105 158614 299631 158616
rect 299105 158611 299171 158614
rect 299565 158611 299631 158614
rect 315798 158612 315804 158676
rect 315868 158674 315874 158676
rect 316033 158674 316099 158677
rect 315868 158672 316099 158674
rect 315868 158616 316038 158672
rect 316094 158616 316099 158672
rect 315868 158614 316099 158616
rect 315868 158612 315874 158614
rect 316033 158611 316099 158614
rect 316677 158674 316743 158677
rect 319437 158676 319503 158677
rect 320541 158676 320607 158677
rect 323117 158676 323183 158677
rect 324221 158676 324287 158677
rect 326429 158676 326495 158677
rect 328269 158676 328335 158677
rect 328637 158676 328703 158677
rect 329925 158676 329991 158677
rect 317086 158674 317092 158676
rect 316677 158672 317092 158674
rect 316677 158616 316682 158672
rect 316738 158616 317092 158672
rect 316677 158614 317092 158616
rect 316677 158611 316743 158614
rect 317086 158612 317092 158614
rect 317156 158612 317162 158676
rect 319437 158672 319484 158676
rect 319548 158674 319554 158676
rect 319437 158616 319442 158672
rect 319437 158612 319484 158616
rect 319548 158614 319594 158674
rect 320541 158672 320588 158676
rect 320652 158674 320658 158676
rect 320541 158616 320546 158672
rect 319548 158612 319554 158614
rect 320541 158612 320588 158616
rect 320652 158614 320698 158674
rect 323117 158672 323164 158676
rect 323228 158674 323234 158676
rect 323117 158616 323122 158672
rect 320652 158612 320658 158614
rect 323117 158612 323164 158616
rect 323228 158614 323274 158674
rect 324221 158672 324268 158676
rect 324332 158674 324338 158676
rect 324221 158616 324226 158672
rect 323228 158612 323234 158614
rect 324221 158612 324268 158616
rect 324332 158614 324378 158674
rect 326429 158672 326476 158676
rect 326540 158674 326546 158676
rect 326429 158616 326434 158672
rect 324332 158612 324338 158614
rect 326429 158612 326476 158616
rect 326540 158614 326586 158674
rect 328269 158672 328316 158676
rect 328380 158674 328386 158676
rect 328269 158616 328274 158672
rect 326540 158612 326546 158614
rect 328269 158612 328316 158616
rect 328380 158614 328426 158674
rect 328637 158672 328684 158676
rect 328748 158674 328754 158676
rect 328637 158616 328642 158672
rect 328380 158612 328386 158614
rect 328637 158612 328684 158616
rect 328748 158614 328794 158674
rect 329925 158672 329972 158676
rect 330036 158674 330042 158676
rect 330477 158674 330543 158677
rect 330702 158674 330708 158676
rect 329925 158616 329930 158672
rect 328748 158612 328754 158614
rect 329925 158612 329972 158616
rect 330036 158614 330082 158674
rect 330477 158672 330708 158674
rect 330477 158616 330482 158672
rect 330538 158616 330708 158672
rect 330477 158614 330708 158616
rect 330036 158612 330042 158614
rect 319437 158611 319503 158612
rect 320541 158611 320607 158612
rect 323117 158611 323183 158612
rect 324221 158611 324287 158612
rect 326429 158611 326495 158612
rect 328269 158611 328335 158612
rect 328637 158611 328703 158612
rect 329925 158611 329991 158612
rect 330477 158611 330543 158614
rect 330702 158612 330708 158614
rect 330772 158612 330778 158676
rect 332225 158674 332291 158677
rect 333605 158676 333671 158677
rect 334525 158676 334591 158677
rect 332358 158674 332364 158676
rect 332225 158672 332364 158674
rect 332225 158616 332230 158672
rect 332286 158616 332364 158672
rect 332225 158614 332364 158616
rect 332225 158611 332291 158614
rect 332358 158612 332364 158614
rect 332428 158612 332434 158676
rect 333605 158672 333652 158676
rect 333716 158674 333722 158676
rect 333605 158616 333610 158672
rect 333605 158612 333652 158616
rect 333716 158614 333762 158674
rect 334525 158672 334572 158676
rect 334636 158674 334642 158676
rect 335629 158674 335695 158677
rect 335997 158676 336063 158677
rect 335854 158674 335860 158676
rect 334525 158616 334530 158672
rect 333716 158612 333722 158614
rect 334525 158612 334572 158616
rect 334636 158614 334682 158674
rect 335629 158672 335860 158674
rect 335629 158616 335634 158672
rect 335690 158616 335860 158672
rect 335629 158614 335860 158616
rect 334636 158612 334642 158614
rect 333605 158611 333671 158612
rect 334525 158611 334591 158612
rect 335629 158611 335695 158614
rect 335854 158612 335860 158614
rect 335924 158612 335930 158676
rect 335997 158672 336044 158676
rect 336108 158674 336114 158676
rect 336825 158674 336891 158677
rect 338389 158676 338455 158677
rect 336958 158674 336964 158676
rect 335997 158616 336002 158672
rect 335997 158612 336044 158616
rect 336108 158614 336154 158674
rect 336825 158672 336964 158674
rect 336825 158616 336830 158672
rect 336886 158616 336964 158672
rect 336825 158614 336964 158616
rect 336108 158612 336114 158614
rect 335997 158611 336063 158612
rect 336825 158611 336891 158614
rect 336958 158612 336964 158614
rect 337028 158612 337034 158676
rect 338389 158672 338436 158676
rect 338500 158674 338506 158676
rect 338757 158674 338823 158677
rect 340965 158676 341031 158677
rect 343541 158676 343607 158677
rect 349797 158676 349863 158677
rect 339350 158674 339356 158676
rect 338389 158616 338394 158672
rect 338389 158612 338436 158616
rect 338500 158614 338546 158674
rect 338757 158672 339356 158674
rect 338757 158616 338762 158672
rect 338818 158616 339356 158672
rect 338757 158614 339356 158616
rect 338500 158612 338506 158614
rect 338389 158611 338455 158612
rect 338757 158611 338823 158614
rect 339350 158612 339356 158614
rect 339420 158612 339426 158676
rect 340965 158672 341012 158676
rect 341076 158674 341082 158676
rect 340965 158616 340970 158672
rect 340965 158612 341012 158616
rect 341076 158614 341122 158674
rect 343541 158672 343588 158676
rect 343652 158674 343658 158676
rect 343541 158616 343546 158672
rect 341076 158612 341082 158614
rect 343541 158612 343588 158616
rect 343652 158614 343698 158674
rect 349797 158672 349844 158676
rect 349908 158674 349914 158676
rect 355225 158674 355291 158677
rect 356973 158676 357039 158677
rect 360837 158676 360903 158677
rect 363413 158676 363479 158677
rect 368197 158676 368263 158677
rect 371049 158676 371115 158677
rect 373441 158676 373507 158677
rect 376017 158676 376083 158677
rect 378593 158676 378659 158677
rect 380985 158676 381051 158677
rect 383561 158676 383627 158677
rect 385953 158676 386019 158677
rect 388529 158676 388595 158677
rect 355726 158674 355732 158676
rect 349797 158616 349802 158672
rect 343652 158612 343658 158614
rect 349797 158612 349844 158616
rect 349908 158614 349954 158674
rect 355225 158672 355732 158674
rect 355225 158616 355230 158672
rect 355286 158616 355732 158672
rect 355225 158614 355732 158616
rect 349908 158612 349914 158614
rect 340965 158611 341031 158612
rect 343541 158611 343607 158612
rect 349797 158611 349863 158612
rect 355225 158611 355291 158614
rect 355726 158612 355732 158614
rect 355796 158612 355802 158676
rect 356973 158672 357020 158676
rect 357084 158674 357090 158676
rect 356973 158616 356978 158672
rect 356973 158612 357020 158616
rect 357084 158614 357130 158674
rect 360837 158672 360884 158676
rect 360948 158674 360954 158676
rect 360837 158616 360842 158672
rect 357084 158612 357090 158614
rect 360837 158612 360884 158616
rect 360948 158614 360994 158674
rect 363413 158672 363460 158676
rect 363524 158674 363530 158676
rect 363413 158616 363418 158672
rect 360948 158612 360954 158614
rect 363413 158612 363460 158616
rect 363524 158614 363570 158674
rect 368197 158672 368244 158676
rect 368308 158674 368314 158676
rect 370998 158674 371004 158676
rect 368197 158616 368202 158672
rect 363524 158612 363530 158614
rect 368197 158612 368244 158616
rect 368308 158614 368354 158674
rect 370958 158614 371004 158674
rect 371068 158672 371115 158676
rect 373390 158674 373396 158676
rect 371110 158616 371115 158672
rect 368308 158612 368314 158614
rect 370998 158612 371004 158614
rect 371068 158612 371115 158616
rect 373350 158614 373396 158674
rect 373460 158672 373507 158676
rect 375966 158674 375972 158676
rect 373502 158616 373507 158672
rect 373390 158612 373396 158614
rect 373460 158612 373507 158616
rect 375926 158614 375972 158674
rect 376036 158672 376083 158676
rect 378542 158674 378548 158676
rect 376078 158616 376083 158672
rect 375966 158612 375972 158614
rect 376036 158612 376083 158616
rect 378502 158614 378548 158674
rect 378612 158672 378659 158676
rect 380934 158674 380940 158676
rect 378654 158616 378659 158672
rect 378542 158612 378548 158614
rect 378612 158612 378659 158616
rect 380894 158614 380940 158674
rect 381004 158672 381051 158676
rect 383510 158674 383516 158676
rect 381046 158616 381051 158672
rect 380934 158612 380940 158614
rect 381004 158612 381051 158616
rect 383470 158614 383516 158674
rect 383580 158672 383627 158676
rect 385902 158674 385908 158676
rect 383622 158616 383627 158672
rect 383510 158612 383516 158614
rect 383580 158612 383627 158616
rect 385862 158614 385908 158674
rect 385972 158672 386019 158676
rect 388478 158674 388484 158676
rect 386014 158616 386019 158672
rect 385902 158612 385908 158614
rect 385972 158612 386019 158616
rect 388438 158614 388484 158674
rect 388548 158672 388595 158676
rect 388590 158616 388595 158672
rect 388478 158612 388484 158614
rect 388548 158612 388595 158616
rect 391054 158612 391060 158676
rect 391124 158674 391130 158676
rect 391473 158674 391539 158677
rect 393497 158676 393563 158677
rect 395889 158676 395955 158677
rect 398465 158676 398531 158677
rect 393446 158674 393452 158676
rect 391124 158672 391539 158674
rect 391124 158616 391478 158672
rect 391534 158616 391539 158672
rect 391124 158614 391539 158616
rect 393406 158614 393452 158674
rect 393516 158672 393563 158676
rect 395838 158674 395844 158676
rect 393558 158616 393563 158672
rect 391124 158612 391130 158614
rect 356973 158611 357039 158612
rect 360837 158611 360903 158612
rect 363413 158611 363479 158612
rect 368197 158611 368263 158612
rect 371049 158611 371115 158612
rect 373441 158611 373507 158612
rect 376017 158611 376083 158612
rect 378593 158611 378659 158612
rect 380985 158611 381051 158612
rect 383561 158611 383627 158612
rect 385953 158611 386019 158612
rect 388529 158611 388595 158612
rect 391473 158611 391539 158614
rect 393446 158612 393452 158614
rect 393516 158612 393563 158616
rect 395798 158614 395844 158674
rect 395908 158672 395955 158676
rect 398414 158674 398420 158676
rect 395950 158616 395955 158672
rect 395838 158612 395844 158614
rect 395908 158612 395955 158616
rect 398374 158614 398420 158674
rect 398484 158672 398531 158676
rect 398526 158616 398531 158672
rect 398414 158612 398420 158614
rect 398484 158612 398531 158616
rect 400990 158612 400996 158676
rect 401060 158674 401066 158676
rect 401409 158674 401475 158677
rect 401060 158672 401475 158674
rect 401060 158616 401414 158672
rect 401470 158616 401475 158672
rect 401060 158614 401475 158616
rect 401060 158612 401066 158614
rect 393497 158611 393563 158612
rect 395889 158611 395955 158612
rect 398465 158611 398531 158612
rect 401409 158611 401475 158614
rect 403382 158612 403388 158676
rect 403452 158674 403458 158676
rect 403801 158674 403867 158677
rect 403452 158672 403867 158674
rect 403452 158616 403806 158672
rect 403862 158616 403867 158672
rect 403452 158614 403867 158616
rect 403452 158612 403458 158614
rect 403801 158611 403867 158614
rect 405958 158612 405964 158676
rect 406028 158674 406034 158676
rect 406745 158674 406811 158677
rect 406028 158672 406811 158674
rect 406028 158616 406750 158672
rect 406806 158616 406811 158672
rect 406028 158614 406811 158616
rect 406028 158612 406034 158614
rect 406745 158611 406811 158614
rect 135897 158540 135963 158541
rect 137001 158540 137067 158541
rect 135846 158538 135852 158540
rect 135806 158478 135852 158538
rect 135916 158536 135963 158540
rect 136950 158538 136956 158540
rect 135958 158480 135963 158536
rect 135846 158476 135852 158478
rect 135916 158476 135963 158480
rect 136910 158478 136956 158538
rect 137020 158536 137067 158540
rect 137062 158480 137067 158536
rect 136950 158476 136956 158478
rect 137020 158476 137067 158480
rect 138054 158476 138060 158540
rect 138124 158538 138130 158540
rect 139209 158538 139275 158541
rect 138124 158536 139275 158538
rect 138124 158480 139214 158536
rect 139270 158480 139275 158536
rect 138124 158478 139275 158480
rect 138124 158476 138130 158478
rect 135897 158475 135963 158476
rect 137001 158475 137067 158476
rect 139209 158475 139275 158478
rect 139526 158476 139532 158540
rect 139596 158538 139602 158540
rect 140681 158538 140747 158541
rect 139596 158536 140747 158538
rect 139596 158480 140686 158536
rect 140742 158480 140747 158536
rect 139596 158478 140747 158480
rect 139596 158476 139602 158478
rect 140681 158475 140747 158478
rect 175958 158476 175964 158540
rect 176028 158538 176034 158540
rect 282361 158538 282427 158541
rect 176028 158536 282427 158538
rect 176028 158480 282366 158536
rect 282422 158480 282427 158536
rect 176028 158478 282427 158480
rect 176028 158476 176034 158478
rect 282361 158475 282427 158478
rect 284661 158538 284727 158541
rect 284845 158538 284911 158541
rect 359222 158538 359228 158540
rect 284661 158536 359228 158538
rect 284661 158480 284666 158536
rect 284722 158480 284850 158536
rect 284906 158480 359228 158536
rect 284661 158478 359228 158480
rect 284661 158475 284727 158478
rect 284845 158475 284911 158478
rect 359222 158476 359228 158478
rect 359292 158476 359298 158540
rect 149830 158340 149836 158404
rect 149900 158402 149906 158404
rect 150249 158402 150315 158405
rect 149900 158400 150315 158402
rect 149900 158344 150254 158400
rect 150310 158344 150315 158400
rect 149900 158342 150315 158344
rect 149900 158340 149906 158342
rect 150249 158339 150315 158342
rect 178534 158340 178540 158404
rect 178604 158402 178610 158404
rect 178953 158402 179019 158405
rect 178604 158400 179019 158402
rect 178604 158344 178958 158400
rect 179014 158344 179019 158400
rect 178604 158342 179019 158344
rect 178604 158340 178610 158342
rect 178953 158339 179019 158342
rect 180926 158340 180932 158404
rect 180996 158402 181002 158404
rect 181713 158402 181779 158405
rect 195881 158404 195947 158405
rect 198457 158404 198523 158405
rect 195830 158402 195836 158404
rect 180996 158400 181779 158402
rect 180996 158344 181718 158400
rect 181774 158344 181779 158400
rect 180996 158342 181779 158344
rect 195790 158342 195836 158402
rect 195900 158400 195947 158404
rect 198406 158402 198412 158404
rect 195942 158344 195947 158400
rect 180996 158340 181002 158342
rect 181713 158339 181779 158342
rect 195830 158340 195836 158342
rect 195900 158340 195947 158344
rect 198366 158342 198412 158402
rect 198476 158400 198523 158404
rect 198518 158344 198523 158400
rect 198406 158340 198412 158342
rect 198476 158340 198523 158344
rect 195881 158339 195947 158340
rect 198457 158339 198523 158340
rect 276013 158402 276079 158405
rect 277301 158402 277367 158405
rect 338113 158404 338179 158405
rect 331254 158402 331260 158404
rect 276013 158400 331260 158402
rect 276013 158344 276018 158400
rect 276074 158344 277306 158400
rect 277362 158344 331260 158400
rect 276013 158342 331260 158344
rect 276013 158339 276079 158342
rect 277301 158339 277367 158342
rect 331254 158340 331260 158342
rect 331324 158340 331330 158404
rect 338062 158402 338068 158404
rect 338022 158342 338068 158402
rect 338132 158400 338179 158404
rect 338174 158344 338179 158400
rect 338062 158340 338068 158342
rect 338132 158340 338179 158344
rect 338113 158339 338179 158340
rect 117078 158204 117084 158268
rect 117148 158266 117154 158268
rect 117221 158266 117287 158269
rect 117148 158264 117287 158266
rect 117148 158208 117226 158264
rect 117282 158208 117287 158264
rect 117148 158206 117287 158208
rect 117148 158204 117154 158206
rect 117221 158203 117287 158206
rect 141182 158204 141188 158268
rect 141252 158266 141258 158268
rect 141417 158266 141483 158269
rect 141785 158268 141851 158269
rect 146017 158268 146083 158269
rect 146385 158268 146451 158269
rect 150985 158268 151051 158269
rect 141734 158266 141740 158268
rect 141252 158264 141483 158266
rect 141252 158208 141422 158264
rect 141478 158208 141483 158264
rect 141252 158206 141483 158208
rect 141694 158206 141740 158266
rect 141804 158264 141851 158268
rect 145966 158266 145972 158268
rect 141846 158208 141851 158264
rect 141252 158204 141258 158206
rect 141417 158203 141483 158206
rect 141734 158204 141740 158206
rect 141804 158204 141851 158208
rect 145926 158206 145972 158266
rect 146036 158264 146083 158268
rect 146334 158266 146340 158268
rect 146078 158208 146083 158264
rect 145966 158204 145972 158206
rect 146036 158204 146083 158208
rect 146294 158206 146340 158266
rect 146404 158264 146451 158268
rect 150934 158266 150940 158268
rect 146446 158208 146451 158264
rect 146334 158204 146340 158206
rect 146404 158204 146451 158208
rect 150894 158206 150940 158266
rect 151004 158264 151051 158268
rect 151046 158208 151051 158264
rect 150934 158204 150940 158206
rect 151004 158204 151051 158208
rect 170990 158204 170996 158268
rect 171060 158266 171066 158268
rect 238201 158266 238267 158269
rect 171060 158264 238267 158266
rect 171060 158208 238206 158264
rect 238262 158208 238267 158264
rect 171060 158206 238267 158208
rect 171060 158204 171066 158206
rect 141785 158203 141851 158204
rect 146017 158203 146083 158204
rect 146385 158203 146451 158204
rect 150985 158203 151051 158204
rect 238201 158203 238267 158206
rect 274633 158266 274699 158269
rect 275921 158266 275987 158269
rect 343909 158268 343975 158269
rect 348693 158268 348759 158269
rect 353293 158268 353359 158269
rect 327574 158266 327580 158268
rect 274633 158264 327580 158266
rect 274633 158208 274638 158264
rect 274694 158208 275926 158264
rect 275982 158208 327580 158264
rect 274633 158206 327580 158208
rect 274633 158203 274699 158206
rect 275921 158203 275987 158206
rect 327574 158204 327580 158206
rect 327644 158204 327650 158268
rect 343909 158264 343956 158268
rect 344020 158266 344026 158268
rect 343909 158208 343914 158264
rect 343909 158204 343956 158208
rect 344020 158206 344066 158266
rect 348693 158264 348740 158268
rect 348804 158266 348810 158268
rect 348693 158208 348698 158264
rect 344020 158204 344026 158206
rect 348693 158204 348740 158208
rect 348804 158206 348850 158266
rect 353293 158264 353340 158268
rect 353404 158266 353410 158268
rect 353293 158208 353298 158264
rect 348804 158204 348810 158206
rect 353293 158204 353340 158208
rect 353404 158206 353450 158266
rect 353404 158204 353410 158206
rect 343909 158203 343975 158204
rect 348693 158203 348759 158204
rect 353293 158203 353359 158204
rect 185945 158132 186011 158133
rect 185894 158130 185900 158132
rect 185854 158070 185900 158130
rect 185964 158128 186011 158132
rect 186006 158072 186011 158128
rect 185894 158068 185900 158070
rect 185964 158068 186011 158072
rect 188654 158068 188660 158132
rect 188724 158130 188730 158132
rect 238385 158130 238451 158133
rect 188724 158128 238451 158130
rect 188724 158072 238390 158128
rect 238446 158072 238451 158128
rect 188724 158070 238451 158072
rect 188724 158068 188730 158070
rect 185945 158067 186011 158068
rect 238385 158067 238451 158070
rect 284569 158130 284635 158133
rect 285305 158130 285371 158133
rect 333462 158130 333468 158132
rect 284569 158128 333468 158130
rect 284569 158072 284574 158128
rect 284630 158072 285310 158128
rect 285366 158072 333468 158128
rect 284569 158070 333468 158072
rect 284569 158067 284635 158070
rect 285305 158067 285371 158070
rect 333462 158068 333468 158070
rect 333532 158068 333538 158132
rect 125409 157996 125475 157997
rect 125358 157994 125364 157996
rect 125318 157934 125364 157994
rect 125428 157992 125475 157996
rect 125470 157936 125475 157992
rect 125358 157932 125364 157934
rect 125428 157932 125475 157936
rect 125409 157931 125475 157932
rect 140589 157996 140655 157997
rect 140589 157992 140636 157996
rect 140700 157994 140706 157996
rect 289629 157994 289695 157997
rect 322054 157994 322060 157996
rect 140589 157936 140594 157992
rect 140589 157932 140636 157936
rect 140700 157934 140746 157994
rect 289629 157992 322060 157994
rect 289629 157936 289634 157992
rect 289690 157936 322060 157992
rect 289629 157934 322060 157936
rect 140700 157932 140706 157934
rect 140589 157931 140655 157932
rect 289629 157931 289695 157934
rect 322054 157932 322060 157934
rect 322124 157932 322130 157996
rect 325141 157994 325207 157997
rect 346393 157996 346459 157997
rect 325366 157994 325372 157996
rect 325141 157992 325372 157994
rect 325141 157936 325146 157992
rect 325202 157936 325372 157992
rect 325141 157934 325372 157936
rect 325141 157931 325207 157934
rect 325366 157932 325372 157934
rect 325436 157932 325442 157996
rect 346342 157994 346348 157996
rect 346302 157934 346348 157994
rect 346412 157992 346459 157996
rect 346454 157936 346459 157992
rect 346342 157932 346348 157934
rect 346412 157932 346459 157936
rect 346393 157931 346459 157932
rect 143942 157796 143948 157860
rect 144012 157858 144018 157860
rect 144269 157858 144335 157861
rect 145281 157860 145347 157861
rect 148777 157860 148843 157861
rect 145230 157858 145236 157860
rect 144012 157856 144335 157858
rect 144012 157800 144274 157856
rect 144330 157800 144335 157856
rect 144012 157798 144335 157800
rect 145190 157798 145236 157858
rect 145300 157856 145347 157860
rect 148726 157858 148732 157860
rect 145342 157800 145347 157856
rect 144012 157796 144018 157798
rect 144269 157795 144335 157798
rect 145230 157796 145236 157798
rect 145300 157796 145347 157800
rect 148686 157798 148732 157858
rect 148796 157856 148843 157860
rect 148838 157800 148843 157856
rect 148726 157796 148732 157798
rect 148796 157796 148843 157800
rect 193438 157796 193444 157860
rect 193508 157858 193514 157860
rect 193949 157858 194015 157861
rect 193508 157856 194015 157858
rect 193508 157800 193954 157856
rect 194010 157800 194015 157856
rect 193508 157798 194015 157800
rect 193508 157796 193514 157798
rect 145281 157795 145347 157796
rect 148777 157795 148843 157796
rect 193949 157795 194015 157798
rect 339493 157858 339559 157861
rect 340638 157858 340644 157860
rect 339493 157856 340644 157858
rect 339493 157800 339498 157856
rect 339554 157800 340644 157856
rect 339493 157798 340644 157800
rect 339493 157795 339559 157798
rect 340638 157796 340644 157798
rect 340708 157796 340714 157860
rect 341149 157858 341215 157861
rect 342805 157860 342871 157861
rect 341742 157858 341748 157860
rect 341149 157856 341748 157858
rect 341149 157800 341154 157856
rect 341210 157800 341748 157856
rect 341149 157798 341748 157800
rect 341149 157795 341215 157798
rect 341742 157796 341748 157798
rect 341812 157796 341818 157860
rect 342805 157856 342852 157860
rect 342916 157858 342922 157860
rect 345105 157858 345171 157861
rect 345238 157858 345244 157860
rect 342805 157800 342810 157856
rect 342805 157796 342852 157800
rect 342916 157798 342962 157858
rect 345105 157856 345244 157858
rect 345105 157800 345110 157856
rect 345166 157800 345244 157856
rect 345105 157798 345244 157800
rect 342916 157796 342922 157798
rect 342805 157795 342871 157796
rect 345105 157795 345171 157798
rect 345238 157796 345244 157798
rect 345308 157796 345314 157860
rect 346853 157858 346919 157861
rect 347630 157858 347636 157860
rect 346853 157856 347636 157858
rect 346853 157800 346858 157856
rect 346914 157800 347636 157856
rect 346853 157798 347636 157800
rect 346853 157795 346919 157798
rect 347630 157796 347636 157798
rect 347700 157796 347706 157860
rect 130694 157660 130700 157724
rect 130764 157722 130770 157724
rect 282494 157722 282500 157724
rect 130764 157662 282500 157722
rect 130764 157660 130770 157662
rect 282494 157660 282500 157662
rect 282564 157660 282570 157724
rect 142838 157524 142844 157588
rect 142908 157586 142914 157588
rect 143073 157586 143139 157589
rect 142908 157584 143139 157586
rect 142908 157528 143078 157584
rect 143134 157528 143139 157584
rect 142908 157526 143139 157528
rect 142908 157524 142914 157526
rect 143073 157523 143139 157526
rect 147622 157524 147628 157588
rect 147692 157586 147698 157588
rect 147765 157586 147831 157589
rect 201033 157588 201099 157589
rect 200982 157586 200988 157588
rect 147692 157584 147831 157586
rect 147692 157528 147770 157584
rect 147826 157528 147831 157584
rect 147692 157526 147831 157528
rect 200942 157526 200988 157586
rect 201052 157584 201099 157588
rect 201094 157528 201099 157584
rect 147692 157524 147698 157526
rect 147765 157523 147831 157526
rect 200982 157524 200988 157526
rect 201052 157524 201099 157528
rect 205950 157524 205956 157588
rect 206020 157586 206026 157588
rect 206277 157586 206343 157589
rect 206020 157584 206343 157586
rect 206020 157528 206282 157584
rect 206338 157528 206343 157584
rect 206020 157526 206343 157528
rect 206020 157524 206026 157526
rect 201033 157523 201099 157524
rect 206277 157523 206343 157526
rect 278681 157586 278747 157589
rect 358118 157586 358124 157588
rect 278681 157584 358124 157586
rect 278681 157528 278686 157584
rect 278742 157528 358124 157584
rect 278681 157526 358124 157528
rect 278681 157523 278747 157526
rect 358118 157524 358124 157526
rect 358188 157524 358194 157588
rect 118233 157452 118299 157453
rect 136081 157452 136147 157453
rect 118182 157450 118188 157452
rect 118142 157390 118188 157450
rect 118252 157448 118299 157452
rect 118294 157392 118299 157448
rect 118182 157388 118188 157390
rect 118252 157388 118299 157392
rect 133638 157388 133644 157452
rect 133708 157388 133714 157452
rect 136030 157450 136036 157452
rect 135990 157390 136036 157450
rect 136100 157448 136147 157452
rect 136142 157392 136147 157448
rect 136030 157388 136036 157390
rect 136100 157388 136147 157392
rect 138606 157388 138612 157452
rect 138676 157450 138682 157452
rect 138933 157450 138999 157453
rect 138676 157448 138999 157450
rect 138676 157392 138938 157448
rect 138994 157392 138999 157448
rect 138676 157390 138999 157392
rect 138676 157388 138682 157390
rect 118233 157387 118299 157388
rect 133646 157314 133706 157388
rect 136081 157387 136147 157388
rect 138933 157387 138999 157390
rect 143574 157388 143580 157452
rect 143644 157450 143650 157452
rect 144361 157450 144427 157453
rect 148409 157452 148475 157453
rect 151353 157452 151419 157453
rect 148358 157450 148364 157452
rect 143644 157448 144427 157450
rect 143644 157392 144366 157448
rect 144422 157392 144427 157448
rect 143644 157390 144427 157392
rect 148318 157390 148364 157450
rect 148428 157448 148475 157452
rect 151302 157450 151308 157452
rect 148470 157392 148475 157448
rect 143644 157388 143650 157390
rect 144361 157387 144427 157390
rect 148358 157388 148364 157390
rect 148428 157388 148475 157392
rect 151262 157390 151308 157450
rect 151372 157448 151419 157452
rect 151414 157392 151419 157448
rect 151302 157388 151308 157390
rect 151372 157388 151419 157392
rect 152222 157388 152228 157452
rect 152292 157450 152298 157452
rect 152641 157450 152707 157453
rect 152292 157448 152707 157450
rect 152292 157392 152646 157448
rect 152702 157392 152707 157448
rect 152292 157390 152707 157392
rect 152292 157388 152298 157390
rect 148409 157387 148475 157388
rect 151353 157387 151419 157388
rect 152641 157387 152707 157390
rect 153326 157388 153332 157452
rect 153396 157450 153402 157452
rect 153929 157450 153995 157453
rect 154481 157452 154547 157453
rect 155769 157452 155835 157453
rect 157057 157452 157123 157453
rect 154430 157450 154436 157452
rect 153396 157448 153995 157450
rect 153396 157392 153934 157448
rect 153990 157392 153995 157448
rect 153396 157390 153995 157392
rect 154390 157390 154436 157450
rect 154500 157448 154547 157452
rect 155718 157450 155724 157452
rect 154542 157392 154547 157448
rect 153396 157388 153402 157390
rect 153929 157387 153995 157390
rect 154430 157388 154436 157390
rect 154500 157388 154547 157392
rect 155678 157390 155724 157450
rect 155788 157448 155835 157452
rect 157006 157450 157012 157452
rect 155830 157392 155835 157448
rect 155718 157388 155724 157390
rect 155788 157388 155835 157392
rect 156966 157390 157012 157450
rect 157076 157448 157123 157452
rect 157118 157392 157123 157448
rect 157006 157388 157012 157390
rect 157076 157388 157123 157392
rect 183502 157388 183508 157452
rect 183572 157450 183578 157452
rect 279366 157450 279372 157452
rect 183572 157390 279372 157450
rect 183572 157388 183578 157390
rect 279366 157388 279372 157390
rect 279436 157388 279442 157452
rect 317689 157450 317755 157453
rect 351085 157452 351151 157453
rect 352189 157452 352255 157453
rect 354397 157452 354463 157453
rect 318190 157450 318196 157452
rect 317689 157448 318196 157450
rect 317689 157392 317694 157448
rect 317750 157392 318196 157448
rect 317689 157390 318196 157392
rect 154481 157387 154547 157388
rect 155769 157387 155835 157388
rect 157057 157387 157123 157388
rect 317689 157387 317755 157390
rect 318190 157388 318196 157390
rect 318260 157388 318266 157452
rect 351085 157448 351132 157452
rect 351196 157450 351202 157452
rect 351085 157392 351090 157448
rect 351085 157388 351132 157392
rect 351196 157390 351242 157450
rect 352189 157448 352236 157452
rect 352300 157450 352306 157452
rect 352189 157392 352194 157448
rect 351196 157388 351202 157390
rect 352189 157388 352236 157392
rect 352300 157390 352346 157450
rect 354397 157448 354444 157452
rect 354508 157450 354514 157452
rect 354397 157392 354402 157448
rect 352300 157388 352306 157390
rect 354397 157388 354444 157392
rect 354508 157390 354554 157450
rect 354508 157388 354514 157390
rect 351085 157387 351151 157388
rect 352189 157387 352255 157388
rect 354397 157387 354463 157388
rect 273989 157314 274055 157317
rect 133646 157312 274055 157314
rect 133646 157256 273994 157312
rect 274050 157256 274055 157312
rect 133646 157254 274055 157256
rect 273989 157251 274055 157254
rect 202873 156906 202939 156909
rect 266813 156906 266879 156909
rect 202873 156904 266879 156906
rect 202873 156848 202878 156904
rect 202934 156848 266818 156904
rect 266874 156848 266879 156904
rect 202873 156846 266879 156848
rect 202873 156843 202939 156846
rect 266813 156843 266879 156846
rect 178033 156770 178099 156773
rect 255957 156770 256023 156773
rect 178033 156768 256023 156770
rect 178033 156712 178038 156768
rect 178094 156712 255962 156768
rect 256018 156712 256023 156768
rect 178033 156710 256023 156712
rect 178033 156707 178099 156710
rect 255957 156707 256023 156710
rect 125593 156634 125659 156637
rect 252829 156634 252895 156637
rect 125593 156632 252895 156634
rect 125593 156576 125598 156632
rect 125654 156576 252834 156632
rect 252890 156576 252895 156632
rect 125593 156574 252895 156576
rect 125593 156571 125659 156574
rect 252829 156571 252895 156574
rect 185945 155954 186011 155957
rect 279550 155954 279556 155956
rect 185945 155952 279556 155954
rect 185945 155896 185950 155952
rect 186006 155896 279556 155952
rect 185945 155894 279556 155896
rect 185945 155891 186011 155894
rect 279550 155892 279556 155894
rect 279620 155892 279626 155956
rect 220813 155546 220879 155549
rect 270953 155546 271019 155549
rect 220813 155544 271019 155546
rect 220813 155488 220818 155544
rect 220874 155488 270958 155544
rect 271014 155488 271019 155544
rect 220813 155486 271019 155488
rect 220813 155483 220879 155486
rect 270953 155483 271019 155486
rect 182173 155410 182239 155413
rect 262489 155410 262555 155413
rect 182173 155408 262555 155410
rect 182173 155352 182178 155408
rect 182234 155352 262494 155408
rect 262550 155352 262555 155408
rect 182173 155350 262555 155352
rect 182173 155347 182239 155350
rect 262489 155347 262555 155350
rect 160093 155274 160159 155277
rect 259913 155274 259979 155277
rect 160093 155272 259979 155274
rect 160093 155216 160098 155272
rect 160154 155216 259918 155272
rect 259974 155216 259979 155272
rect 160093 155214 259979 155216
rect 160093 155211 160159 155214
rect 259913 155211 259979 155214
rect 286726 153716 286732 153780
rect 286796 153778 286802 153780
rect 309133 153778 309199 153781
rect 286796 153776 309199 153778
rect 286796 153720 309138 153776
rect 309194 153720 309199 153776
rect 286796 153718 309199 153720
rect 286796 153716 286802 153718
rect 309133 153715 309199 153718
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect 284886 150996 284892 151060
rect 284956 151058 284962 151060
rect 300853 151058 300919 151061
rect 284956 151056 300919 151058
rect 284956 151000 300858 151056
rect 300914 151000 300919 151056
rect 284956 150998 300919 151000
rect 284956 150996 284962 150998
rect 300853 150995 300919 150998
rect 269757 150378 269823 150381
rect 277158 150378 277164 150380
rect 269757 150376 277164 150378
rect 269757 150320 269762 150376
rect 269818 150320 277164 150376
rect 269757 150318 277164 150320
rect 269757 150315 269823 150318
rect 277158 150316 277164 150318
rect 277228 150316 277234 150380
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3141 136778 3207 136781
rect -960 136776 3207 136778
rect -960 136720 3146 136776
rect 3202 136720 3207 136776
rect -960 136718 3207 136720
rect -960 136628 480 136718
rect 3141 136715 3207 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3693 97610 3759 97613
rect -960 97608 3759 97610
rect -960 97552 3698 97608
rect 3754 97552 3759 97608
rect -960 97550 3759 97552
rect -960 97460 480 97550
rect 3693 97547 3759 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 298318 75108 298324 75172
rect 298388 75170 298394 75172
rect 375373 75170 375439 75173
rect 298388 75168 375439 75170
rect 298388 75112 375378 75168
rect 375434 75112 375439 75168
rect 298388 75110 375439 75112
rect 298388 75108 298394 75110
rect 375373 75107 375439 75110
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 439446 71844 439452 71908
rect 439516 71906 439522 71908
rect 583526 71906 583586 72798
rect 439516 71846 583586 71906
rect 439516 71844 439522 71846
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 283966 9556 283972 9620
rect 284036 9618 284042 9620
rect 374085 9618 374151 9621
rect 284036 9616 374151 9618
rect 284036 9560 374090 9616
rect 374146 9560 374151 9616
rect 284036 9558 374151 9560
rect 284036 9556 284042 9558
rect 374085 9555 374151 9558
rect 293350 9420 293356 9484
rect 293420 9482 293426 9484
rect 387149 9482 387215 9485
rect 293420 9480 387215 9482
rect 293420 9424 387154 9480
rect 387210 9424 387215 9480
rect 293420 9422 387215 9424
rect 293420 9420 293426 9422
rect 387149 9419 387215 9422
rect 289302 9284 289308 9348
rect 289372 9346 289378 9348
rect 394233 9346 394299 9349
rect 289372 9344 394299 9346
rect 289372 9288 394238 9344
rect 394294 9288 394299 9344
rect 289372 9286 394299 9288
rect 289372 9284 289378 9286
rect 394233 9283 394299 9286
rect 295190 9148 295196 9212
rect 295260 9210 295266 9212
rect 408401 9210 408467 9213
rect 295260 9208 408467 9210
rect 295260 9152 408406 9208
rect 408462 9152 408467 9208
rect 295260 9150 408467 9152
rect 295260 9148 295266 9150
rect 408401 9147 408467 9150
rect 285070 9012 285076 9076
rect 285140 9074 285146 9076
rect 397729 9074 397795 9077
rect 285140 9072 397795 9074
rect 285140 9016 397734 9072
rect 397790 9016 397795 9072
rect 285140 9014 397795 9016
rect 285140 9012 285146 9014
rect 397729 9011 397795 9014
rect 286910 8876 286916 8940
rect 286980 8938 286986 8940
rect 404813 8938 404879 8941
rect 286980 8936 404879 8938
rect 286980 8880 404818 8936
rect 404874 8880 404879 8936
rect 286980 8878 404879 8880
rect 286980 8876 286986 8878
rect 404813 8875 404879 8878
rect 289486 8740 289492 8804
rect 289556 8802 289562 8804
rect 379973 8802 380039 8805
rect 289556 8800 380039 8802
rect 289556 8744 379978 8800
rect 380034 8744 380039 8800
rect 289556 8742 380039 8744
rect 289556 8740 289562 8742
rect 379973 8739 380039 8742
rect 298502 6836 298508 6900
rect 298572 6898 298578 6900
rect 372889 6898 372955 6901
rect 298572 6896 372955 6898
rect 298572 6840 372894 6896
rect 372950 6840 372955 6896
rect 298572 6838 372955 6840
rect 298572 6836 298578 6838
rect 372889 6835 372955 6838
rect 292430 6700 292436 6764
rect 292500 6762 292506 6764
rect 382365 6762 382431 6765
rect 292500 6760 382431 6762
rect 292500 6704 382370 6760
rect 382426 6704 382431 6760
rect 292500 6702 382431 6704
rect 292500 6700 292506 6702
rect 382365 6699 382431 6702
rect -960 6490 480 6580
rect 292246 6564 292252 6628
rect 292316 6626 292322 6628
rect 389449 6626 389515 6629
rect 292316 6624 389515 6626
rect 292316 6568 389454 6624
rect 389510 6568 389515 6624
rect 292316 6566 389515 6568
rect 292316 6564 292322 6566
rect 389449 6563 389515 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 290958 6428 290964 6492
rect 291028 6490 291034 6492
rect 393037 6490 393103 6493
rect 291028 6488 393103 6490
rect 291028 6432 393042 6488
rect 393098 6432 393103 6488
rect 583520 6476 584960 6716
rect 291028 6430 393103 6432
rect 291028 6428 291034 6430
rect 393037 6427 393103 6430
rect 288198 6292 288204 6356
rect 288268 6354 288274 6356
rect 390645 6354 390711 6357
rect 288268 6352 390711 6354
rect 288268 6296 390650 6352
rect 390706 6296 390711 6352
rect 288268 6294 390711 6296
rect 288268 6292 288274 6294
rect 390645 6291 390711 6294
rect 292062 6156 292068 6220
rect 292132 6218 292138 6220
rect 396533 6218 396599 6221
rect 292132 6216 396599 6218
rect 292132 6160 396538 6216
rect 396594 6160 396599 6216
rect 292132 6158 396599 6160
rect 292132 6156 292138 6158
rect 396533 6155 396599 6158
rect 297582 6020 297588 6084
rect 297652 6082 297658 6084
rect 369393 6082 369459 6085
rect 297652 6080 369459 6082
rect 297652 6024 369398 6080
rect 369454 6024 369459 6080
rect 297652 6022 369459 6024
rect 297652 6020 297658 6022
rect 369393 6019 369459 6022
rect 297950 4932 297956 4996
rect 298020 4994 298026 4996
rect 368197 4994 368263 4997
rect 298020 4992 368263 4994
rect 298020 4936 368202 4992
rect 368258 4936 368263 4992
rect 298020 4934 368263 4936
rect 298020 4932 298026 4934
rect 368197 4931 368263 4934
rect 297766 4796 297772 4860
rect 297836 4858 297842 4860
rect 370589 4858 370655 4861
rect 297836 4856 370655 4858
rect 297836 4800 370594 4856
rect 370650 4800 370655 4856
rect 297836 4798 370655 4800
rect 297836 4796 297842 4798
rect 370589 4795 370655 4798
rect 295926 3980 295932 4044
rect 295996 4042 296002 4044
rect 381169 4042 381235 4045
rect 295996 4040 381235 4042
rect 295996 3984 381174 4040
rect 381230 3984 381235 4040
rect 295996 3982 381235 3984
rect 295996 3980 296002 3982
rect 381169 3979 381235 3982
rect 296110 3844 296116 3908
rect 296180 3906 296186 3908
rect 383561 3906 383627 3909
rect 296180 3904 383627 3906
rect 296180 3848 383566 3904
rect 383622 3848 383627 3904
rect 296180 3846 383627 3848
rect 296180 3844 296186 3846
rect 383561 3843 383627 3846
rect 296478 3708 296484 3772
rect 296548 3770 296554 3772
rect 388253 3770 388319 3773
rect 296548 3768 388319 3770
rect 296548 3712 388258 3768
rect 388314 3712 388319 3768
rect 296548 3710 388319 3712
rect 296548 3708 296554 3710
rect 388253 3707 388319 3710
rect 435541 3770 435607 3773
rect 439262 3770 439268 3772
rect 435541 3768 439268 3770
rect 435541 3712 435546 3768
rect 435602 3712 439268 3768
rect 435541 3710 439268 3712
rect 435541 3707 435607 3710
rect 439262 3708 439268 3710
rect 439332 3708 439338 3772
rect 296294 3572 296300 3636
rect 296364 3634 296370 3636
rect 391841 3634 391907 3637
rect 296364 3632 391907 3634
rect 296364 3576 391846 3632
rect 391902 3576 391907 3632
rect 296364 3574 391907 3576
rect 296364 3572 296370 3574
rect 391841 3571 391907 3574
rect 433241 3634 433307 3637
rect 437606 3634 437612 3636
rect 433241 3632 437612 3634
rect 433241 3576 433246 3632
rect 433302 3576 437612 3632
rect 433241 3574 437612 3576
rect 433241 3571 433307 3574
rect 437606 3572 437612 3574
rect 437676 3572 437682 3636
rect 293534 3436 293540 3500
rect 293604 3498 293610 3500
rect 395337 3498 395403 3501
rect 293604 3496 395403 3498
rect 293604 3440 395342 3496
rect 395398 3440 395403 3496
rect 293604 3438 395403 3440
rect 293604 3436 293610 3438
rect 395337 3435 395403 3438
rect 437422 3436 437428 3500
rect 437492 3498 437498 3500
rect 437933 3498 437999 3501
rect 439129 3500 439195 3501
rect 437492 3496 437999 3498
rect 437492 3440 437938 3496
rect 437994 3440 437999 3496
rect 437492 3438 437999 3440
rect 437492 3436 437498 3438
rect 437933 3435 437999 3438
rect 439078 3436 439084 3500
rect 439148 3498 439195 3500
rect 439148 3496 439240 3498
rect 439190 3440 439240 3496
rect 439148 3438 439240 3440
rect 439148 3436 439195 3438
rect 439129 3435 439195 3436
rect 293718 3300 293724 3364
rect 293788 3362 293794 3364
rect 398925 3362 398991 3365
rect 293788 3360 398991 3362
rect 293788 3304 398930 3360
rect 398986 3304 398991 3360
rect 293788 3302 398991 3304
rect 293788 3300 293794 3302
rect 398925 3299 398991 3302
rect 432045 3362 432111 3365
rect 437790 3362 437796 3364
rect 432045 3360 437796 3362
rect 432045 3304 432050 3360
rect 432106 3304 437796 3360
rect 432045 3302 437796 3304
rect 432045 3299 432111 3302
rect 437790 3300 437796 3302
rect 437860 3300 437866 3364
rect 284150 3164 284156 3228
rect 284220 3226 284226 3228
rect 363505 3226 363571 3229
rect 284220 3224 363571 3226
rect 284220 3168 363510 3224
rect 363566 3168 363571 3224
rect 284220 3166 363571 3168
rect 284220 3164 284226 3166
rect 363505 3163 363571 3166
<< via3 >>
rect 247540 477396 247604 477460
rect 250116 477396 250180 477460
rect 251404 477396 251468 477460
rect 253428 477396 253492 477460
rect 268332 477260 268396 477324
rect 243124 476988 243188 477052
rect 248644 476988 248708 477052
rect 256188 476988 256252 477052
rect 258028 477048 258092 477052
rect 258028 476992 258078 477048
rect 258078 476992 258092 477048
rect 258028 476988 258092 476992
rect 270908 476988 270972 477052
rect 305868 476988 305932 477052
rect 308444 476988 308508 477052
rect 245332 476852 245396 476916
rect 303476 476852 303540 476916
rect 311020 476852 311084 476916
rect 323348 476852 323412 476916
rect 325924 476852 325988 476916
rect 257108 476716 257172 476780
rect 258396 476716 258460 476780
rect 248276 476580 248340 476644
rect 253612 476580 253676 476644
rect 260972 476580 261036 476644
rect 263548 476640 263612 476644
rect 263548 476584 263598 476640
rect 263598 476584 263612 476640
rect 263548 476580 263612 476584
rect 265940 476580 266004 476644
rect 278452 476580 278516 476644
rect 239628 476444 239692 476508
rect 244412 476444 244476 476508
rect 250668 476444 250732 476508
rect 262812 476444 262876 476508
rect 273484 476444 273548 476508
rect 313412 476444 313476 476508
rect 315804 476444 315868 476508
rect 235948 476368 236012 476372
rect 235948 476312 235998 476368
rect 235998 476312 236012 476368
rect 235948 476308 236012 476312
rect 254532 476308 254596 476372
rect 260788 476308 260852 476372
rect 263916 476308 263980 476372
rect 267596 476368 267660 476372
rect 267596 476312 267610 476368
rect 267610 476312 267660 476368
rect 267596 476308 267660 476312
rect 273300 476308 273364 476372
rect 276060 476368 276124 476372
rect 276060 476312 276074 476368
rect 276074 476312 276124 476368
rect 276060 476308 276124 476312
rect 318380 476308 318444 476372
rect 320956 476308 321020 476372
rect 237052 476172 237116 476236
rect 238156 476172 238220 476236
rect 240548 476172 240612 476236
rect 241836 476172 241900 476236
rect 246436 476172 246500 476236
rect 252324 476232 252388 476236
rect 252324 476176 252374 476232
rect 252374 476176 252388 476232
rect 252324 476172 252388 476176
rect 255820 476172 255884 476236
rect 259500 476172 259564 476236
rect 261708 476172 261772 476236
rect 265388 476172 265452 476236
rect 266492 476172 266556 476236
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 274404 476172 274468 476236
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278084 476172 278148 476236
rect 279188 476172 279252 476236
rect 280844 476172 280908 476236
rect 283420 476172 283484 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293356 476172 293420 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476232 300964 476236
rect 300900 476176 300914 476232
rect 300914 476176 300964 476232
rect 300900 476172 300964 476176
rect 439452 442988 439516 443052
rect 358860 442716 358924 442780
rect 295196 309028 295260 309092
rect 296300 308892 296364 308956
rect 282132 308756 282196 308820
rect 286180 308620 286244 308684
rect 296484 308212 296548 308276
rect 297956 308076 298020 308140
rect 277348 307940 277412 308004
rect 297772 307940 297836 308004
rect 298140 307940 298204 308004
rect 277532 307804 277596 307868
rect 284892 307804 284956 307868
rect 286732 307804 286796 307868
rect 297404 307804 297468 307868
rect 297588 307804 297652 307868
rect 298508 307864 298572 307868
rect 298508 307808 298522 307864
rect 298522 307808 298572 307864
rect 298508 307804 298572 307808
rect 282500 306308 282564 306372
rect 279372 306172 279436 306236
rect 279556 303316 279620 303380
rect 439084 287676 439148 287740
rect 437428 275164 437492 275228
rect 293356 248236 293420 248300
rect 289492 248100 289556 248164
rect 288204 247964 288268 248028
rect 289308 247828 289372 247892
rect 288020 247692 288084 247756
rect 285076 247556 285140 247620
rect 437612 247556 437676 247620
rect 296116 247420 296180 247484
rect 284524 247148 284588 247212
rect 287652 247148 287716 247212
rect 288940 247148 289004 247212
rect 284708 247072 284772 247076
rect 284708 247016 284758 247072
rect 284758 247016 284772 247072
rect 284708 247012 284772 247016
rect 286364 247012 286428 247076
rect 286916 247072 286980 247076
rect 286916 247016 286966 247072
rect 286966 247016 286980 247072
rect 286916 247012 286980 247016
rect 287836 247072 287900 247076
rect 287836 247016 287886 247072
rect 287886 247016 287900 247072
rect 287836 247012 287900 247016
rect 289124 247072 289188 247076
rect 289124 247016 289174 247072
rect 289174 247016 289188 247072
rect 289124 247012 289188 247016
rect 358860 245516 358924 245580
rect 293540 245244 293604 245308
rect 290964 245108 291028 245172
rect 437796 245108 437860 245172
rect 284156 244972 284220 245036
rect 439268 244972 439332 245036
rect 283972 244836 284036 244900
rect 292436 244700 292500 244764
rect 295932 244564 295996 244628
rect 297404 244564 297468 244628
rect 292252 244428 292316 244492
rect 290596 244352 290660 244356
rect 290596 244296 290646 244352
rect 290646 244296 290660 244352
rect 290596 244292 290660 244296
rect 291700 244352 291764 244356
rect 291700 244296 291750 244352
rect 291750 244296 291764 244352
rect 291700 244292 291764 244296
rect 292068 244352 292132 244356
rect 292068 244296 292118 244352
rect 292118 244296 292132 244352
rect 292068 244292 292132 244296
rect 293172 244292 293236 244356
rect 293724 244352 293788 244356
rect 293724 244296 293774 244352
rect 293774 244296 293788 244352
rect 293724 244292 293788 244296
rect 295012 244352 295076 244356
rect 295012 244296 295062 244352
rect 295062 244296 295076 244352
rect 295012 244292 295076 244296
rect 297220 244292 297284 244356
rect 298692 244428 298756 244492
rect 298324 244352 298388 244356
rect 298324 244296 298374 244352
rect 298374 244296 298388 244352
rect 298324 244292 298388 244296
rect 293172 196012 293236 196076
rect 284524 169764 284588 169828
rect 295012 168404 295076 168468
rect 297220 167044 297284 167108
rect 298692 167044 298756 167108
rect 277532 160652 277596 160716
rect 160934 159896 160998 159900
rect 160934 159840 160982 159896
rect 160982 159840 160998 159896
rect 160934 159836 160998 159840
rect 163518 159896 163582 159900
rect 163518 159840 163558 159896
rect 163558 159840 163582 159896
rect 163518 159836 163582 159840
rect 165966 159896 166030 159900
rect 165966 159840 165986 159896
rect 165986 159840 166030 159896
rect 165966 159836 166030 159840
rect 203366 159836 203430 159900
rect 345974 159896 346038 159900
rect 345974 159840 345994 159896
rect 345994 159840 346038 159896
rect 345974 159836 346038 159840
rect 348286 159896 348350 159900
rect 348286 159840 348294 159896
rect 348294 159840 348350 159896
rect 348286 159836 348350 159840
rect 353590 159896 353654 159900
rect 353590 159840 353630 159896
rect 353630 159840 353654 159896
rect 353590 159836 353654 159840
rect 365966 159836 366030 159900
rect 351006 159760 351070 159764
rect 351006 159704 351054 159760
rect 351054 159704 351070 159760
rect 351006 159700 351070 159704
rect 356038 159624 356102 159628
rect 356038 159568 356058 159624
rect 356058 159568 356102 159624
rect 356038 159564 356102 159568
rect 358486 159624 358550 159628
rect 358486 159568 358506 159624
rect 358506 159568 358550 159624
rect 358486 159564 358550 159568
rect 298140 159292 298204 159356
rect 153700 159156 153764 159220
rect 128308 159020 128372 159084
rect 287652 159020 287716 159084
rect 173388 158884 173452 158948
rect 286180 158884 286244 158948
rect 287836 158884 287900 158948
rect 288940 158884 289004 158948
rect 156092 158748 156156 158812
rect 282132 158748 282196 158812
rect 284708 158748 284772 158812
rect 286364 158748 286428 158812
rect 288020 158748 288084 158812
rect 289124 158748 289188 158812
rect 290596 158808 290660 158812
rect 290596 158752 290646 158808
rect 290646 158752 290660 158808
rect 290596 158748 290660 158752
rect 291700 158748 291764 158812
rect 116164 158612 116228 158676
rect 119660 158672 119724 158676
rect 119660 158616 119710 158672
rect 119710 158616 119724 158672
rect 119660 158612 119724 158616
rect 120580 158612 120644 158676
rect 121868 158612 121932 158676
rect 123156 158672 123220 158676
rect 123156 158616 123206 158672
rect 123206 158616 123220 158672
rect 123156 158612 123220 158616
rect 124260 158612 124324 158676
rect 126468 158672 126532 158676
rect 126468 158616 126518 158672
rect 126518 158616 126532 158672
rect 126468 158612 126532 158616
rect 127572 158672 127636 158676
rect 127572 158616 127622 158672
rect 127622 158616 127636 158672
rect 127572 158612 127636 158616
rect 128676 158672 128740 158676
rect 128676 158616 128726 158672
rect 128726 158616 128740 158672
rect 128676 158612 128740 158616
rect 130148 158672 130212 158676
rect 130148 158616 130198 158672
rect 130198 158616 130212 158672
rect 130148 158612 130212 158616
rect 131252 158672 131316 158676
rect 131252 158616 131302 158672
rect 131302 158616 131316 158672
rect 131252 158612 131316 158616
rect 132356 158672 132420 158676
rect 132356 158616 132406 158672
rect 132406 158616 132420 158672
rect 132356 158612 132420 158616
rect 133460 158672 133524 158676
rect 133460 158616 133510 158672
rect 133510 158616 133524 158672
rect 133460 158612 133524 158616
rect 134564 158612 134628 158676
rect 158116 158672 158180 158676
rect 158116 158616 158166 158672
rect 158166 158616 158180 158672
rect 158116 158612 158180 158616
rect 158484 158672 158548 158676
rect 158484 158616 158534 158672
rect 158534 158616 158548 158672
rect 158484 158612 158548 158616
rect 159220 158612 159284 158676
rect 168236 158672 168300 158676
rect 168236 158616 168286 158672
rect 168286 158616 168300 158672
rect 168236 158612 168300 158616
rect 191052 158672 191116 158676
rect 191052 158616 191102 158672
rect 191102 158616 191116 158672
rect 191052 158612 191116 158616
rect 315804 158612 315868 158676
rect 317092 158612 317156 158676
rect 319484 158672 319548 158676
rect 319484 158616 319498 158672
rect 319498 158616 319548 158672
rect 319484 158612 319548 158616
rect 320588 158672 320652 158676
rect 320588 158616 320602 158672
rect 320602 158616 320652 158672
rect 320588 158612 320652 158616
rect 323164 158672 323228 158676
rect 323164 158616 323178 158672
rect 323178 158616 323228 158672
rect 323164 158612 323228 158616
rect 324268 158672 324332 158676
rect 324268 158616 324282 158672
rect 324282 158616 324332 158672
rect 324268 158612 324332 158616
rect 326476 158672 326540 158676
rect 326476 158616 326490 158672
rect 326490 158616 326540 158672
rect 326476 158612 326540 158616
rect 328316 158672 328380 158676
rect 328316 158616 328330 158672
rect 328330 158616 328380 158672
rect 328316 158612 328380 158616
rect 328684 158672 328748 158676
rect 328684 158616 328698 158672
rect 328698 158616 328748 158672
rect 328684 158612 328748 158616
rect 329972 158672 330036 158676
rect 329972 158616 329986 158672
rect 329986 158616 330036 158672
rect 329972 158612 330036 158616
rect 330708 158612 330772 158676
rect 332364 158612 332428 158676
rect 333652 158672 333716 158676
rect 333652 158616 333666 158672
rect 333666 158616 333716 158672
rect 333652 158612 333716 158616
rect 334572 158672 334636 158676
rect 334572 158616 334586 158672
rect 334586 158616 334636 158672
rect 334572 158612 334636 158616
rect 335860 158612 335924 158676
rect 336044 158672 336108 158676
rect 336044 158616 336058 158672
rect 336058 158616 336108 158672
rect 336044 158612 336108 158616
rect 336964 158612 337028 158676
rect 338436 158672 338500 158676
rect 338436 158616 338450 158672
rect 338450 158616 338500 158672
rect 338436 158612 338500 158616
rect 339356 158612 339420 158676
rect 341012 158672 341076 158676
rect 341012 158616 341026 158672
rect 341026 158616 341076 158672
rect 341012 158612 341076 158616
rect 343588 158672 343652 158676
rect 343588 158616 343602 158672
rect 343602 158616 343652 158672
rect 343588 158612 343652 158616
rect 349844 158672 349908 158676
rect 349844 158616 349858 158672
rect 349858 158616 349908 158672
rect 349844 158612 349908 158616
rect 355732 158612 355796 158676
rect 357020 158672 357084 158676
rect 357020 158616 357034 158672
rect 357034 158616 357084 158672
rect 357020 158612 357084 158616
rect 360884 158672 360948 158676
rect 360884 158616 360898 158672
rect 360898 158616 360948 158672
rect 360884 158612 360948 158616
rect 363460 158672 363524 158676
rect 363460 158616 363474 158672
rect 363474 158616 363524 158672
rect 363460 158612 363524 158616
rect 368244 158672 368308 158676
rect 368244 158616 368258 158672
rect 368258 158616 368308 158672
rect 368244 158612 368308 158616
rect 371004 158672 371068 158676
rect 371004 158616 371054 158672
rect 371054 158616 371068 158672
rect 371004 158612 371068 158616
rect 373396 158672 373460 158676
rect 373396 158616 373446 158672
rect 373446 158616 373460 158672
rect 373396 158612 373460 158616
rect 375972 158672 376036 158676
rect 375972 158616 376022 158672
rect 376022 158616 376036 158672
rect 375972 158612 376036 158616
rect 378548 158672 378612 158676
rect 378548 158616 378598 158672
rect 378598 158616 378612 158672
rect 378548 158612 378612 158616
rect 380940 158672 381004 158676
rect 380940 158616 380990 158672
rect 380990 158616 381004 158672
rect 380940 158612 381004 158616
rect 383516 158672 383580 158676
rect 383516 158616 383566 158672
rect 383566 158616 383580 158672
rect 383516 158612 383580 158616
rect 385908 158672 385972 158676
rect 385908 158616 385958 158672
rect 385958 158616 385972 158672
rect 385908 158612 385972 158616
rect 388484 158672 388548 158676
rect 388484 158616 388534 158672
rect 388534 158616 388548 158672
rect 388484 158612 388548 158616
rect 391060 158612 391124 158676
rect 393452 158672 393516 158676
rect 393452 158616 393502 158672
rect 393502 158616 393516 158672
rect 393452 158612 393516 158616
rect 395844 158672 395908 158676
rect 395844 158616 395894 158672
rect 395894 158616 395908 158672
rect 395844 158612 395908 158616
rect 398420 158672 398484 158676
rect 398420 158616 398470 158672
rect 398470 158616 398484 158672
rect 398420 158612 398484 158616
rect 400996 158612 401060 158676
rect 403388 158612 403452 158676
rect 405964 158612 406028 158676
rect 135852 158536 135916 158540
rect 135852 158480 135902 158536
rect 135902 158480 135916 158536
rect 135852 158476 135916 158480
rect 136956 158536 137020 158540
rect 136956 158480 137006 158536
rect 137006 158480 137020 158536
rect 136956 158476 137020 158480
rect 138060 158476 138124 158540
rect 139532 158476 139596 158540
rect 175964 158476 176028 158540
rect 359228 158476 359292 158540
rect 149836 158340 149900 158404
rect 178540 158340 178604 158404
rect 180932 158340 180996 158404
rect 195836 158400 195900 158404
rect 195836 158344 195886 158400
rect 195886 158344 195900 158400
rect 195836 158340 195900 158344
rect 198412 158400 198476 158404
rect 198412 158344 198462 158400
rect 198462 158344 198476 158400
rect 198412 158340 198476 158344
rect 331260 158340 331324 158404
rect 338068 158400 338132 158404
rect 338068 158344 338118 158400
rect 338118 158344 338132 158400
rect 338068 158340 338132 158344
rect 117084 158204 117148 158268
rect 141188 158204 141252 158268
rect 141740 158264 141804 158268
rect 141740 158208 141790 158264
rect 141790 158208 141804 158264
rect 141740 158204 141804 158208
rect 145972 158264 146036 158268
rect 145972 158208 146022 158264
rect 146022 158208 146036 158264
rect 145972 158204 146036 158208
rect 146340 158264 146404 158268
rect 146340 158208 146390 158264
rect 146390 158208 146404 158264
rect 146340 158204 146404 158208
rect 150940 158264 151004 158268
rect 150940 158208 150990 158264
rect 150990 158208 151004 158264
rect 150940 158204 151004 158208
rect 170996 158204 171060 158268
rect 327580 158204 327644 158268
rect 343956 158264 344020 158268
rect 343956 158208 343970 158264
rect 343970 158208 344020 158264
rect 343956 158204 344020 158208
rect 348740 158264 348804 158268
rect 348740 158208 348754 158264
rect 348754 158208 348804 158264
rect 348740 158204 348804 158208
rect 353340 158264 353404 158268
rect 353340 158208 353354 158264
rect 353354 158208 353404 158264
rect 353340 158204 353404 158208
rect 185900 158128 185964 158132
rect 185900 158072 185950 158128
rect 185950 158072 185964 158128
rect 185900 158068 185964 158072
rect 188660 158068 188724 158132
rect 333468 158068 333532 158132
rect 125364 157992 125428 157996
rect 125364 157936 125414 157992
rect 125414 157936 125428 157992
rect 125364 157932 125428 157936
rect 140636 157992 140700 157996
rect 140636 157936 140650 157992
rect 140650 157936 140700 157992
rect 140636 157932 140700 157936
rect 322060 157932 322124 157996
rect 325372 157932 325436 157996
rect 346348 157992 346412 157996
rect 346348 157936 346398 157992
rect 346398 157936 346412 157992
rect 346348 157932 346412 157936
rect 143948 157796 144012 157860
rect 145236 157856 145300 157860
rect 145236 157800 145286 157856
rect 145286 157800 145300 157856
rect 145236 157796 145300 157800
rect 148732 157856 148796 157860
rect 148732 157800 148782 157856
rect 148782 157800 148796 157856
rect 148732 157796 148796 157800
rect 193444 157796 193508 157860
rect 340644 157796 340708 157860
rect 341748 157796 341812 157860
rect 342852 157856 342916 157860
rect 342852 157800 342866 157856
rect 342866 157800 342916 157856
rect 342852 157796 342916 157800
rect 345244 157796 345308 157860
rect 347636 157796 347700 157860
rect 130700 157660 130764 157724
rect 282500 157660 282564 157724
rect 142844 157524 142908 157588
rect 147628 157524 147692 157588
rect 200988 157584 201052 157588
rect 200988 157528 201038 157584
rect 201038 157528 201052 157584
rect 200988 157524 201052 157528
rect 205956 157524 206020 157588
rect 358124 157524 358188 157588
rect 118188 157448 118252 157452
rect 118188 157392 118238 157448
rect 118238 157392 118252 157448
rect 118188 157388 118252 157392
rect 133644 157388 133708 157452
rect 136036 157448 136100 157452
rect 136036 157392 136086 157448
rect 136086 157392 136100 157448
rect 136036 157388 136100 157392
rect 138612 157388 138676 157452
rect 143580 157388 143644 157452
rect 148364 157448 148428 157452
rect 148364 157392 148414 157448
rect 148414 157392 148428 157448
rect 148364 157388 148428 157392
rect 151308 157448 151372 157452
rect 151308 157392 151358 157448
rect 151358 157392 151372 157448
rect 151308 157388 151372 157392
rect 152228 157388 152292 157452
rect 153332 157388 153396 157452
rect 154436 157448 154500 157452
rect 154436 157392 154486 157448
rect 154486 157392 154500 157448
rect 154436 157388 154500 157392
rect 155724 157448 155788 157452
rect 155724 157392 155774 157448
rect 155774 157392 155788 157448
rect 155724 157388 155788 157392
rect 157012 157448 157076 157452
rect 157012 157392 157062 157448
rect 157062 157392 157076 157448
rect 157012 157388 157076 157392
rect 183508 157388 183572 157452
rect 279372 157388 279436 157452
rect 318196 157388 318260 157452
rect 351132 157448 351196 157452
rect 351132 157392 351146 157448
rect 351146 157392 351196 157448
rect 351132 157388 351196 157392
rect 352236 157448 352300 157452
rect 352236 157392 352250 157448
rect 352250 157392 352300 157448
rect 352236 157388 352300 157392
rect 354444 157448 354508 157452
rect 354444 157392 354458 157448
rect 354458 157392 354508 157448
rect 354444 157388 354508 157392
rect 279556 155892 279620 155956
rect 286732 153716 286796 153780
rect 284892 150996 284956 151060
rect 277164 150316 277228 150380
rect 298324 75108 298388 75172
rect 439452 71844 439516 71908
rect 283972 9556 284036 9620
rect 293356 9420 293420 9484
rect 289308 9284 289372 9348
rect 295196 9148 295260 9212
rect 285076 9012 285140 9076
rect 286916 8876 286980 8940
rect 289492 8740 289556 8804
rect 298508 6836 298572 6900
rect 292436 6700 292500 6764
rect 292252 6564 292316 6628
rect 290964 6428 291028 6492
rect 288204 6292 288268 6356
rect 292068 6156 292132 6220
rect 297588 6020 297652 6084
rect 297956 4932 298020 4996
rect 297772 4796 297836 4860
rect 295932 3980 295996 4044
rect 296116 3844 296180 3908
rect 296484 3708 296548 3772
rect 439268 3708 439332 3772
rect 296300 3572 296364 3636
rect 437612 3572 437676 3636
rect 293540 3436 293604 3500
rect 437428 3436 437492 3500
rect 439084 3496 439148 3500
rect 439084 3440 439134 3496
rect 439134 3440 439148 3496
rect 439084 3436 439148 3440
rect 293724 3300 293788 3364
rect 437796 3300 437860 3364
rect 284156 3164 284220 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 245308 101414 245898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 245308 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 245308 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 245308 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 245308 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 245308 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 245308 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 245308 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 245308 137414 245898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 245308 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 245308 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 245308 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 245308 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 245308 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 245308 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 245308 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 245308 173414 245898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 245308 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 245308 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 245308 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 245308 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 245308 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 245308 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 245308 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 245308 209414 245898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 235950 479710 236116 479770
rect 237054 479710 237204 479770
rect 238158 479710 238292 479770
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 245308 213914 250398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 245308 218414 254898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 235950 476373 236010 479710
rect 235947 476372 236013 476373
rect 235947 476308 235948 476372
rect 236012 476308 236013 476372
rect 235947 476307 236013 476308
rect 237054 476237 237114 479710
rect 238158 476237 238218 479710
rect 239630 476509 239690 479710
rect 239627 476508 239693 476509
rect 239627 476444 239628 476508
rect 239692 476444 239693 476508
rect 239627 476443 239693 476444
rect 240550 476237 240610 479710
rect 241838 476237 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244474 479770
rect 243126 477053 243186 479710
rect 243123 477052 243189 477053
rect 243123 476988 243124 477052
rect 243188 476988 243189 477052
rect 243123 476987 243189 476988
rect 244414 476509 244474 479710
rect 245334 479710 245500 479770
rect 246438 479710 246588 479770
rect 247542 479710 247676 479770
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 250064 479710 250178 479770
rect 245334 476917 245394 479710
rect 245331 476916 245397 476917
rect 245331 476852 245332 476916
rect 245396 476852 245397 476916
rect 245331 476851 245397 476852
rect 244411 476508 244477 476509
rect 244411 476444 244412 476508
rect 244476 476444 244477 476508
rect 244411 476443 244477 476444
rect 246438 476237 246498 479710
rect 247542 477461 247602 479710
rect 247539 477460 247605 477461
rect 247539 477396 247540 477460
rect 247604 477396 247605 477460
rect 247539 477395 247605 477396
rect 248278 476645 248338 479710
rect 248646 477053 248706 479710
rect 250118 477461 250178 479710
rect 250670 479710 250804 479770
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 251288 479710 251466 479770
rect 250115 477460 250181 477461
rect 250115 477396 250116 477460
rect 250180 477396 250181 477460
rect 250115 477395 250181 477396
rect 248643 477052 248709 477053
rect 248643 476988 248644 477052
rect 248708 476988 248709 477052
rect 248643 476987 248709 476988
rect 248275 476644 248341 476645
rect 248275 476580 248276 476644
rect 248340 476580 248341 476644
rect 248275 476579 248341 476580
rect 250670 476509 250730 479710
rect 251406 477461 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 251403 477460 251469 477461
rect 251403 477396 251404 477460
rect 251468 477396 251469 477460
rect 251403 477395 251469 477396
rect 250667 476508 250733 476509
rect 250667 476444 250668 476508
rect 250732 476444 250733 476508
rect 250667 476443 250733 476444
rect 252326 476237 252386 479710
rect 253430 477461 253490 479710
rect 253427 477460 253493 477461
rect 253427 477396 253428 477460
rect 253492 477396 253493 477460
rect 253427 477395 253493 477396
rect 253614 476645 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 258496 479770 258556 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 253611 476644 253677 476645
rect 253611 476580 253612 476644
rect 253676 476580 253677 476644
rect 253611 476579 253677 476580
rect 254534 476373 254594 479710
rect 254531 476372 254597 476373
rect 254531 476308 254532 476372
rect 254596 476308 254597 476372
rect 254531 476307 254597 476308
rect 255822 476237 255882 479710
rect 256190 477053 256250 479710
rect 256187 477052 256253 477053
rect 256187 476988 256188 477052
rect 256252 476988 256253 477052
rect 256187 476987 256253 476988
rect 257110 476781 257170 479710
rect 257846 479710 258148 479770
rect 258398 479710 258556 479770
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 259448 479710 259562 479770
rect 260672 479710 260850 479770
rect 257846 477050 257906 479710
rect 258027 477052 258093 477053
rect 258027 477050 258028 477052
rect 257846 476990 258028 477050
rect 258027 476988 258028 476990
rect 258092 476988 258093 477052
rect 258027 476987 258093 476988
rect 258398 476781 258458 479710
rect 257107 476780 257173 476781
rect 257107 476716 257108 476780
rect 257172 476716 257173 476780
rect 257107 476715 257173 476716
rect 258395 476780 258461 476781
rect 258395 476716 258396 476780
rect 258460 476716 258461 476780
rect 258395 476715 258461 476716
rect 259502 476237 259562 479710
rect 260790 476373 260850 479710
rect 260974 479710 261140 479770
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 260974 476645 261034 479710
rect 260971 476644 261037 476645
rect 260971 476580 260972 476644
rect 261036 476580 261037 476644
rect 260971 476579 261037 476580
rect 260787 476372 260853 476373
rect 260787 476308 260788 476372
rect 260852 476308 260853 476372
rect 260787 476307 260853 476308
rect 261710 476237 261770 479710
rect 262814 476509 262874 479710
rect 263550 476645 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476644 263613 476645
rect 263547 476580 263548 476644
rect 263612 476580 263613 476644
rect 263547 476579 263613 476580
rect 262811 476508 262877 476509
rect 262811 476444 262812 476508
rect 262876 476444 262877 476508
rect 262811 476443 262877 476444
rect 263918 476373 263978 479710
rect 263915 476372 263981 476373
rect 263915 476308 263916 476372
rect 263980 476308 263981 476372
rect 263915 476307 263981 476308
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 476645 266002 479710
rect 265939 476644 266005 476645
rect 265939 476580 265940 476644
rect 266004 476580 266005 476644
rect 265939 476579 266005 476580
rect 266494 476237 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 267598 476373 267658 479710
rect 268334 477325 268394 479710
rect 268331 477324 268397 477325
rect 268331 477260 268332 477324
rect 268396 477260 268397 477324
rect 268331 477259 268397 477260
rect 267595 476372 267661 476373
rect 267595 476308 267596 476372
rect 267660 476308 267661 476372
rect 267595 476307 267661 476308
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 271144 479710 271338 479770
rect 270910 477053 270970 479710
rect 270907 477052 270973 477053
rect 270907 476988 270908 477052
rect 270972 476988 270973 477052
rect 270907 476987 270973 476988
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273486 479710 273652 479770
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 272198 476237 272258 479710
rect 273302 476373 273362 479710
rect 273486 476509 273546 479710
rect 273483 476508 273549 476509
rect 273483 476444 273484 476508
rect 273548 476444 273549 476508
rect 273483 476443 273549 476444
rect 273299 476372 273365 476373
rect 273299 476308 273300 476372
rect 273364 476308 273365 476372
rect 273299 476307 273365 476308
rect 274406 476237 274466 479710
rect 275878 476237 275938 479710
rect 276062 476373 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476372 276125 476373
rect 276059 476308 276060 476372
rect 276124 476308 276125 476372
rect 276059 476307 276125 476308
rect 276982 476237 277042 479710
rect 278086 476237 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 279168 479710 279250 479770
rect 278454 476645 278514 479710
rect 278451 476644 278517 476645
rect 278451 476580 278452 476644
rect 278516 476580 278517 476644
rect 278451 476579 278517 476580
rect 279190 476237 279250 479710
rect 280846 479710 280996 479770
rect 283422 479710 283580 479770
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 293448 479770 293508 480080
rect 285968 479710 286058 479770
rect 280846 476237 280906 479710
rect 283422 476237 283482 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293358 479710 293508 479770
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293358 476237 293418 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305870 479710 306020 479770
rect 308446 479710 308604 479770
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 318472 479770 318532 480080
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476917 303538 479710
rect 305870 477053 305930 479710
rect 308446 477053 308506 479710
rect 305867 477052 305933 477053
rect 305867 476988 305868 477052
rect 305932 476988 305933 477052
rect 305867 476987 305933 476988
rect 308443 477052 308509 477053
rect 308443 476988 308444 477052
rect 308508 476988 308509 477052
rect 308443 476987 308509 476988
rect 311022 476917 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318382 479710 318532 479770
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 320920 479710 321018 479770
rect 303475 476916 303541 476917
rect 303475 476852 303476 476916
rect 303540 476852 303541 476916
rect 303475 476851 303541 476852
rect 311019 476916 311085 476917
rect 311019 476852 311020 476916
rect 311084 476852 311085 476916
rect 311019 476851 311085 476852
rect 313414 476509 313474 479710
rect 315806 476509 315866 479710
rect 313411 476508 313477 476509
rect 313411 476444 313412 476508
rect 313476 476444 313477 476508
rect 313411 476443 313477 476444
rect 315803 476508 315869 476509
rect 315803 476444 315804 476508
rect 315868 476444 315869 476508
rect 315803 476443 315869 476444
rect 318382 476373 318442 479710
rect 320958 476373 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 476917 323410 479710
rect 325926 476917 325986 479710
rect 323347 476916 323413 476917
rect 323347 476852 323348 476916
rect 323412 476852 323413 476916
rect 323347 476851 323413 476852
rect 325923 476916 325989 476917
rect 325923 476852 325924 476916
rect 325988 476852 325989 476916
rect 325923 476851 325989 476852
rect 318379 476372 318445 476373
rect 318379 476308 318380 476372
rect 318444 476308 318445 476372
rect 318379 476307 318445 476308
rect 320955 476372 321021 476373
rect 320955 476308 320956 476372
rect 321020 476308 321021 476372
rect 320955 476307 321021 476308
rect 237051 476236 237117 476237
rect 237051 476172 237052 476236
rect 237116 476172 237117 476236
rect 237051 476171 237117 476172
rect 238155 476236 238221 476237
rect 238155 476172 238156 476236
rect 238220 476172 238221 476236
rect 238155 476171 238221 476172
rect 240547 476236 240613 476237
rect 240547 476172 240548 476236
rect 240612 476172 240613 476236
rect 240547 476171 240613 476172
rect 241835 476236 241901 476237
rect 241835 476172 241836 476236
rect 241900 476172 241901 476236
rect 241835 476171 241901 476172
rect 246435 476236 246501 476237
rect 246435 476172 246436 476236
rect 246500 476172 246501 476236
rect 246435 476171 246501 476172
rect 252323 476236 252389 476237
rect 252323 476172 252324 476236
rect 252388 476172 252389 476236
rect 252323 476171 252389 476172
rect 255819 476236 255885 476237
rect 255819 476172 255820 476236
rect 255884 476172 255885 476236
rect 255819 476171 255885 476172
rect 259499 476236 259565 476237
rect 259499 476172 259500 476236
rect 259564 476172 259565 476236
rect 259499 476171 259565 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 266491 476236 266557 476237
rect 266491 476172 266492 476236
rect 266556 476172 266557 476236
rect 266491 476171 266557 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 274403 476236 274469 476237
rect 274403 476172 274404 476236
rect 274468 476172 274469 476236
rect 274403 476171 274469 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278083 476236 278149 476237
rect 278083 476172 278084 476236
rect 278148 476172 278149 476236
rect 278083 476171 278149 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 280843 476236 280909 476237
rect 280843 476172 280844 476236
rect 280908 476172 280909 476236
rect 280843 476171 280909 476172
rect 283419 476236 283485 476237
rect 283419 476172 283420 476236
rect 283484 476172 283485 476236
rect 283419 476171 283485 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293355 476236 293421 476237
rect 293355 476172 293356 476236
rect 293420 476172 293421 476236
rect 293355 476171 293421 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 445423 362414 470898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 358859 442780 358925 442781
rect 358859 442716 358860 442780
rect 358924 442716 358925 442780
rect 358859 442715 358925 442716
rect 249568 439954 249888 439986
rect 249568 439718 249610 439954
rect 249846 439718 249888 439954
rect 249568 439634 249888 439718
rect 249568 439398 249610 439634
rect 249846 439398 249888 439634
rect 249568 439366 249888 439398
rect 280288 439954 280608 439986
rect 280288 439718 280330 439954
rect 280566 439718 280608 439954
rect 280288 439634 280608 439718
rect 280288 439398 280330 439634
rect 280566 439398 280608 439634
rect 280288 439366 280608 439398
rect 311008 439954 311328 439986
rect 311008 439718 311050 439954
rect 311286 439718 311328 439954
rect 311008 439634 311328 439718
rect 311008 439398 311050 439634
rect 311286 439398 311328 439634
rect 311008 439366 311328 439398
rect 341728 439954 342048 439986
rect 341728 439718 341770 439954
rect 342006 439718 342048 439954
rect 341728 439634 342048 439718
rect 341728 439398 341770 439634
rect 342006 439398 342048 439634
rect 341728 439366 342048 439398
rect 234208 435454 234528 435486
rect 234208 435218 234250 435454
rect 234486 435218 234528 435454
rect 234208 435134 234528 435218
rect 234208 434898 234250 435134
rect 234486 434898 234528 435134
rect 234208 434866 234528 434898
rect 264928 435454 265248 435486
rect 264928 435218 264970 435454
rect 265206 435218 265248 435454
rect 264928 435134 265248 435218
rect 264928 434898 264970 435134
rect 265206 434898 265248 435134
rect 264928 434866 265248 434898
rect 295648 435454 295968 435486
rect 295648 435218 295690 435454
rect 295926 435218 295968 435454
rect 295648 435134 295968 435218
rect 295648 434898 295690 435134
rect 295926 434898 295968 435134
rect 295648 434866 295968 434898
rect 326368 435454 326688 435486
rect 326368 435218 326410 435454
rect 326646 435218 326688 435454
rect 326368 435134 326688 435218
rect 326368 434898 326410 435134
rect 326646 434898 326688 435134
rect 326368 434866 326688 434898
rect 357088 435454 357408 435486
rect 357088 435218 357130 435454
rect 357366 435218 357408 435454
rect 357088 435134 357408 435218
rect 357088 434898 357130 435134
rect 357366 434898 357408 435134
rect 357088 434866 357408 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 249568 403954 249888 403986
rect 249568 403718 249610 403954
rect 249846 403718 249888 403954
rect 249568 403634 249888 403718
rect 249568 403398 249610 403634
rect 249846 403398 249888 403634
rect 249568 403366 249888 403398
rect 280288 403954 280608 403986
rect 280288 403718 280330 403954
rect 280566 403718 280608 403954
rect 280288 403634 280608 403718
rect 280288 403398 280330 403634
rect 280566 403398 280608 403634
rect 280288 403366 280608 403398
rect 311008 403954 311328 403986
rect 311008 403718 311050 403954
rect 311286 403718 311328 403954
rect 311008 403634 311328 403718
rect 311008 403398 311050 403634
rect 311286 403398 311328 403634
rect 311008 403366 311328 403398
rect 341728 403954 342048 403986
rect 341728 403718 341770 403954
rect 342006 403718 342048 403954
rect 341728 403634 342048 403718
rect 341728 403398 341770 403634
rect 342006 403398 342048 403634
rect 341728 403366 342048 403398
rect 234208 399454 234528 399486
rect 234208 399218 234250 399454
rect 234486 399218 234528 399454
rect 234208 399134 234528 399218
rect 234208 398898 234250 399134
rect 234486 398898 234528 399134
rect 234208 398866 234528 398898
rect 264928 399454 265248 399486
rect 264928 399218 264970 399454
rect 265206 399218 265248 399454
rect 264928 399134 265248 399218
rect 264928 398898 264970 399134
rect 265206 398898 265248 399134
rect 264928 398866 265248 398898
rect 295648 399454 295968 399486
rect 295648 399218 295690 399454
rect 295926 399218 295968 399454
rect 295648 399134 295968 399218
rect 295648 398898 295690 399134
rect 295926 398898 295968 399134
rect 295648 398866 295968 398898
rect 326368 399454 326688 399486
rect 326368 399218 326410 399454
rect 326646 399218 326688 399454
rect 326368 399134 326688 399218
rect 326368 398898 326410 399134
rect 326646 398898 326688 399134
rect 326368 398866 326688 398898
rect 357088 399454 357408 399486
rect 357088 399218 357130 399454
rect 357366 399218 357408 399454
rect 357088 399134 357408 399218
rect 357088 398898 357130 399134
rect 357366 398898 357408 399134
rect 357088 398866 357408 398898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 249568 367954 249888 367986
rect 249568 367718 249610 367954
rect 249846 367718 249888 367954
rect 249568 367634 249888 367718
rect 249568 367398 249610 367634
rect 249846 367398 249888 367634
rect 249568 367366 249888 367398
rect 280288 367954 280608 367986
rect 280288 367718 280330 367954
rect 280566 367718 280608 367954
rect 280288 367634 280608 367718
rect 280288 367398 280330 367634
rect 280566 367398 280608 367634
rect 280288 367366 280608 367398
rect 311008 367954 311328 367986
rect 311008 367718 311050 367954
rect 311286 367718 311328 367954
rect 311008 367634 311328 367718
rect 311008 367398 311050 367634
rect 311286 367398 311328 367634
rect 311008 367366 311328 367398
rect 341728 367954 342048 367986
rect 341728 367718 341770 367954
rect 342006 367718 342048 367954
rect 341728 367634 342048 367718
rect 341728 367398 341770 367634
rect 342006 367398 342048 367634
rect 341728 367366 342048 367398
rect 234208 363454 234528 363486
rect 234208 363218 234250 363454
rect 234486 363218 234528 363454
rect 234208 363134 234528 363218
rect 234208 362898 234250 363134
rect 234486 362898 234528 363134
rect 234208 362866 234528 362898
rect 264928 363454 265248 363486
rect 264928 363218 264970 363454
rect 265206 363218 265248 363454
rect 264928 363134 265248 363218
rect 264928 362898 264970 363134
rect 265206 362898 265248 363134
rect 264928 362866 265248 362898
rect 295648 363454 295968 363486
rect 295648 363218 295690 363454
rect 295926 363218 295968 363454
rect 295648 363134 295968 363218
rect 295648 362898 295690 363134
rect 295926 362898 295968 363134
rect 295648 362866 295968 362898
rect 326368 363454 326688 363486
rect 326368 363218 326410 363454
rect 326646 363218 326688 363454
rect 326368 363134 326688 363218
rect 326368 362898 326410 363134
rect 326646 362898 326688 363134
rect 326368 362866 326688 362898
rect 357088 363454 357408 363486
rect 357088 363218 357130 363454
rect 357366 363218 357408 363454
rect 357088 363134 357408 363218
rect 357088 362898 357130 363134
rect 357366 362898 357408 363134
rect 357088 362866 357408 362898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 249568 331954 249888 331986
rect 249568 331718 249610 331954
rect 249846 331718 249888 331954
rect 249568 331634 249888 331718
rect 249568 331398 249610 331634
rect 249846 331398 249888 331634
rect 249568 331366 249888 331398
rect 280288 331954 280608 331986
rect 280288 331718 280330 331954
rect 280566 331718 280608 331954
rect 280288 331634 280608 331718
rect 280288 331398 280330 331634
rect 280566 331398 280608 331634
rect 280288 331366 280608 331398
rect 311008 331954 311328 331986
rect 311008 331718 311050 331954
rect 311286 331718 311328 331954
rect 311008 331634 311328 331718
rect 311008 331398 311050 331634
rect 311286 331398 311328 331634
rect 311008 331366 311328 331398
rect 341728 331954 342048 331986
rect 341728 331718 341770 331954
rect 342006 331718 342048 331954
rect 341728 331634 342048 331718
rect 341728 331398 341770 331634
rect 342006 331398 342048 331634
rect 341728 331366 342048 331398
rect 234208 327454 234528 327486
rect 234208 327218 234250 327454
rect 234486 327218 234528 327454
rect 234208 327134 234528 327218
rect 234208 326898 234250 327134
rect 234486 326898 234528 327134
rect 234208 326866 234528 326898
rect 264928 327454 265248 327486
rect 264928 327218 264970 327454
rect 265206 327218 265248 327454
rect 264928 327134 265248 327218
rect 264928 326898 264970 327134
rect 265206 326898 265248 327134
rect 264928 326866 265248 326898
rect 295648 327454 295968 327486
rect 295648 327218 295690 327454
rect 295926 327218 295968 327454
rect 295648 327134 295968 327218
rect 295648 326898 295690 327134
rect 295926 326898 295968 327134
rect 295648 326866 295968 326898
rect 326368 327454 326688 327486
rect 326368 327218 326410 327454
rect 326646 327218 326688 327454
rect 326368 327134 326688 327218
rect 326368 326898 326410 327134
rect 326646 326898 326688 327134
rect 326368 326866 326688 326898
rect 357088 327454 357408 327486
rect 357088 327218 357130 327454
rect 357366 327218 357408 327454
rect 357088 327134 357408 327218
rect 357088 326898 357130 327134
rect 357366 326898 357408 327134
rect 357088 326866 357408 326898
rect 295195 309092 295261 309093
rect 295195 309028 295196 309092
rect 295260 309028 295261 309092
rect 295195 309027 295261 309028
rect 282131 308820 282197 308821
rect 282131 308756 282132 308820
rect 282196 308756 282197 308820
rect 282131 308755 282197 308756
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 240294 277954 240914 308400
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 100272 223954 100620 223986
rect 100272 223718 100328 223954
rect 100564 223718 100620 223954
rect 100272 223634 100620 223718
rect 100272 223398 100328 223634
rect 100564 223398 100620 223634
rect 100272 223366 100620 223398
rect 236000 223954 236348 223986
rect 236000 223718 236056 223954
rect 236292 223718 236348 223954
rect 236000 223634 236348 223718
rect 236000 223398 236056 223634
rect 236292 223398 236348 223634
rect 236000 223366 236348 223398
rect 100952 219454 101300 219486
rect 100952 219218 101008 219454
rect 101244 219218 101300 219454
rect 100952 219134 101300 219218
rect 100952 218898 101008 219134
rect 101244 218898 101300 219134
rect 100952 218866 101300 218898
rect 235320 219454 235668 219486
rect 235320 219218 235376 219454
rect 235612 219218 235668 219454
rect 235320 219134 235668 219218
rect 235320 218898 235376 219134
rect 235612 218898 235668 219134
rect 235320 218866 235668 218898
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 100272 187954 100620 187986
rect 100272 187718 100328 187954
rect 100564 187718 100620 187954
rect 100272 187634 100620 187718
rect 100272 187398 100328 187634
rect 100564 187398 100620 187634
rect 100272 187366 100620 187398
rect 236000 187954 236348 187986
rect 236000 187718 236056 187954
rect 236292 187718 236348 187954
rect 236000 187634 236348 187718
rect 236000 187398 236056 187634
rect 236292 187398 236348 187634
rect 236000 187366 236348 187398
rect 100952 183454 101300 183486
rect 100952 183218 101008 183454
rect 101244 183218 101300 183454
rect 100952 183134 101300 183218
rect 100952 182898 101008 183134
rect 101244 182898 101300 183134
rect 100952 182866 101300 182898
rect 235320 183454 235668 183486
rect 235320 183218 235376 183454
rect 235612 183218 235668 183454
rect 235320 183134 235668 183218
rect 235320 182898 235376 183134
rect 235612 182898 235668 183134
rect 235320 182866 235668 182898
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 116056 159490 116116 160106
rect 117144 159490 117204 160106
rect 118232 159490 118292 160106
rect 116056 159430 116226 159490
rect 116166 158677 116226 159430
rect 117086 159430 117204 159490
rect 118190 159430 118292 159490
rect 119592 159490 119652 160106
rect 120544 159490 120604 160106
rect 121768 159490 121828 160106
rect 123128 159490 123188 160106
rect 124216 159490 124276 160106
rect 125440 159490 125500 160106
rect 126528 159490 126588 160106
rect 127616 159490 127676 160106
rect 119592 159430 119722 159490
rect 120544 159430 120642 159490
rect 121768 159430 121930 159490
rect 123128 159430 123218 159490
rect 124216 159430 124322 159490
rect 116163 158676 116229 158677
rect 116163 158612 116164 158676
rect 116228 158612 116229 158676
rect 116163 158611 116229 158612
rect 117086 158269 117146 159430
rect 117083 158268 117149 158269
rect 117083 158204 117084 158268
rect 117148 158204 117149 158268
rect 117083 158203 117149 158204
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 138454 101414 158000
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 142954 105914 158000
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 147454 110414 158000
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 151954 114914 158000
rect 118190 157453 118250 159430
rect 119662 158677 119722 159430
rect 120582 158677 120642 159430
rect 121870 158677 121930 159430
rect 123158 158677 123218 159430
rect 124262 158677 124322 159430
rect 125366 159430 125500 159490
rect 126470 159430 126588 159490
rect 127574 159430 127676 159490
rect 128296 159490 128356 160106
rect 128704 159490 128764 160106
rect 128296 159430 128370 159490
rect 119659 158676 119725 158677
rect 119659 158612 119660 158676
rect 119724 158612 119725 158676
rect 119659 158611 119725 158612
rect 120579 158676 120645 158677
rect 120579 158612 120580 158676
rect 120644 158612 120645 158676
rect 120579 158611 120645 158612
rect 121867 158676 121933 158677
rect 121867 158612 121868 158676
rect 121932 158612 121933 158676
rect 121867 158611 121933 158612
rect 123155 158676 123221 158677
rect 123155 158612 123156 158676
rect 123220 158612 123221 158676
rect 123155 158611 123221 158612
rect 124259 158676 124325 158677
rect 124259 158612 124260 158676
rect 124324 158612 124325 158676
rect 124259 158611 124325 158612
rect 118187 157452 118253 157453
rect 118187 157388 118188 157452
rect 118252 157388 118253 157452
rect 118187 157387 118253 157388
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 156454 119414 158000
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 124954 123914 158000
rect 125366 157997 125426 159430
rect 126470 158677 126530 159430
rect 127574 158677 127634 159430
rect 128310 159085 128370 159430
rect 128678 159430 128764 159490
rect 130064 159490 130124 160106
rect 130744 159490 130804 160106
rect 131288 159490 131348 160106
rect 132376 159490 132436 160106
rect 133464 159490 133524 160106
rect 130064 159430 130210 159490
rect 128307 159084 128373 159085
rect 128307 159020 128308 159084
rect 128372 159020 128373 159084
rect 128307 159019 128373 159020
rect 128678 158677 128738 159430
rect 130150 158677 130210 159430
rect 130702 159430 130804 159490
rect 131254 159430 131348 159490
rect 132358 159430 132436 159490
rect 133462 159430 133524 159490
rect 133600 159490 133660 160106
rect 134552 159490 134612 160106
rect 135912 159490 135972 160106
rect 136048 159490 136108 160106
rect 137000 159490 137060 160106
rect 138088 159490 138148 160106
rect 133600 159430 133706 159490
rect 134552 159430 134626 159490
rect 126467 158676 126533 158677
rect 126467 158612 126468 158676
rect 126532 158612 126533 158676
rect 126467 158611 126533 158612
rect 127571 158676 127637 158677
rect 127571 158612 127572 158676
rect 127636 158612 127637 158676
rect 127571 158611 127637 158612
rect 128675 158676 128741 158677
rect 128675 158612 128676 158676
rect 128740 158612 128741 158676
rect 128675 158611 128741 158612
rect 130147 158676 130213 158677
rect 130147 158612 130148 158676
rect 130212 158612 130213 158676
rect 130147 158611 130213 158612
rect 125363 157996 125429 157997
rect 125363 157932 125364 157996
rect 125428 157932 125429 157996
rect 125363 157931 125429 157932
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 129454 128414 158000
rect 130702 157725 130762 159430
rect 131254 158677 131314 159430
rect 132358 158677 132418 159430
rect 133462 158677 133522 159430
rect 131251 158676 131317 158677
rect 131251 158612 131252 158676
rect 131316 158612 131317 158676
rect 131251 158611 131317 158612
rect 132355 158676 132421 158677
rect 132355 158612 132356 158676
rect 132420 158612 132421 158676
rect 132355 158611 132421 158612
rect 133459 158676 133525 158677
rect 133459 158612 133460 158676
rect 133524 158612 133525 158676
rect 133459 158611 133525 158612
rect 130699 157724 130765 157725
rect 130699 157660 130700 157724
rect 130764 157660 130765 157724
rect 130699 157659 130765 157660
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 133954 132914 158000
rect 133646 157453 133706 159430
rect 134566 158677 134626 159430
rect 135854 159430 135972 159490
rect 136038 159430 136108 159490
rect 136958 159430 137060 159490
rect 138062 159430 138148 159490
rect 138496 159490 138556 160106
rect 139448 159490 139508 160106
rect 140672 159490 140732 160106
rect 138496 159430 138674 159490
rect 139448 159430 139594 159490
rect 134563 158676 134629 158677
rect 134563 158612 134564 158676
rect 134628 158612 134629 158676
rect 134563 158611 134629 158612
rect 135854 158541 135914 159430
rect 135851 158540 135917 158541
rect 135851 158476 135852 158540
rect 135916 158476 135917 158540
rect 135851 158475 135917 158476
rect 136038 157453 136098 159430
rect 136958 158541 137018 159430
rect 138062 158541 138122 159430
rect 136955 158540 137021 158541
rect 136955 158476 136956 158540
rect 137020 158476 137021 158540
rect 136955 158475 137021 158476
rect 138059 158540 138125 158541
rect 138059 158476 138060 158540
rect 138124 158476 138125 158540
rect 138059 158475 138125 158476
rect 133643 157452 133709 157453
rect 133643 157388 133644 157452
rect 133708 157388 133709 157452
rect 133643 157387 133709 157388
rect 136035 157452 136101 157453
rect 136035 157388 136036 157452
rect 136100 157388 136101 157452
rect 136035 157387 136101 157388
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 138454 137414 158000
rect 138614 157453 138674 159430
rect 139534 158541 139594 159430
rect 140638 159430 140732 159490
rect 141080 159490 141140 160106
rect 141760 159490 141820 160106
rect 142848 159490 142908 160106
rect 141080 159430 141250 159490
rect 139531 158540 139597 158541
rect 139531 158476 139532 158540
rect 139596 158476 139597 158540
rect 139531 158475 139597 158476
rect 140638 157997 140698 159430
rect 141190 158269 141250 159430
rect 141742 159430 141820 159490
rect 142846 159430 142908 159490
rect 143528 159490 143588 160106
rect 143936 159490 143996 160106
rect 145296 159490 145356 160106
rect 145976 159490 146036 160106
rect 146384 159490 146444 160106
rect 143528 159430 143642 159490
rect 143936 159430 144010 159490
rect 141742 158269 141802 159430
rect 141187 158268 141253 158269
rect 141187 158204 141188 158268
rect 141252 158204 141253 158268
rect 141187 158203 141253 158204
rect 141739 158268 141805 158269
rect 141739 158204 141740 158268
rect 141804 158204 141805 158268
rect 141739 158203 141805 158204
rect 140635 157996 140701 157997
rect 140635 157932 140636 157996
rect 140700 157932 140701 157996
rect 140635 157931 140701 157932
rect 138611 157452 138677 157453
rect 138611 157388 138612 157452
rect 138676 157388 138677 157452
rect 138611 157387 138677 157388
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 142954 141914 158000
rect 142846 157589 142906 159430
rect 142843 157588 142909 157589
rect 142843 157524 142844 157588
rect 142908 157524 142909 157588
rect 142843 157523 142909 157524
rect 143582 157453 143642 159430
rect 143950 157861 144010 159430
rect 145238 159430 145356 159490
rect 145974 159430 146036 159490
rect 146342 159430 146444 159490
rect 147608 159490 147668 160106
rect 148288 159490 148348 160106
rect 148696 159490 148756 160106
rect 149784 159490 149844 160106
rect 151008 159490 151068 160106
rect 147608 159430 147690 159490
rect 148288 159430 148426 159490
rect 148696 159430 148794 159490
rect 149784 159430 149898 159490
rect 145238 157861 145298 159430
rect 145974 158269 146034 159430
rect 146342 158269 146402 159430
rect 145971 158268 146037 158269
rect 145971 158204 145972 158268
rect 146036 158204 146037 158268
rect 145971 158203 146037 158204
rect 146339 158268 146405 158269
rect 146339 158204 146340 158268
rect 146404 158204 146405 158268
rect 146339 158203 146405 158204
rect 143947 157860 144013 157861
rect 143947 157796 143948 157860
rect 144012 157796 144013 157860
rect 143947 157795 144013 157796
rect 145235 157860 145301 157861
rect 145235 157796 145236 157860
rect 145300 157796 145301 157860
rect 145235 157795 145301 157796
rect 143579 157452 143645 157453
rect 143579 157388 143580 157452
rect 143644 157388 143645 157452
rect 143579 157387 143645 157388
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 147454 146414 158000
rect 147630 157589 147690 159430
rect 147627 157588 147693 157589
rect 147627 157524 147628 157588
rect 147692 157524 147693 157588
rect 147627 157523 147693 157524
rect 148366 157453 148426 159430
rect 148734 157861 148794 159430
rect 149838 158405 149898 159430
rect 150942 159430 151068 159490
rect 151144 159490 151204 160106
rect 152232 159490 152292 160106
rect 151144 159430 151370 159490
rect 149835 158404 149901 158405
rect 149835 158340 149836 158404
rect 149900 158340 149901 158404
rect 149835 158339 149901 158340
rect 150942 158269 151002 159430
rect 150939 158268 151005 158269
rect 150939 158204 150940 158268
rect 151004 158204 151005 158268
rect 150939 158203 151005 158204
rect 148731 157860 148797 157861
rect 148731 157796 148732 157860
rect 148796 157796 148797 157860
rect 148731 157795 148797 157796
rect 148363 157452 148429 157453
rect 148363 157388 148364 157452
rect 148428 157388 148429 157452
rect 148363 157387 148429 157388
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 151954 150914 158000
rect 151310 157453 151370 159430
rect 152230 159430 152292 159490
rect 153320 159490 153380 160106
rect 153592 159490 153652 160106
rect 154408 159490 154468 160106
rect 155768 159490 155828 160106
rect 153320 159430 153394 159490
rect 153592 159430 153762 159490
rect 154408 159430 154498 159490
rect 152230 157453 152290 159430
rect 153334 157453 153394 159430
rect 153702 159221 153762 159430
rect 153699 159220 153765 159221
rect 153699 159156 153700 159220
rect 153764 159156 153765 159220
rect 153699 159155 153765 159156
rect 154438 157453 154498 159430
rect 155726 159430 155828 159490
rect 156040 159490 156100 160106
rect 156992 159490 157052 160106
rect 158080 159490 158140 160106
rect 158488 159490 158548 160106
rect 156040 159430 156154 159490
rect 156992 159430 157074 159490
rect 158080 159430 158178 159490
rect 151307 157452 151373 157453
rect 151307 157388 151308 157452
rect 151372 157388 151373 157452
rect 151307 157387 151373 157388
rect 152227 157452 152293 157453
rect 152227 157388 152228 157452
rect 152292 157388 152293 157452
rect 152227 157387 152293 157388
rect 153331 157452 153397 157453
rect 153331 157388 153332 157452
rect 153396 157388 153397 157452
rect 153331 157387 153397 157388
rect 154435 157452 154501 157453
rect 154435 157388 154436 157452
rect 154500 157388 154501 157452
rect 154435 157387 154501 157388
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 156454 155414 158000
rect 155726 157453 155786 159430
rect 156094 158813 156154 159430
rect 156091 158812 156157 158813
rect 156091 158748 156092 158812
rect 156156 158748 156157 158812
rect 156091 158747 156157 158748
rect 157014 157453 157074 159430
rect 158118 158677 158178 159430
rect 158486 159430 158548 159490
rect 159168 159490 159228 160106
rect 160936 159901 160996 160106
rect 163520 159901 163580 160106
rect 165968 159901 166028 160106
rect 160933 159900 160999 159901
rect 160933 159836 160934 159900
rect 160998 159836 160999 159900
rect 160933 159835 160999 159836
rect 163517 159900 163583 159901
rect 163517 159836 163518 159900
rect 163582 159836 163583 159900
rect 163517 159835 163583 159836
rect 165965 159900 166031 159901
rect 165965 159836 165966 159900
rect 166030 159836 166031 159900
rect 165965 159835 166031 159836
rect 168280 159490 168340 160106
rect 171000 159490 171060 160106
rect 173448 159490 173508 160106
rect 159168 159430 159282 159490
rect 158486 158677 158546 159430
rect 159222 158677 159282 159430
rect 168238 159430 168340 159490
rect 170998 159430 171060 159490
rect 173390 159430 173508 159490
rect 175896 159490 175956 160106
rect 178480 159490 178540 160106
rect 180928 159490 180988 160106
rect 183512 159490 183572 160106
rect 185960 159490 186020 160106
rect 175896 159430 176026 159490
rect 178480 159430 178602 159490
rect 180928 159430 180994 159490
rect 168238 158677 168298 159430
rect 158115 158676 158181 158677
rect 158115 158612 158116 158676
rect 158180 158612 158181 158676
rect 158115 158611 158181 158612
rect 158483 158676 158549 158677
rect 158483 158612 158484 158676
rect 158548 158612 158549 158676
rect 158483 158611 158549 158612
rect 159219 158676 159285 158677
rect 159219 158612 159220 158676
rect 159284 158612 159285 158676
rect 159219 158611 159285 158612
rect 168235 158676 168301 158677
rect 168235 158612 168236 158676
rect 168300 158612 168301 158676
rect 168235 158611 168301 158612
rect 170998 158269 171058 159430
rect 173390 158949 173450 159430
rect 173387 158948 173453 158949
rect 173387 158884 173388 158948
rect 173452 158884 173453 158948
rect 173387 158883 173453 158884
rect 175966 158541 176026 159430
rect 175963 158540 176029 158541
rect 175963 158476 175964 158540
rect 176028 158476 176029 158540
rect 175963 158475 176029 158476
rect 178542 158405 178602 159430
rect 180934 158405 180994 159430
rect 183510 159430 183572 159490
rect 185902 159430 186020 159490
rect 188544 159490 188604 160106
rect 190992 159490 191052 160106
rect 193440 159490 193500 160106
rect 195888 159490 195948 160106
rect 198472 159490 198532 160106
rect 188544 159430 188722 159490
rect 190992 159430 191114 159490
rect 193440 159430 193506 159490
rect 178539 158404 178605 158405
rect 178539 158340 178540 158404
rect 178604 158340 178605 158404
rect 178539 158339 178605 158340
rect 180931 158404 180997 158405
rect 180931 158340 180932 158404
rect 180996 158340 180997 158404
rect 180931 158339 180997 158340
rect 170995 158268 171061 158269
rect 170995 158204 170996 158268
rect 171060 158204 171061 158268
rect 170995 158203 171061 158204
rect 155723 157452 155789 157453
rect 155723 157388 155724 157452
rect 155788 157388 155789 157452
rect 155723 157387 155789 157388
rect 157011 157452 157077 157453
rect 157011 157388 157012 157452
rect 157076 157388 157077 157452
rect 157011 157387 157077 157388
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 124954 159914 158000
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 129454 164414 158000
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 133954 168914 158000
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 138454 173414 158000
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 142954 177914 158000
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 147454 182414 158000
rect 183510 157453 183570 159430
rect 185902 158133 185962 159430
rect 188662 158133 188722 159430
rect 191054 158677 191114 159430
rect 191051 158676 191117 158677
rect 191051 158612 191052 158676
rect 191116 158612 191117 158676
rect 191051 158611 191117 158612
rect 185899 158132 185965 158133
rect 185899 158068 185900 158132
rect 185964 158068 185965 158132
rect 185899 158067 185965 158068
rect 188659 158132 188725 158133
rect 188659 158068 188660 158132
rect 188724 158068 188725 158132
rect 188659 158067 188725 158068
rect 183507 157452 183573 157453
rect 183507 157388 183508 157452
rect 183572 157388 183573 157452
rect 183507 157387 183573 157388
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 151954 186914 158000
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 156454 191414 158000
rect 193446 157861 193506 159430
rect 195838 159430 195948 159490
rect 198414 159430 198532 159490
rect 200920 159490 200980 160106
rect 203368 159901 203428 160106
rect 203365 159900 203431 159901
rect 203365 159836 203366 159900
rect 203430 159836 203431 159900
rect 203365 159835 203431 159836
rect 205952 159490 206012 160106
rect 200920 159430 201050 159490
rect 205952 159430 206018 159490
rect 195838 158405 195898 159430
rect 198414 158405 198474 159430
rect 195835 158404 195901 158405
rect 195835 158340 195836 158404
rect 195900 158340 195901 158404
rect 195835 158339 195901 158340
rect 198411 158404 198477 158405
rect 198411 158340 198412 158404
rect 198476 158340 198477 158404
rect 198411 158339 198477 158340
rect 193443 157860 193509 157861
rect 193443 157796 193444 157860
rect 193508 157796 193509 157860
rect 193443 157795 193509 157796
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 124954 195914 158000
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 129454 200414 158000
rect 200990 157589 201050 159430
rect 200987 157588 201053 157589
rect 200987 157524 200988 157588
rect 201052 157524 201053 157588
rect 200987 157523 201053 157524
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 133954 204914 158000
rect 205958 157589 206018 159430
rect 205955 157588 206021 157589
rect 205955 157524 205956 157588
rect 206020 157524 206021 157588
rect 205955 157523 206021 157524
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 138454 209414 158000
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 142954 213914 158000
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 129454 236414 158000
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 273454 272414 308400
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 277954 276914 308400
rect 277347 308004 277413 308005
rect 277347 307940 277348 308004
rect 277412 307940 277413 308004
rect 277347 307939 277413 307940
rect 277350 302250 277410 307939
rect 277531 307868 277597 307869
rect 277531 307804 277532 307868
rect 277596 307804 277597 307868
rect 277531 307803 277597 307804
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 277166 302190 277410 302250
rect 277166 150381 277226 302190
rect 277534 160717 277594 307803
rect 279371 306236 279437 306237
rect 279371 306172 279372 306236
rect 279436 306172 279437 306236
rect 279371 306171 279437 306172
rect 277531 160716 277597 160717
rect 277531 160652 277532 160716
rect 277596 160652 277597 160716
rect 277531 160651 277597 160652
rect 279374 157453 279434 306171
rect 279555 303380 279621 303381
rect 279555 303316 279556 303380
rect 279620 303316 279621 303380
rect 279555 303315 279621 303316
rect 279371 157452 279437 157453
rect 279371 157388 279372 157452
rect 279436 157388 279437 157452
rect 279371 157387 279437 157388
rect 279558 155957 279618 303315
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 279555 155956 279621 155957
rect 279555 155892 279556 155956
rect 279620 155892 279621 155956
rect 279555 155891 279621 155892
rect 277163 150380 277229 150381
rect 277163 150316 277164 150380
rect 277228 150316 277229 150380
rect 277163 150315 277229 150316
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 138454 281414 173898
rect 282134 158813 282194 308755
rect 286179 308684 286245 308685
rect 286179 308620 286180 308684
rect 286244 308620 286245 308684
rect 286179 308619 286245 308620
rect 284891 307868 284957 307869
rect 284891 307804 284892 307868
rect 284956 307804 284957 307868
rect 284891 307803 284957 307804
rect 282499 306372 282565 306373
rect 282499 306308 282500 306372
rect 282564 306308 282565 306372
rect 282499 306307 282565 306308
rect 282131 158812 282197 158813
rect 282131 158748 282132 158812
rect 282196 158748 282197 158812
rect 282131 158747 282197 158748
rect 282502 157725 282562 306307
rect 284523 247212 284589 247213
rect 284523 247148 284524 247212
rect 284588 247148 284589 247212
rect 284523 247147 284589 247148
rect 284155 245036 284221 245037
rect 284155 244972 284156 245036
rect 284220 244972 284221 245036
rect 284155 244971 284221 244972
rect 283971 244900 284037 244901
rect 283971 244836 283972 244900
rect 284036 244836 284037 244900
rect 283971 244835 284037 244836
rect 282499 157724 282565 157725
rect 282499 157660 282500 157724
rect 282564 157660 282565 157724
rect 282499 157659 282565 157660
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 283974 9621 284034 244835
rect 283971 9620 284037 9621
rect 283971 9556 283972 9620
rect 284036 9556 284037 9620
rect 283971 9555 284037 9556
rect 284158 3229 284218 244971
rect 284526 169829 284586 247147
rect 284707 247076 284773 247077
rect 284707 247012 284708 247076
rect 284772 247012 284773 247076
rect 284707 247011 284773 247012
rect 284523 169828 284589 169829
rect 284523 169764 284524 169828
rect 284588 169764 284589 169828
rect 284523 169763 284589 169764
rect 284710 158813 284770 247011
rect 284707 158812 284773 158813
rect 284707 158748 284708 158812
rect 284772 158748 284773 158812
rect 284707 158747 284773 158748
rect 284894 151061 284954 307803
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285075 247620 285141 247621
rect 285075 247556 285076 247620
rect 285140 247556 285141 247620
rect 285075 247555 285141 247556
rect 284891 151060 284957 151061
rect 284891 150996 284892 151060
rect 284956 150996 284957 151060
rect 284891 150995 284957 150996
rect 285078 9077 285138 247555
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 286182 158949 286242 308619
rect 286731 307868 286797 307869
rect 286731 307804 286732 307868
rect 286796 307804 286797 307868
rect 286731 307803 286797 307804
rect 286363 247076 286429 247077
rect 286363 247012 286364 247076
rect 286428 247012 286429 247076
rect 286363 247011 286429 247012
rect 286179 158948 286245 158949
rect 286179 158884 286180 158948
rect 286244 158884 286245 158948
rect 286179 158883 286245 158884
rect 286366 158813 286426 247011
rect 286363 158812 286429 158813
rect 286363 158748 286364 158812
rect 286428 158748 286429 158812
rect 286363 158747 286429 158748
rect 286734 153781 286794 307803
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289491 248164 289557 248165
rect 289491 248100 289492 248164
rect 289556 248100 289557 248164
rect 289491 248099 289557 248100
rect 288203 248028 288269 248029
rect 288203 247964 288204 248028
rect 288268 247964 288269 248028
rect 288203 247963 288269 247964
rect 288019 247756 288085 247757
rect 288019 247692 288020 247756
rect 288084 247692 288085 247756
rect 288019 247691 288085 247692
rect 287651 247212 287717 247213
rect 287651 247148 287652 247212
rect 287716 247148 287717 247212
rect 287651 247147 287717 247148
rect 286915 247076 286981 247077
rect 286915 247012 286916 247076
rect 286980 247012 286981 247076
rect 286915 247011 286981 247012
rect 286731 153780 286797 153781
rect 286731 153716 286732 153780
rect 286796 153716 286797 153780
rect 286731 153715 286797 153716
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285075 9076 285141 9077
rect 285075 9012 285076 9076
rect 285140 9012 285141 9076
rect 285075 9011 285141 9012
rect 284155 3228 284221 3229
rect 284155 3164 284156 3228
rect 284220 3164 284221 3228
rect 284155 3163 284221 3164
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 -7066 285914 34398
rect 286918 8941 286978 247011
rect 287654 159085 287714 247147
rect 287835 247076 287901 247077
rect 287835 247012 287836 247076
rect 287900 247012 287901 247076
rect 287835 247011 287901 247012
rect 287651 159084 287717 159085
rect 287651 159020 287652 159084
rect 287716 159020 287717 159084
rect 287651 159019 287717 159020
rect 287838 158949 287898 247011
rect 287835 158948 287901 158949
rect 287835 158884 287836 158948
rect 287900 158884 287901 158948
rect 287835 158883 287901 158884
rect 288022 158813 288082 247691
rect 288019 158812 288085 158813
rect 288019 158748 288020 158812
rect 288084 158748 288085 158812
rect 288019 158747 288085 158748
rect 286915 8940 286981 8941
rect 286915 8876 286916 8940
rect 286980 8876 286981 8940
rect 286915 8875 286981 8876
rect 288206 6357 288266 247963
rect 289307 247892 289373 247893
rect 289307 247828 289308 247892
rect 289372 247828 289373 247892
rect 289307 247827 289373 247828
rect 288939 247212 289005 247213
rect 288939 247148 288940 247212
rect 289004 247148 289005 247212
rect 288939 247147 289005 247148
rect 288942 158949 289002 247147
rect 289123 247076 289189 247077
rect 289123 247012 289124 247076
rect 289188 247012 289189 247076
rect 289123 247011 289189 247012
rect 288939 158948 289005 158949
rect 288939 158884 288940 158948
rect 289004 158884 289005 158948
rect 288939 158883 289005 158884
rect 289126 158813 289186 247011
rect 289123 158812 289189 158813
rect 289123 158748 289124 158812
rect 289188 158748 289189 158812
rect 289123 158747 289189 158748
rect 289310 9349 289370 247827
rect 289307 9348 289373 9349
rect 289307 9284 289308 9348
rect 289372 9284 289373 9348
rect 289307 9283 289373 9284
rect 289494 8805 289554 248099
rect 289794 219454 290414 254898
rect 294294 295954 294914 308400
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 293355 248300 293421 248301
rect 293355 248236 293356 248300
rect 293420 248236 293421 248300
rect 293355 248235 293421 248236
rect 290963 245172 291029 245173
rect 290963 245108 290964 245172
rect 291028 245108 291029 245172
rect 290963 245107 291029 245108
rect 290595 244356 290661 244357
rect 290595 244292 290596 244356
rect 290660 244292 290661 244356
rect 290595 244291 290661 244292
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 290598 158813 290658 244291
rect 290595 158812 290661 158813
rect 290595 158748 290596 158812
rect 290660 158748 290661 158812
rect 290595 158747 290661 158748
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289491 8804 289557 8805
rect 289491 8740 289492 8804
rect 289556 8740 289557 8804
rect 289491 8739 289557 8740
rect 288203 6356 288269 6357
rect 288203 6292 288204 6356
rect 288268 6292 288269 6356
rect 288203 6291 288269 6292
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 3454 290414 38898
rect 290966 6493 291026 245107
rect 292435 244764 292501 244765
rect 292435 244700 292436 244764
rect 292500 244700 292501 244764
rect 292435 244699 292501 244700
rect 292251 244492 292317 244493
rect 292251 244428 292252 244492
rect 292316 244428 292317 244492
rect 292251 244427 292317 244428
rect 291699 244356 291765 244357
rect 291699 244292 291700 244356
rect 291764 244292 291765 244356
rect 291699 244291 291765 244292
rect 292067 244356 292133 244357
rect 292067 244292 292068 244356
rect 292132 244292 292133 244356
rect 292067 244291 292133 244292
rect 291702 158813 291762 244291
rect 291699 158812 291765 158813
rect 291699 158748 291700 158812
rect 291764 158748 291765 158812
rect 291699 158747 291765 158748
rect 290963 6492 291029 6493
rect 290963 6428 290964 6492
rect 291028 6428 291029 6492
rect 290963 6427 291029 6428
rect 292070 6221 292130 244291
rect 292254 6629 292314 244427
rect 292438 6765 292498 244699
rect 293171 244356 293237 244357
rect 293171 244292 293172 244356
rect 293236 244292 293237 244356
rect 293171 244291 293237 244292
rect 293174 196077 293234 244291
rect 293171 196076 293237 196077
rect 293171 196012 293172 196076
rect 293236 196012 293237 196076
rect 293171 196011 293237 196012
rect 293358 9485 293418 248235
rect 293539 245308 293605 245309
rect 293539 245244 293540 245308
rect 293604 245244 293605 245308
rect 293539 245243 293605 245244
rect 293355 9484 293421 9485
rect 293355 9420 293356 9484
rect 293420 9420 293421 9484
rect 293355 9419 293421 9420
rect 292435 6764 292501 6765
rect 292435 6700 292436 6764
rect 292500 6700 292501 6764
rect 292435 6699 292501 6700
rect 292251 6628 292317 6629
rect 292251 6564 292252 6628
rect 292316 6564 292317 6628
rect 292251 6563 292317 6564
rect 292067 6220 292133 6221
rect 292067 6156 292068 6220
rect 292132 6156 292133 6220
rect 292067 6155 292133 6156
rect 293542 3501 293602 245243
rect 293723 244356 293789 244357
rect 293723 244292 293724 244356
rect 293788 244292 293789 244356
rect 293723 244291 293789 244292
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 293539 3500 293605 3501
rect 293539 3436 293540 3500
rect 293604 3436 293605 3500
rect 293539 3435 293605 3436
rect 293726 3365 293786 244291
rect 294294 223954 294914 259398
rect 295011 244356 295077 244357
rect 295011 244292 295012 244356
rect 295076 244292 295077 244356
rect 295011 244291 295077 244292
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 295014 168469 295074 244291
rect 295011 168468 295077 168469
rect 295011 168404 295012 168468
rect 295076 168404 295077 168468
rect 295011 168403 295077 168404
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 295198 9213 295258 309027
rect 296299 308956 296365 308957
rect 296299 308892 296300 308956
rect 296364 308892 296365 308956
rect 296299 308891 296365 308892
rect 296115 247484 296181 247485
rect 296115 247420 296116 247484
rect 296180 247420 296181 247484
rect 296115 247419 296181 247420
rect 295931 244628 295997 244629
rect 295931 244564 295932 244628
rect 295996 244564 295997 244628
rect 295931 244563 295997 244564
rect 295195 9212 295261 9213
rect 295195 9148 295196 9212
rect 295260 9148 295261 9212
rect 295195 9147 295261 9148
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 293723 3364 293789 3365
rect 293723 3300 293724 3364
rect 293788 3300 293789 3364
rect 293723 3299 293789 3300
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 -1306 294914 7398
rect 295934 4045 295994 244563
rect 295931 4044 295997 4045
rect 295931 3980 295932 4044
rect 295996 3980 295997 4044
rect 295931 3979 295997 3980
rect 296118 3909 296178 247419
rect 296115 3908 296181 3909
rect 296115 3844 296116 3908
rect 296180 3844 296181 3908
rect 296115 3843 296181 3844
rect 296302 3637 296362 308891
rect 296483 308276 296549 308277
rect 296483 308212 296484 308276
rect 296548 308212 296549 308276
rect 296483 308211 296549 308212
rect 296486 3773 296546 308211
rect 297955 308140 298021 308141
rect 297955 308076 297956 308140
rect 298020 308076 298021 308140
rect 297955 308075 298021 308076
rect 297771 308004 297837 308005
rect 297771 307940 297772 308004
rect 297836 307940 297837 308004
rect 297771 307939 297837 307940
rect 297403 307868 297469 307869
rect 297403 307804 297404 307868
rect 297468 307804 297469 307868
rect 297403 307803 297469 307804
rect 297587 307868 297653 307869
rect 297587 307804 297588 307868
rect 297652 307804 297653 307868
rect 297587 307803 297653 307804
rect 297406 244629 297466 307803
rect 297403 244628 297469 244629
rect 297403 244564 297404 244628
rect 297468 244564 297469 244628
rect 297403 244563 297469 244564
rect 297219 244356 297285 244357
rect 297219 244292 297220 244356
rect 297284 244292 297285 244356
rect 297219 244291 297285 244292
rect 297222 167109 297282 244291
rect 297219 167108 297285 167109
rect 297219 167044 297220 167108
rect 297284 167044 297285 167108
rect 297219 167043 297285 167044
rect 297590 6085 297650 307803
rect 297587 6084 297653 6085
rect 297587 6020 297588 6084
rect 297652 6020 297653 6084
rect 297587 6019 297653 6020
rect 297774 4861 297834 307939
rect 297958 4997 298018 308075
rect 298139 308004 298205 308005
rect 298139 307940 298140 308004
rect 298204 307940 298205 308004
rect 298139 307939 298205 307940
rect 298142 159357 298202 307939
rect 298507 307868 298573 307869
rect 298507 307804 298508 307868
rect 298572 307804 298573 307868
rect 298507 307803 298573 307804
rect 298323 244356 298389 244357
rect 298323 244292 298324 244356
rect 298388 244292 298389 244356
rect 298323 244291 298389 244292
rect 298139 159356 298205 159357
rect 298139 159292 298140 159356
rect 298204 159292 298205 159356
rect 298139 159291 298205 159292
rect 298326 75173 298386 244291
rect 298323 75172 298389 75173
rect 298323 75108 298324 75172
rect 298388 75108 298389 75172
rect 298323 75107 298389 75108
rect 298510 6901 298570 307803
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 358862 245581 358922 442715
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 358859 245580 358925 245581
rect 358859 245516 358860 245580
rect 358924 245516 358925 245580
rect 358859 245515 358925 245516
rect 361794 245308 362414 254898
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 245308 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 245308 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 245308 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 245308 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 245308 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 245308 389414 245898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 245308 393914 250398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 245308 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 245308 402914 259398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 245308 407414 263898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 245308 411914 268398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 245308 416414 272898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 245308 420914 277398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 245308 425414 245898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 245308 429914 250398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 439451 443052 439517 443053
rect 439451 442988 439452 443052
rect 439516 442988 439517 443052
rect 439451 442987 439517 442988
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 437427 275228 437493 275229
rect 437427 275164 437428 275228
rect 437492 275164 437493 275228
rect 437427 275163 437493 275164
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 245308 434414 254898
rect 298691 244492 298757 244493
rect 298691 244428 298692 244492
rect 298756 244428 298757 244492
rect 298691 244427 298757 244428
rect 298694 167109 298754 244427
rect 300272 223954 300620 223986
rect 300272 223718 300328 223954
rect 300564 223718 300620 223954
rect 300272 223634 300620 223718
rect 300272 223398 300328 223634
rect 300564 223398 300620 223634
rect 300272 223366 300620 223398
rect 436000 223954 436348 223986
rect 436000 223718 436056 223954
rect 436292 223718 436348 223954
rect 436000 223634 436348 223718
rect 436000 223398 436056 223634
rect 436292 223398 436348 223634
rect 436000 223366 436348 223398
rect 300952 219454 301300 219486
rect 300952 219218 301008 219454
rect 301244 219218 301300 219454
rect 300952 219134 301300 219218
rect 300952 218898 301008 219134
rect 301244 218898 301300 219134
rect 300952 218866 301300 218898
rect 435320 219454 435668 219486
rect 435320 219218 435376 219454
rect 435612 219218 435668 219454
rect 435320 219134 435668 219218
rect 435320 218898 435376 219134
rect 435612 218898 435668 219134
rect 435320 218866 435668 218898
rect 300272 187954 300620 187986
rect 300272 187718 300328 187954
rect 300564 187718 300620 187954
rect 300272 187634 300620 187718
rect 300272 187398 300328 187634
rect 300564 187398 300620 187634
rect 300272 187366 300620 187398
rect 436000 187954 436348 187986
rect 436000 187718 436056 187954
rect 436292 187718 436348 187954
rect 436000 187634 436348 187718
rect 436000 187398 436056 187634
rect 436292 187398 436348 187634
rect 436000 187366 436348 187398
rect 300952 183454 301300 183486
rect 300952 183218 301008 183454
rect 301244 183218 301300 183454
rect 300952 183134 301300 183218
rect 300952 182898 301008 183134
rect 301244 182898 301300 183134
rect 300952 182866 301300 182898
rect 435320 183454 435668 183486
rect 435320 183218 435376 183454
rect 435612 183218 435668 183454
rect 435320 183134 435668 183218
rect 435320 182898 435376 183134
rect 435612 182898 435668 183134
rect 435320 182866 435668 182898
rect 298691 167108 298757 167109
rect 298691 167044 298692 167108
rect 298756 167044 298757 167108
rect 298691 167043 298757 167044
rect 316056 159490 316116 160106
rect 317144 159490 317204 160106
rect 318232 159490 318292 160106
rect 319592 159490 319652 160106
rect 315806 159430 316116 159490
rect 317094 159430 317204 159490
rect 318198 159430 318292 159490
rect 319486 159430 319652 159490
rect 320544 159490 320604 160106
rect 321768 159490 321828 160106
rect 323128 159490 323188 160106
rect 324216 159490 324276 160106
rect 325440 159490 325500 160106
rect 326528 159490 326588 160106
rect 327616 159490 327676 160106
rect 320544 159430 320650 159490
rect 321768 159430 322122 159490
rect 323128 159430 323226 159490
rect 324216 159430 324330 159490
rect 315806 158677 315866 159430
rect 317094 158677 317154 159430
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 317091 158676 317157 158677
rect 317091 158612 317092 158676
rect 317156 158612 317157 158676
rect 317091 158611 317157 158612
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298507 6900 298573 6901
rect 298507 6836 298508 6900
rect 298572 6836 298573 6900
rect 298507 6835 298573 6836
rect 297955 4996 298021 4997
rect 297955 4932 297956 4996
rect 298020 4932 298021 4996
rect 297955 4931 298021 4932
rect 297771 4860 297837 4861
rect 297771 4796 297772 4860
rect 297836 4796 297837 4860
rect 297771 4795 297837 4796
rect 296483 3772 296549 3773
rect 296483 3708 296484 3772
rect 296548 3708 296549 3772
rect 296483 3707 296549 3708
rect 296299 3636 296365 3637
rect 296299 3572 296300 3636
rect 296364 3572 296365 3636
rect 296299 3571 296365 3572
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 138454 317414 158000
rect 318198 157453 318258 159430
rect 319486 158677 319546 159430
rect 320590 158677 320650 159430
rect 319483 158676 319549 158677
rect 319483 158612 319484 158676
rect 319548 158612 319549 158676
rect 319483 158611 319549 158612
rect 320587 158676 320653 158677
rect 320587 158612 320588 158676
rect 320652 158612 320653 158676
rect 320587 158611 320653 158612
rect 318195 157452 318261 157453
rect 318195 157388 318196 157452
rect 318260 157388 318261 157452
rect 318195 157387 318261 157388
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 142954 321914 158000
rect 322062 157997 322122 159430
rect 323166 158677 323226 159430
rect 324270 158677 324330 159430
rect 325374 159430 325500 159490
rect 326478 159430 326588 159490
rect 327582 159430 327676 159490
rect 328296 159490 328356 160106
rect 328704 159490 328764 160106
rect 330064 159490 330124 160106
rect 330744 159490 330804 160106
rect 331288 159490 331348 160106
rect 332376 159490 332436 160106
rect 328296 159430 328378 159490
rect 323163 158676 323229 158677
rect 323163 158612 323164 158676
rect 323228 158612 323229 158676
rect 323163 158611 323229 158612
rect 324267 158676 324333 158677
rect 324267 158612 324268 158676
rect 324332 158612 324333 158676
rect 324267 158611 324333 158612
rect 325374 157997 325434 159430
rect 326478 158677 326538 159430
rect 326475 158676 326541 158677
rect 326475 158612 326476 158676
rect 326540 158612 326541 158676
rect 326475 158611 326541 158612
rect 327582 158269 327642 159430
rect 328318 158677 328378 159430
rect 328686 159430 328764 159490
rect 329974 159430 330124 159490
rect 330710 159430 330804 159490
rect 331262 159430 331348 159490
rect 332366 159430 332436 159490
rect 333464 159490 333524 160106
rect 333600 159490 333660 160106
rect 334552 159490 334612 160106
rect 335912 159490 335972 160106
rect 336048 159490 336108 160106
rect 337000 159490 337060 160106
rect 338088 159490 338148 160106
rect 338496 159490 338556 160106
rect 339448 159490 339508 160106
rect 340672 159490 340732 160106
rect 341080 159490 341140 160106
rect 341760 159490 341820 160106
rect 333464 159430 333530 159490
rect 333600 159430 333714 159490
rect 334552 159430 334634 159490
rect 328686 158677 328746 159430
rect 329974 158677 330034 159430
rect 330710 158677 330770 159430
rect 328315 158676 328381 158677
rect 328315 158612 328316 158676
rect 328380 158612 328381 158676
rect 328315 158611 328381 158612
rect 328683 158676 328749 158677
rect 328683 158612 328684 158676
rect 328748 158612 328749 158676
rect 328683 158611 328749 158612
rect 329971 158676 330037 158677
rect 329971 158612 329972 158676
rect 330036 158612 330037 158676
rect 329971 158611 330037 158612
rect 330707 158676 330773 158677
rect 330707 158612 330708 158676
rect 330772 158612 330773 158676
rect 330707 158611 330773 158612
rect 331262 158405 331322 159430
rect 332366 158677 332426 159430
rect 332363 158676 332429 158677
rect 332363 158612 332364 158676
rect 332428 158612 332429 158676
rect 332363 158611 332429 158612
rect 331259 158404 331325 158405
rect 331259 158340 331260 158404
rect 331324 158340 331325 158404
rect 331259 158339 331325 158340
rect 327579 158268 327645 158269
rect 327579 158204 327580 158268
rect 327644 158204 327645 158268
rect 327579 158203 327645 158204
rect 333470 158133 333530 159430
rect 333654 158677 333714 159430
rect 334574 158677 334634 159430
rect 335862 159430 335972 159490
rect 336046 159430 336108 159490
rect 336966 159430 337060 159490
rect 338070 159430 338148 159490
rect 338438 159430 338556 159490
rect 339358 159430 339508 159490
rect 340646 159430 340732 159490
rect 341014 159430 341140 159490
rect 341750 159430 341820 159490
rect 342848 159490 342908 160106
rect 343528 159490 343588 160106
rect 343936 159490 343996 160106
rect 345296 159490 345356 160106
rect 345976 159901 346036 160106
rect 345973 159900 346039 159901
rect 345973 159836 345974 159900
rect 346038 159836 346039 159900
rect 345973 159835 346039 159836
rect 346384 159490 346444 160106
rect 342848 159430 342914 159490
rect 343528 159430 343650 159490
rect 343936 159430 344018 159490
rect 335862 158677 335922 159430
rect 336046 158677 336106 159430
rect 336966 158677 337026 159430
rect 333651 158676 333717 158677
rect 333651 158612 333652 158676
rect 333716 158612 333717 158676
rect 333651 158611 333717 158612
rect 334571 158676 334637 158677
rect 334571 158612 334572 158676
rect 334636 158612 334637 158676
rect 334571 158611 334637 158612
rect 335859 158676 335925 158677
rect 335859 158612 335860 158676
rect 335924 158612 335925 158676
rect 335859 158611 335925 158612
rect 336043 158676 336109 158677
rect 336043 158612 336044 158676
rect 336108 158612 336109 158676
rect 336043 158611 336109 158612
rect 336963 158676 337029 158677
rect 336963 158612 336964 158676
rect 337028 158612 337029 158676
rect 336963 158611 337029 158612
rect 338070 158405 338130 159430
rect 338438 158677 338498 159430
rect 339358 158677 339418 159430
rect 338435 158676 338501 158677
rect 338435 158612 338436 158676
rect 338500 158612 338501 158676
rect 338435 158611 338501 158612
rect 339355 158676 339421 158677
rect 339355 158612 339356 158676
rect 339420 158612 339421 158676
rect 339355 158611 339421 158612
rect 338067 158404 338133 158405
rect 338067 158340 338068 158404
rect 338132 158340 338133 158404
rect 338067 158339 338133 158340
rect 333467 158132 333533 158133
rect 333467 158068 333468 158132
rect 333532 158068 333533 158132
rect 333467 158067 333533 158068
rect 322059 157996 322125 157997
rect 322059 157932 322060 157996
rect 322124 157932 322125 157996
rect 322059 157931 322125 157932
rect 325371 157996 325437 157997
rect 325371 157932 325372 157996
rect 325436 157932 325437 157996
rect 325371 157931 325437 157932
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 124954 339914 158000
rect 340646 157861 340706 159430
rect 341014 158677 341074 159430
rect 341011 158676 341077 158677
rect 341011 158612 341012 158676
rect 341076 158612 341077 158676
rect 341011 158611 341077 158612
rect 341750 157861 341810 159430
rect 342854 157861 342914 159430
rect 343590 158677 343650 159430
rect 343587 158676 343653 158677
rect 343587 158612 343588 158676
rect 343652 158612 343653 158676
rect 343587 158611 343653 158612
rect 343958 158269 344018 159430
rect 345246 159430 345356 159490
rect 346350 159430 346444 159490
rect 347608 159490 347668 160106
rect 348288 159901 348348 160106
rect 348285 159900 348351 159901
rect 348285 159836 348286 159900
rect 348350 159836 348351 159900
rect 348285 159835 348351 159836
rect 348696 159490 348756 160106
rect 349784 159490 349844 160106
rect 351008 159765 351068 160106
rect 351005 159764 351071 159765
rect 351005 159700 351006 159764
rect 351070 159700 351071 159764
rect 351005 159699 351071 159700
rect 351144 159490 351204 160106
rect 347608 159430 347698 159490
rect 348696 159430 348802 159490
rect 349784 159430 349906 159490
rect 343955 158268 344021 158269
rect 343955 158204 343956 158268
rect 344020 158204 344021 158268
rect 343955 158203 344021 158204
rect 340643 157860 340709 157861
rect 340643 157796 340644 157860
rect 340708 157796 340709 157860
rect 340643 157795 340709 157796
rect 341747 157860 341813 157861
rect 341747 157796 341748 157860
rect 341812 157796 341813 157860
rect 341747 157795 341813 157796
rect 342851 157860 342917 157861
rect 342851 157796 342852 157860
rect 342916 157796 342917 157860
rect 342851 157795 342917 157796
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 129454 344414 158000
rect 345246 157861 345306 159430
rect 346350 157997 346410 159430
rect 346347 157996 346413 157997
rect 346347 157932 346348 157996
rect 346412 157932 346413 157996
rect 346347 157931 346413 157932
rect 347638 157861 347698 159430
rect 348742 158269 348802 159430
rect 349846 158677 349906 159430
rect 351134 159430 351204 159490
rect 352232 159490 352292 160106
rect 353320 159490 353380 160106
rect 353592 159901 353652 160106
rect 353589 159900 353655 159901
rect 353589 159836 353590 159900
rect 353654 159836 353655 159900
rect 353589 159835 353655 159836
rect 354408 159490 354468 160106
rect 355768 159490 355828 160106
rect 356040 159629 356100 160106
rect 356037 159628 356103 159629
rect 356037 159564 356038 159628
rect 356102 159564 356103 159628
rect 356037 159563 356103 159564
rect 352232 159430 352298 159490
rect 353320 159430 353402 159490
rect 354408 159430 354506 159490
rect 349843 158676 349909 158677
rect 349843 158612 349844 158676
rect 349908 158612 349909 158676
rect 349843 158611 349909 158612
rect 348739 158268 348805 158269
rect 348739 158204 348740 158268
rect 348804 158204 348805 158268
rect 348739 158203 348805 158204
rect 345243 157860 345309 157861
rect 345243 157796 345244 157860
rect 345308 157796 345309 157860
rect 345243 157795 345309 157796
rect 347635 157860 347701 157861
rect 347635 157796 347636 157860
rect 347700 157796 347701 157860
rect 347635 157795 347701 157796
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 133954 348914 158000
rect 351134 157453 351194 159430
rect 352238 157453 352298 159430
rect 353342 158269 353402 159430
rect 353339 158268 353405 158269
rect 353339 158204 353340 158268
rect 353404 158204 353405 158268
rect 353339 158203 353405 158204
rect 351131 157452 351197 157453
rect 351131 157388 351132 157452
rect 351196 157388 351197 157452
rect 351131 157387 351197 157388
rect 352235 157452 352301 157453
rect 352235 157388 352236 157452
rect 352300 157388 352301 157452
rect 352235 157387 352301 157388
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 138454 353414 158000
rect 354446 157453 354506 159430
rect 355734 159430 355828 159490
rect 356992 159490 357052 160106
rect 358080 159490 358140 160106
rect 358488 159629 358548 160106
rect 358485 159628 358551 159629
rect 358485 159564 358486 159628
rect 358550 159564 358551 159628
rect 358485 159563 358551 159564
rect 359168 159490 359228 160106
rect 360936 159490 360996 160106
rect 363520 159490 363580 160106
rect 365968 159901 366028 160106
rect 365965 159900 366031 159901
rect 365965 159836 365966 159900
rect 366030 159836 366031 159900
rect 365965 159835 366031 159836
rect 368280 159490 368340 160106
rect 356992 159430 357082 159490
rect 358080 159430 358186 159490
rect 359168 159430 359290 159490
rect 355734 158677 355794 159430
rect 357022 158677 357082 159430
rect 355731 158676 355797 158677
rect 355731 158612 355732 158676
rect 355796 158612 355797 158676
rect 355731 158611 355797 158612
rect 357019 158676 357085 158677
rect 357019 158612 357020 158676
rect 357084 158612 357085 158676
rect 357019 158611 357085 158612
rect 354443 157452 354509 157453
rect 354443 157388 354444 157452
rect 354508 157388 354509 157452
rect 354443 157387 354509 157388
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 142954 357914 158000
rect 358126 157589 358186 159430
rect 359230 158541 359290 159430
rect 360886 159430 360996 159490
rect 363462 159430 363580 159490
rect 368246 159430 368340 159490
rect 371000 159490 371060 160106
rect 373448 159490 373508 160106
rect 371000 159430 371066 159490
rect 360886 158677 360946 159430
rect 363462 158677 363522 159430
rect 368246 158677 368306 159430
rect 371006 158677 371066 159430
rect 373398 159430 373508 159490
rect 375896 159490 375956 160106
rect 378480 159490 378540 160106
rect 380928 159490 380988 160106
rect 383512 159490 383572 160106
rect 385960 159490 386020 160106
rect 388544 159490 388604 160106
rect 375896 159430 376034 159490
rect 378480 159430 378610 159490
rect 380928 159430 381002 159490
rect 383512 159430 383578 159490
rect 373398 158677 373458 159430
rect 375974 158677 376034 159430
rect 378550 158677 378610 159430
rect 380942 158677 381002 159430
rect 383518 158677 383578 159430
rect 385910 159430 386020 159490
rect 388486 159430 388604 159490
rect 390992 159490 391052 160106
rect 393440 159490 393500 160106
rect 395888 159490 395948 160106
rect 398472 159490 398532 160106
rect 390992 159430 391122 159490
rect 393440 159430 393514 159490
rect 385910 158677 385970 159430
rect 388486 158677 388546 159430
rect 391062 158677 391122 159430
rect 393454 158677 393514 159430
rect 395846 159430 395948 159490
rect 398422 159430 398532 159490
rect 400920 159490 400980 160106
rect 403368 159490 403428 160106
rect 405952 159490 406012 160106
rect 400920 159430 401058 159490
rect 403368 159430 403450 159490
rect 405952 159430 406026 159490
rect 395846 158677 395906 159430
rect 398422 158677 398482 159430
rect 400998 158677 401058 159430
rect 403390 158677 403450 159430
rect 405966 158677 406026 159430
rect 360883 158676 360949 158677
rect 360883 158612 360884 158676
rect 360948 158612 360949 158676
rect 360883 158611 360949 158612
rect 363459 158676 363525 158677
rect 363459 158612 363460 158676
rect 363524 158612 363525 158676
rect 363459 158611 363525 158612
rect 368243 158676 368309 158677
rect 368243 158612 368244 158676
rect 368308 158612 368309 158676
rect 368243 158611 368309 158612
rect 371003 158676 371069 158677
rect 371003 158612 371004 158676
rect 371068 158612 371069 158676
rect 371003 158611 371069 158612
rect 373395 158676 373461 158677
rect 373395 158612 373396 158676
rect 373460 158612 373461 158676
rect 373395 158611 373461 158612
rect 375971 158676 376037 158677
rect 375971 158612 375972 158676
rect 376036 158612 376037 158676
rect 375971 158611 376037 158612
rect 378547 158676 378613 158677
rect 378547 158612 378548 158676
rect 378612 158612 378613 158676
rect 378547 158611 378613 158612
rect 380939 158676 381005 158677
rect 380939 158612 380940 158676
rect 381004 158612 381005 158676
rect 380939 158611 381005 158612
rect 383515 158676 383581 158677
rect 383515 158612 383516 158676
rect 383580 158612 383581 158676
rect 383515 158611 383581 158612
rect 385907 158676 385973 158677
rect 385907 158612 385908 158676
rect 385972 158612 385973 158676
rect 385907 158611 385973 158612
rect 388483 158676 388549 158677
rect 388483 158612 388484 158676
rect 388548 158612 388549 158676
rect 388483 158611 388549 158612
rect 391059 158676 391125 158677
rect 391059 158612 391060 158676
rect 391124 158612 391125 158676
rect 391059 158611 391125 158612
rect 393451 158676 393517 158677
rect 393451 158612 393452 158676
rect 393516 158612 393517 158676
rect 393451 158611 393517 158612
rect 395843 158676 395909 158677
rect 395843 158612 395844 158676
rect 395908 158612 395909 158676
rect 395843 158611 395909 158612
rect 398419 158676 398485 158677
rect 398419 158612 398420 158676
rect 398484 158612 398485 158676
rect 398419 158611 398485 158612
rect 400995 158676 401061 158677
rect 400995 158612 400996 158676
rect 401060 158612 401061 158676
rect 400995 158611 401061 158612
rect 403387 158676 403453 158677
rect 403387 158612 403388 158676
rect 403452 158612 403453 158676
rect 403387 158611 403453 158612
rect 405963 158676 406029 158677
rect 405963 158612 405964 158676
rect 406028 158612 406029 158676
rect 405963 158611 406029 158612
rect 359227 158540 359293 158541
rect 359227 158476 359228 158540
rect 359292 158476 359293 158540
rect 359227 158475 359293 158476
rect 358123 157588 358189 157589
rect 358123 157524 358124 157588
rect 358188 157524 358189 157588
rect 358123 157523 358189 157524
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 147454 362414 158000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 151954 366914 158000
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 156454 371414 158000
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 124954 375914 158000
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 129454 380414 158000
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 133954 384914 158000
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 138454 389414 158000
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 142954 393914 158000
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 147454 398414 158000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 151954 402914 158000
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 156454 407414 158000
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 124954 411914 158000
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 129454 416414 158000
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 133954 420914 158000
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 138454 425414 158000
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 142954 429914 158000
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 147454 434414 158000
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 437430 3501 437490 275163
rect 438294 259954 438914 295398
rect 439083 287740 439149 287741
rect 439083 287676 439084 287740
rect 439148 287676 439149 287740
rect 439083 287675 439149 287676
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 437611 247620 437677 247621
rect 437611 247556 437612 247620
rect 437676 247556 437677 247620
rect 437611 247555 437677 247556
rect 437614 3637 437674 247555
rect 438294 245308 438914 259398
rect 437795 245172 437861 245173
rect 437795 245108 437796 245172
rect 437860 245108 437861 245172
rect 437795 245107 437861 245108
rect 437611 3636 437677 3637
rect 437611 3572 437612 3636
rect 437676 3572 437677 3636
rect 437611 3571 437677 3572
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 437427 3500 437493 3501
rect 437427 3436 437428 3500
rect 437492 3436 437493 3500
rect 437427 3435 437493 3436
rect 437798 3365 437858 245107
rect 438294 151954 438914 158000
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 437795 3364 437861 3365
rect 437795 3300 437796 3364
rect 437860 3300 437861 3364
rect 437795 3299 437861 3300
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 -1306 438914 7398
rect 439086 3501 439146 287675
rect 439267 245036 439333 245037
rect 439267 244972 439268 245036
rect 439332 244972 439333 245036
rect 439267 244971 439333 244972
rect 439270 3773 439330 244971
rect 439454 71909 439514 442987
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 439451 71908 439517 71909
rect 439451 71844 439452 71908
rect 439516 71844 439517 71908
rect 439451 71843 439517 71844
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 439267 3772 439333 3773
rect 439267 3708 439268 3772
rect 439332 3708 439333 3772
rect 439267 3707 439333 3708
rect 439083 3500 439149 3501
rect 439083 3436 439084 3500
rect 439148 3436 439149 3500
rect 439083 3435 439149 3436
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 249610 439718 249846 439954
rect 249610 439398 249846 439634
rect 280330 439718 280566 439954
rect 280330 439398 280566 439634
rect 311050 439718 311286 439954
rect 311050 439398 311286 439634
rect 341770 439718 342006 439954
rect 341770 439398 342006 439634
rect 234250 435218 234486 435454
rect 234250 434898 234486 435134
rect 264970 435218 265206 435454
rect 264970 434898 265206 435134
rect 295690 435218 295926 435454
rect 295690 434898 295926 435134
rect 326410 435218 326646 435454
rect 326410 434898 326646 435134
rect 357130 435218 357366 435454
rect 357130 434898 357366 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 249610 403718 249846 403954
rect 249610 403398 249846 403634
rect 280330 403718 280566 403954
rect 280330 403398 280566 403634
rect 311050 403718 311286 403954
rect 311050 403398 311286 403634
rect 341770 403718 342006 403954
rect 341770 403398 342006 403634
rect 234250 399218 234486 399454
rect 234250 398898 234486 399134
rect 264970 399218 265206 399454
rect 264970 398898 265206 399134
rect 295690 399218 295926 399454
rect 295690 398898 295926 399134
rect 326410 399218 326646 399454
rect 326410 398898 326646 399134
rect 357130 399218 357366 399454
rect 357130 398898 357366 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 249610 367718 249846 367954
rect 249610 367398 249846 367634
rect 280330 367718 280566 367954
rect 280330 367398 280566 367634
rect 311050 367718 311286 367954
rect 311050 367398 311286 367634
rect 341770 367718 342006 367954
rect 341770 367398 342006 367634
rect 234250 363218 234486 363454
rect 234250 362898 234486 363134
rect 264970 363218 265206 363454
rect 264970 362898 265206 363134
rect 295690 363218 295926 363454
rect 295690 362898 295926 363134
rect 326410 363218 326646 363454
rect 326410 362898 326646 363134
rect 357130 363218 357366 363454
rect 357130 362898 357366 363134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 249610 331718 249846 331954
rect 249610 331398 249846 331634
rect 280330 331718 280566 331954
rect 280330 331398 280566 331634
rect 311050 331718 311286 331954
rect 311050 331398 311286 331634
rect 341770 331718 342006 331954
rect 341770 331398 342006 331634
rect 234250 327218 234486 327454
rect 234250 326898 234486 327134
rect 264970 327218 265206 327454
rect 264970 326898 265206 327134
rect 295690 327218 295926 327454
rect 295690 326898 295926 327134
rect 326410 327218 326646 327454
rect 326410 326898 326646 327134
rect 357130 327218 357366 327454
rect 357130 326898 357366 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 100328 223718 100564 223954
rect 100328 223398 100564 223634
rect 236056 223718 236292 223954
rect 236056 223398 236292 223634
rect 101008 219218 101244 219454
rect 101008 218898 101244 219134
rect 235376 219218 235612 219454
rect 235376 218898 235612 219134
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 100328 187718 100564 187954
rect 100328 187398 100564 187634
rect 236056 187718 236292 187954
rect 236056 187398 236292 187634
rect 101008 183218 101244 183454
rect 101008 182898 101244 183134
rect 235376 183218 235612 183454
rect 235376 182898 235612 183134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 300328 223718 300564 223954
rect 300328 223398 300564 223634
rect 436056 223718 436292 223954
rect 436056 223398 436292 223634
rect 301008 219218 301244 219454
rect 301008 218898 301244 219134
rect 435376 219218 435612 219454
rect 435376 218898 435612 219134
rect 300328 187718 300564 187954
rect 300328 187398 300564 187634
rect 436056 187718 436292 187954
rect 436056 187398 436292 187634
rect 301008 183218 301244 183454
rect 301008 182898 301244 183134
rect 435376 183218 435612 183454
rect 435376 182898 435612 183134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 249610 439954
rect 249846 439718 280330 439954
rect 280566 439718 311050 439954
rect 311286 439718 341770 439954
rect 342006 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 249610 439634
rect 249846 439398 280330 439634
rect 280566 439398 311050 439634
rect 311286 439398 341770 439634
rect 342006 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 234250 435454
rect 234486 435218 264970 435454
rect 265206 435218 295690 435454
rect 295926 435218 326410 435454
rect 326646 435218 357130 435454
rect 357366 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 234250 435134
rect 234486 434898 264970 435134
rect 265206 434898 295690 435134
rect 295926 434898 326410 435134
rect 326646 434898 357130 435134
rect 357366 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 249610 403954
rect 249846 403718 280330 403954
rect 280566 403718 311050 403954
rect 311286 403718 341770 403954
rect 342006 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 249610 403634
rect 249846 403398 280330 403634
rect 280566 403398 311050 403634
rect 311286 403398 341770 403634
rect 342006 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 234250 399454
rect 234486 399218 264970 399454
rect 265206 399218 295690 399454
rect 295926 399218 326410 399454
rect 326646 399218 357130 399454
rect 357366 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 234250 399134
rect 234486 398898 264970 399134
rect 265206 398898 295690 399134
rect 295926 398898 326410 399134
rect 326646 398898 357130 399134
rect 357366 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 249610 367954
rect 249846 367718 280330 367954
rect 280566 367718 311050 367954
rect 311286 367718 341770 367954
rect 342006 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 249610 367634
rect 249846 367398 280330 367634
rect 280566 367398 311050 367634
rect 311286 367398 341770 367634
rect 342006 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 234250 363454
rect 234486 363218 264970 363454
rect 265206 363218 295690 363454
rect 295926 363218 326410 363454
rect 326646 363218 357130 363454
rect 357366 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 234250 363134
rect 234486 362898 264970 363134
rect 265206 362898 295690 363134
rect 295926 362898 326410 363134
rect 326646 362898 357130 363134
rect 357366 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 249610 331954
rect 249846 331718 280330 331954
rect 280566 331718 311050 331954
rect 311286 331718 341770 331954
rect 342006 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 249610 331634
rect 249846 331398 280330 331634
rect 280566 331398 311050 331634
rect 311286 331398 341770 331634
rect 342006 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 234250 327454
rect 234486 327218 264970 327454
rect 265206 327218 295690 327454
rect 295926 327218 326410 327454
rect 326646 327218 357130 327454
rect 357366 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 234250 327134
rect 234486 326898 264970 327134
rect 265206 326898 295690 327134
rect 295926 326898 326410 327134
rect 326646 326898 357130 327134
rect 357366 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 100328 223954
rect 100564 223718 236056 223954
rect 236292 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 300328 223954
rect 300564 223718 436056 223954
rect 436292 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 100328 223634
rect 100564 223398 236056 223634
rect 236292 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 300328 223634
rect 300564 223398 436056 223634
rect 436292 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 101008 219454
rect 101244 219218 235376 219454
rect 235612 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 301008 219454
rect 301244 219218 435376 219454
rect 435612 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 101008 219134
rect 101244 218898 235376 219134
rect 235612 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 301008 219134
rect 301244 218898 435376 219134
rect 435612 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 100328 187954
rect 100564 187718 236056 187954
rect 236292 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 300328 187954
rect 300564 187718 436056 187954
rect 436292 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 100328 187634
rect 100564 187398 236056 187634
rect 236292 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 300328 187634
rect 300564 187398 436056 187634
rect 436292 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 101008 183454
rect 101244 183218 235376 183454
rect 235612 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 301008 183454
rect 301244 183218 435376 183454
rect 435612 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 101008 183134
rect 101244 182898 235376 183134
rect 235612 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 301008 183134
rect 301244 182898 435376 183134
rect 435612 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst_A
timestamp 0
transform 1 0 100000 0 1 160000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst_B
timestamp 0
transform 1 0 300000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 230000 0 1 310400
box 13 0 130810 133023
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 245308 110414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 245308 146414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 245308 182414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 245308 362414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 445423 362414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 245308 398414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 245308 434414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 245308 119414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 245308 155414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 245308 191414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 245308 371414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 245308 407414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 245308 128414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 245308 164414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 245308 200414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 245308 380414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 245308 416414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 245308 101414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 245308 137414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 245308 173414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 245308 209414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 565308 245414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 565308 281414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 565308 317414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 565308 353414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 245308 389414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 245308 425414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 245308 132914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 245308 168914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 245308 204914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 245308 384914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 245308 420914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 245308 105914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 245308 141914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 245308 177914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 245308 213914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 245308 393914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 245308 429914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 245308 114914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 245308 150914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 245308 186914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 245308 366914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 245308 402914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 245308 438914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 245308 123914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 245308 159914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 245308 195914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 565308 231914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 565308 267914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 565308 303914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 565308 339914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 245308 375914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 245308 411914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
